//num of or = 2675
//num of and = 22275
//num of not = 12199
//num of wire = 37147
module c1126 (in0,in1,in2,O0,O1,O2,O3,O4,O5,clk,rst);

input in0,in1,in2,clk,rst;

output O0,O1,O2,O3,O4,O5;

wire in0,in1,in2,N0,N1,N2,N3,N4,N5,N6,N7,N8,
N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,
N19,N20,N21,N22,N23,N24,N25,N26,N27,N28,
N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,
N39,N40,N41,N42,N43,N44,N45,N46,N47,N48,
N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,
N59,N60,N61,N62,N63,N64,N65,N66,N67,N68,
N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,
N79,N80,N81,N82,N83,N84,N85,N86,N87,N88,
N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,
N99,N100,N101,N102,N103,N104,N105,N106,N107,N108,
N109,N110,N111,N112,N113,N114,N115,N116,N117,N118,
N119,N120,N121,N122,N123,N124,N125,N126,N127,N128,
N129,N130,N131,N132,N133,N134,N135,N136,N137,N138,
N139,N140,N141,N142,N143,N144,N145,N146,N147,N148,
N149,N150,N151,N152,N153,N154,N155,N156,N157,N158,
N159,N160,N161,N162,N163,N164,N165,N166,N167,N168,
N169,N170,N171,N172,N173,N174,N175,N176,N177,N178,
N179,N180,N181,N182,N183,N184,N185,N186,N187,N188,
N189,N190,N191,N192,N193,N194,N195,N196,N197,N198,
N199,N200,N201,N202,N203,N204,N205,N206,N207,N208,
N209,N210,N211,N212,N213,N214,N215,N216,N217,N218,
N219,N220,N221,N222,N223,N224,N225,N226,N227,N228,
N229,N230,N231,N232,N233,N234,N235,N236,N237,N238,
N239,N240,N241,N242,N243,N244,N245,N246,N247,N248,
N249,N250,N251,N252,N253,N254,N255,N256,N257,N258,
N259,N260,N261,N262,N263,N264,N265,N266,N267,N268,
N269,N270,N271,N272,N273,N274,N275,N276,N277,N278,
N279,N280,N281,N282,N283,N284,N285,N286,N287,N288,
N289,N290,N291,N292,N293,N294,N295,N296,N297,N298,
N299,N300,N301,N302,N303,N304,N305,N306,N307,N308,
N309,N310,N311,N312,N313,N314,N315,N316,N317,N318,
N319,N320,N321,N322,N323,N324,N325,N326,N327,N328,
N329,N330,N331,N332,N333,N334,N335,N336,N337,N338,
N339,N340,N341,N342,N343,N344,N345,N346,N347,N348,
N349,N350,N351,N352,N353,N354,N355,N356,N357,N358,
N359,N360,N361,N362,N363,N364,N365,N366,N367,N368,
N369,N370,N371,N372,N373,N374,N375,N376,N377,N378,
N379,N380,N381,N382,N383,N384,N385,N386,N387,N388,
N389,N390,N391,N392,N393,N394,N395,N396,N397,N398,
N399,N400,N401,N402,N403,N404,N405,N406,N407,N408,
N409,N410,N411,N412,N413,N414,N415,N416,N417,N418,
N419,N420,N421,N422,N423,N424,N425,N426,N427,N428,
N429,N430,N431,N432,N433,N434,N435,N436,N437,N438,
N439,N440,N441,N442,N443,N444,N445,N446,N447,N448,
N449,N450,N451,N452,N453,N454,N455,N456,N457,N458,
N459,N460,N461,N462,N463,N464,N465,N466,N467,N468,
N469,N470,N471,N472,N473,N474,N475,N476,N477,N478,
N479,N480,N481,N482,N483,N484,N485,N486,N487,N488,
N489,N490,N491,N492,N493,N494,N495,N496,N497,N498,
N499,N500,N501,N502,N503,N504,N505,N506,N507,N508,
N509,N510,N511,N512,N513,N514,N515,N516,N517,N518,
N519,N520,N521,N522,N523,N524,N525,N526,N527,N528,
N529,N530,N531,N532,N533,N534,N535,N536,N537,N538,
N539,N540,N541,N542,N543,N544,N545,N546,N547,N548,
N549,N550,N551,N552,N553,N554,N555,N556,N557,N558,
N559,N560,N561,N562,N563,N564,N565,N566,N567,N568,
N569,N570,N571,N572,N573,N574,N575,N576,N577,N578,
N579,N580,N581,N582,N583,N584,N585,N586,N587,N588,
N589,N590,N591,N592,N593,N594,N595,N596,N597,N598,
N599,N600,N601,N602,N603,N604,N605,N606,N607,N608,
N609,N610,N611,N612,N613,N614,N615,N616,N617,N618,
N619,N620,N621,N622,N623,N624,N625,N626,N627,N628,
N629,N630,N631,N632,N633,N634,N635,N636,N637,N638,
N639,N640,N641,N642,N643,N644,N645,N646,N647,N648,
N649,N650,N651,N652,N653,N654,N655,N656,N657,N658,
N659,N660,N661,N662,N663,N664,N665,N666,N667,N668,
N669,N670,N671,N672,N673,N674,N675,N676,N677,N678,
N679,N680,N681,N682,N683,N684,N685,N686,N687,N688,
N689,N690,N691,N692,N693,N694,N695,N696,N697,N698,
N699,N700,N701,N702,N703,N704,N705,N706,N707,N708,
N709,N710,N711,N712,N713,N714,N715,N716,N717,N718,
N719,N720,N721,N722,N723,N724,N725,N726,N727,N728,
N729,N730,N731,N732,N733,N734,N735,N736,N737,N738,
N739,N740,N741,N742,N743,N744,N745,N746,N747,N748,
N749,N750,N751,N752,N753,N754,N755,N756,N757,N758,
N759,N760,N761,N762,N763,N764,N765,N766,N767,N768,
N769,N770,N771,N772,N773,N774,N775,N776,N777,N778,
N779,N780,N781,N782,N783,N784,N785,N786,N787,N788,
N789,N790,N791,N792,N793,N794,N795,N796,N797,N798,
N799,N800,N801,N802,N803,N804,N805,N806,N807,N808,
N809,N810,N811,N812,N813,N814,N815,N816,N817,N818,
N819,N820,N821,N822,N823,N824,N825,N826,N827,N828,
N829,N830,N831,N832,N833,N834,N835,N836,N837,N838,
N839,N840,N841,N842,N843,N844,N845,N846,N847,N848,
N849,N850,N851,N852,N853,N854,N855,N856,N857,N858,
N859,N860,N861,N862,N863,N864,N865,N866,N867,N868,
N869,N870,N871,N872,N873,N874,N875,N876,N877,N878,
N879,N880,N881,N882,N883,N884,N885,N886,N887,N888,
N889,N890,N891,N892,N893,N894,N895,N896,N897,N898,
N899,N900,N901,N902,N903,N904,N905,N906,N907,N908,
N909,N910,N911,N912,N913,N914,N915,N916,N917,N918,
N919,N920,N921,N922,N923,N924,N925,N926,N927,N928,
N929,N930,N931,N932,N933,N934,N935,N936,N937,N938,
N939,N940,N941,N942,N943,N944,N945,N946,N947,N948,
N949,N950,N951,N952,N953,N954,N955,N956,N957,N958,
N959,N960,N961,N962,N963,N964,N965,N966,N967,N968,
N969,N970,N971,N972,N973,N974,N975,N976,N977,N978,
N979,N980,N981,N982,N983,N984,N985,N986,N987,N988,
N989,N990,N991,N992,N993,N994,N995,N996,N997,N998,
N999,N1000,N1001,N1002,N1003,N1004,N1005,N1006,N1007,N1008,
N1009,N1010,N1011,N1012,N1013,N1014,N1015,N1016,N1017,N1018,
N1019,N1020,N1021,N1022,N1023,N1024,N1025,N1026,N1027,N1028,
N1029,N1030,N1031,N1032,N1033,N1034,N1035,N1036,N1037,N1038,
N1039,N1040,N1041,N1042,N1043,N1044,N1045,N1046,N1047,N1048,
N1049,N1050,N1051,N1052,N1053,N1054,N1055,N1056,N1057,N1058,
N1059,N1060,N1061,N1062,N1063,N1064,N1065,N1066,N1067,N1068,
N1069,N1070,N1071,N1072,N1073,N1074,N1075,N1076,N1077,N1078,
N1079,N1080,N1081,N1082,N1083,N1084,N1085,N1086,N1087,N1088,
N1089,N1090,N1091,N1092,N1093,N1094,N1095,N1096,N1097,N1098,
N1099,N1100,N1101,N1102,N1103,N1104,N1105,N1106,N1107,N1108,
N1109,N1110,N1111,N1112,N1113,N1114,N1115,N1116,N1117,N1118,
N1119,N1120,N1121,N1122,N1123,N1124,N1125,N1126,N1127,N1128,
N1129,N1130,N1131,N1132,N1133,N1134,N1135,N1136,N1137,N1138,
N1139,N1140,N1141,N1142,N1143,N1144,N1145,N1146,N1147,N1148,
N1149,N1150,N1151,N1152,N1153,N1154,N1155,N1156,N1157,N1158,
N1159,N1160,N1161,N1162,N1163,N1164,N1165,N1166,N1167,N1168,
N1169,N1170,N1171,N1172,N1173,N1174,N1175,N1176,N1177,N1178,
N1179,N1180,N1181,N1182,N1183,N1184,N1185,N1186,N1187,N1188,
N1189,N1190,N1191,N1192,N1193,N1194,N1195,N1196,N1197,N1198,
N1199,N1200,N1201,N1202,N1203,N1204,N1205,N1206,N1207,N1208,
N1209,N1210,N1211,N1212,N1213,N1214,N1215,N1216,N1217,N1218,
N1219,N1220,N1221,N1222,N1223,N1224,N1225,N1226,N1227,N1228,
N1229,N1230,N1231,N1232,N1233,N1234,N1235,N1236,N1237,N1238,
N1239,N1240,N1241,N1242,N1243,N1244,N1245,N1246,N1247,N1248,
N1249,N1250,N1251,N1252,N1253,N1254,N1255,N1256,N1257,N1258,
N1259,N1260,N1261,N1262,N1263,N1264,N1265,N1266,N1267,N1268,
N1269,N1270,N1271,N1272,N1273,N1274,N1275,N1276,N1277,N1278,
N1279,N1280,N1281,N1282,N1283,N1284,N1285,N1286,N1287,N1288,
N1289,N1290,N1291,N1292,N1293,N1294,N1295,N1296,N1297,N1298,
N1299,N1300,N1301,N1302,N1303,N1304,N1305,N1306,N1307,N1308,
N1309,N1310,N1311,N1312,N1313,N1314,N1315,N1316,N1317,N1318,
N1319,N1320,N1321,N1322,N1323,N1324,N1325,N1326,N1327,N1328,
N1329,N1330,N1331,N1332,N1333,N1334,N1335,N1336,N1337,N1338,
N1339,N1340,N1341,N1342,N1343,N1344,N1345,N1346,N1347,N1348,
N1349,N1350,N1351,N1352,N1353,N1354,N1355,N1356,N1357,N1358,
N1359,N1360,N1361,N1362,N1363,N1364,N1365,N1366,N1367,N1368,
N1369,N1370,N1371,N1372,N1373,N1374,N1375,N1376,N1377,N1378,
N1379,N1380,N1381,N1382,N1383,N1384,N1385,N1386,N1387,N1388,
N1389,N1390,N1391,N1392,N1393,N1394,N1395,N1396,N1397,N1398,
N1399,N1400,N1401,N1402,N1403,N1404,N1405,N1406,N1407,N1408,
N1409,N1410,N1411,N1412,N1413,N1414,N1415,N1416,N1417,N1418,
N1419,N1420,N1421,N1422,N1423,N1424,N1425,N1426,N1427,N1428,
N1429,N1430,N1431,N1432,N1433,N1434,N1435,N1436,N1437,N1438,
N1439,N1440,N1441,N1442,N1443,N1444,N1445,N1446,N1447,N1448,
N1449,N1450,N1451,N1452,N1453,N1454,N1455,N1456,N1457,N1458,
N1459,N1460,N1461,N1462,N1463,N1464,N1465,N1466,N1467,N1468,
N1469,N1470,N1471,N1472,N1473,N1474,N1475,N1476,N1477,N1478,
N1479,N1480,N1481,N1482,N1483,N1484,N1485,N1486,N1487,N1488,
N1489,N1490,N1491,N1492,N1493,N1494,N1495,N1496,N1497,N1498,
N1499,N1500,N1501,N1502,N1503,N1504,N1505,N1506,N1507,N1508,
N1509,N1510,N1511,N1512,N1513,N1514,N1515,N1516,N1517,N1518,
N1519,N1520,N1521,N1522,N1523,N1524,N1525,N1526,N1527,N1528,
N1529,N1530,N1531,N1532,N1533,N1534,N1535,N1536,N1537,N1538,
N1539,N1540,N1541,N1542,N1543,N1544,N1545,N1546,N1547,N1548,
N1549,N1550,N1551,N1552,N1553,N1554,N1555,N1556,N1557,N1558,
N1559,N1560,N1561,N1562,N1563,N1564,N1565,N1566,N1567,N1568,
N1569,N1570,N1571,N1572,N1573,N1574,N1575,N1576,N1577,N1578,
N1579,N1580,N1581,N1582,N1583,N1584,N1585,N1586,N1587,N1588,
N1589,N1590,N1591,N1592,N1593,N1594,N1595,N1596,N1597,N1598,
N1599,N1600,N1601,N1602,N1603,N1604,N1605,N1606,N1607,N1608,
N1609,N1610,N1611,N1612,N1613,N1614,N1615,N1616,N1617,N1618,
N1619,N1620,N1621,N1622,N1623,N1624,N1625,N1626,N1627,N1628,
N1629,N1630,N1631,N1632,N1633,N1634,N1635,N1636,N1637,N1638,
N1639,N1640,N1641,N1642,N1643,N1644,N1645,N1646,N1647,N1648,
N1649,N1650,N1651,N1652,N1653,N1654,N1655,N1656,N1657,N1658,
N1659,N1660,N1661,N1662,N1663,N1664,N1665,N1666,N1667,N1668,
N1669,N1670,N1671,N1672,N1673,N1674,N1675,N1676,N1677,N1678,
N1679,N1680,N1681,N1682,N1683,N1684,N1685,N1686,N1687,N1688,
N1689,N1690,N1691,N1692,N1693,N1694,N1695,N1696,N1697,N1698,
N1699,N1700,N1701,N1702,N1703,N1704,N1705,N1706,N1707,N1708,
N1709,N1710,N1711,N1712,N1713,N1714,N1715,N1716,N1717,N1718,
N1719,N1720,N1721,N1722,N1723,N1724,N1725,N1726,N1727,N1728,
N1729,N1730,N1731,N1732,N1733,N1734,N1735,N1736,N1737,N1738,
N1739,N1740,N1741,N1742,N1743,N1744,N1745,N1746,N1747,N1748,
N1749,N1750,N1751,N1752,N1753,N1754,N1755,N1756,N1757,N1758,
N1759,N1760,N1761,N1762,N1763,N1764,N1765,N1766,N1767,N1768,
N1769,N1770,N1771,N1772,N1773,N1774,N1775,N1776,N1777,N1778,
N1779,N1780,N1781,N1782,N1783,N1784,N1785,N1786,N1787,N1788,
N1789,N1790,N1791,N1792,N1793,N1794,N1795,N1796,N1797,N1798,
N1799,N1800,N1801,N1802,N1803,N1804,N1805,N1806,N1807,N1808,
N1809,N1810,N1811,N1812,N1813,N1814,N1815,N1816,N1817,N1818,
N1819,N1820,N1821,N1822,N1823,N1824,N1825,N1826,N1827,N1828,
N1829,N1830,N1831,N1832,N1833,N1834,N1835,N1836,N1837,N1838,
N1839,N1840,N1841,N1842,N1843,N1844,N1845,N1846,N1847,N1848,
N1849,N1850,N1851,N1852,N1853,N1854,N1855,N1856,N1857,N1858,
N1859,N1860,N1861,N1862,N1863,N1864,N1865,N1866,N1867,N1868,
N1869,N1870,N1871,N1872,N1873,N1874,N1875,N1876,N1877,N1878,
N1879,N1880,N1881,N1882,N1883,N1884,N1885,N1886,N1887,N1888,
N1889,N1890,N1891,N1892,N1893,N1894,N1895,N1896,N1897,N1898,
N1899,N1900,N1901,N1902,N1903,N1904,N1905,N1906,N1907,N1908,
N1909,N1910,N1911,N1912,N1913,N1914,N1915,N1916,N1917,N1918,
N1919,N1920,N1921,N1922,N1923,N1924,N1925,N1926,N1927,N1928,
N1929,N1930,N1931,N1932,N1933,N1934,N1935,N1936,N1937,N1938,
N1939,N1940,N1941,N1942,N1943,N1944,N1945,N1946,N1947,N1948,
N1949,N1950,N1951,N1952,N1953,N1954,N1955,N1956,N1957,N1958,
N1959,N1960,N1961,N1962,N1963,N1964,N1965,N1966,N1967,N1968,
N1969,N1970,N1971,N1972,N1973,N1974,N1975,N1976,N1977,N1978,
N1979,N1980,N1981,N1982,N1983,N1984,N1985,N1986,N1987,N1988,
N1989,N1990,N1991,N1992,N1993,N1994,N1995,N1996,N1997,N1998,
N1999,N2000,N2001,N2002,N2003,N2004,N2005,N2006,N2007,N2008,
N2009,N2010,N2011,N2012,N2013,N2014,N2015,N2016,N2017,N2018,
N2019,N2020,N2021,N2022,N2023,N2024,N2025,N2026,N2027,N2028,
N2029,N2030,N2031,N2032,N2033,N2034,N2035,N2036,N2037,N2038,
N2039,N2040,N2041,N2042,N2043,N2044,N2045,N2046,N2047,N2048,
N2049,N2050,N2051,N2052,N2053,N2054,N2055,N2056,N2057,N2058,
N2059,N2060,N2061,N2062,N2063,N2064,N2065,N2066,N2067,N2068,
N2069,N2070,N2071,N2072,N2073,N2074,N2075,N2076,N2077,N2078,
N2079,N2080,N2081,N2082,N2083,N2084,N2085,N2086,N2087,N2088,
N2089,N2090,N2091,N2092,N2093,N2094,N2095,N2096,N2097,N2098,
N2099,N2100,N2101,N2102,N2103,N2104,N2105,N2106,N2107,N2108,
N2109,N2110,N2111,N2112,N2113,N2114,N2115,N2116,N2117,N2118,
N2119,N2120,N2121,N2122,N2123,N2124,N2125,N2126,N2127,N2128,
N2129,N2130,N2131,N2132,N2133,N2134,N2135,N2136,N2137,N2138,
N2139,N2140,N2141,N2142,N2143,N2144,N2145,N2146,N2147,N2148,
N2149,N2150,N2151,N2152,N2153,N2154,N2155,N2156,N2157,N2158,
N2159,N2160,N2161,N2162,N2163,N2164,N2165,N2166,N2167,N2168,
N2169,N2170,N2171,N2172,N2173,N2174,N2175,N2176,N2177,N2178,
N2179,N2180,N2181,N2182,N2183,N2184,N2185,N2186,N2187,N2188,
N2189,N2190,N2191,N2192,N2193,N2194,N2195,N2196,N2197,N2198,
N2199,N2200,N2201,N2202,N2203,N2204,N2205,N2206,N2207,N2208,
N2209,N2210,N2211,N2212,N2213,N2214,N2215,N2216,N2217,N2218,
N2219,N2220,N2221,N2222,N2223,N2224,N2225,N2226,N2227,N2228,
N2229,N2230,N2231,N2232,N2233,N2234,N2235,N2236,N2237,N2238,
N2239,N2240,N2241,N2242,N2243,N2244,N2245,N2246,N2247,N2248,
N2249,N2250,N2251,N2252,N2253,N2254,N2255,N2256,N2257,N2258,
N2259,N2260,N2261,N2262,N2263,N2264,N2265,N2266,N2267,N2268,
N2269,N2270,N2271,N2272,N2273,N2274,N2275,N2276,N2277,N2278,
N2279,N2280,N2281,N2282,N2283,N2284,N2285,N2286,N2287,N2288,
N2289,N2290,N2291,N2292,N2293,N2294,N2295,N2296,N2297,N2298,
N2299,N2300,N2301,N2302,N2303,N2304,N2305,N2306,N2307,N2308,
N2309,N2310,N2311,N2312,N2313,N2314,N2315,N2316,N2317,N2318,
N2319,N2320,N2321,N2322,N2323,N2324,N2325,N2326,N2327,N2328,
N2329,N2330,N2331,N2332,N2333,N2334,N2335,N2336,N2337,N2338,
N2339,N2340,N2341,N2342,N2343,N2344,N2345,N2346,N2347,N2348,
N2349,N2350,N2351,N2352,N2353,N2354,N2355,N2356,N2357,N2358,
N2359,N2360,N2361,N2362,N2363,N2364,N2365,N2366,N2367,N2368,
N2369,N2370,N2371,N2372,N2373,N2374,N2375,N2376,N2377,N2378,
N2379,N2380,N2381,N2382,N2383,N2384,N2385,N2386,N2387,N2388,
N2389,N2390,N2391,N2392,N2393,N2394,N2395,N2396,N2397,N2398,
N2399,N2400,N2401,N2402,N2403,N2404,N2405,N2406,N2407,N2408,
N2409,N2410,N2411,N2412,N2413,N2414,N2415,N2416,N2417,N2418,
N2419,N2420,N2421,N2422,N2423,N2424,N2425,N2426,N2427,N2428,
N2429,N2430,N2431,N2432,N2433,N2434,N2435,N2436,N2437,N2438,
N2439,N2440,N2441,N2442,N2443,N2444,N2445,N2446,N2447,N2448,
N2449,N2450,N2451,N2452,N2453,N2454,N2455,N2456,N2457,N2458,
N2459,N2460,N2461,N2462,N2463,N2464,N2465,N2466,N2467,N2468,
N2469,N2470,N2471,N2472,N2473,N2474,N2475,N2476,N2477,N2478,
N2479,N2480,N2481,N2482,N2483,N2484,N2485,N2486,N2487,N2488,
N2489,N2490,N2491,N2492,N2493,N2494,N2495,N2496,N2497,N2498,
N2499,N2500,N2501,N2502,N2503,N2504,N2505,N2506,N2507,N2508,
N2509,N2510,N2511,N2512,N2513,N2514,N2515,N2516,N2517,N2518,
N2519,N2520,N2521,N2522,N2523,N2524,N2525,N2526,N2527,N2528,
N2529,N2530,N2531,N2532,N2533,N2534,N2535,N2536,N2537,N2538,
N2539,N2540,N2541,N2542,N2543,N2544,N2545,N2546,N2547,N2548,
N2549,N2550,N2551,N2552,N2553,N2554,N2555,N2556,N2557,N2558,
N2559,N2560,N2561,N2562,N2563,N2564,N2565,N2566,N2567,N2568,
N2569,N2570,N2571,N2572,N2573,N2574,N2575,N2576,N2577,N2578,
N2579,N2580,N2581,N2582,N2583,N2584,N2585,N2586,N2587,N2588,
N2589,N2590,N2591,N2592,N2593,N2594,N2595,N2596,N2597,N2598,
N2599,N2600,N2601,N2602,N2603,N2604,N2605,N2606,N2607,N2608,
N2609,N2610,N2611,N2612,N2613,N2614,N2615,N2616,N2617,N2618,
N2619,N2620,N2621,N2622,N2623,N2624,N2625,N2626,N2627,N2628,
N2629,N2630,N2631,N2632,N2633,N2634,N2635,N2636,N2637,N2638,
N2639,N2640,N2641,N2642,N2643,N2644,N2645,N2646,N2647,N2648,
N2649,N2650,N2651,N2652,N2653,N2654,N2655,N2656,N2657,N2658,
N2659,N2660,N2661,N2662,N2663,N2664,N2665,N2666,N2667,N2668,
N2669,N2670,N2671,N2672,N2673,N2674,N2675,N2676,N2677,N2678,
N2679,N2680,N2681,N2682,N2683,N2684,N2685,N2686,N2687,N2688,
N2689,N2690,N2691,N2692,N2693,N2694,N2695,N2696,N2697,N2698,
N2699,N2700,N2701,N2702,N2703,N2704,N2705,N2706,N2707,N2708,
N2709,N2710,N2711,N2712,N2713,N2714,N2715,N2716,N2717,N2718,
N2719,N2720,N2721,N2722,N2723,N2724,N2725,N2726,N2727,N2728,
N2729,N2730,N2731,N2732,N2733,N2734,N2735,N2736,N2737,N2738,
N2739,N2740,N2741,N2742,N2743,N2744,N2745,N2746,N2747,N2748,
N2749,N2750,N2751,N2752,N2753,N2754,N2755,N2756,N2757,N2758,
N2759,N2760,N2761,N2762,N2763,N2764,N2765,N2766,N2767,N2768,
N2769,N2770,N2771,N2772,N2773,N2774,N2775,N2776,N2777,N2778,
N2779,N2780,N2781,N2782,N2783,N2784,N2785,N2786,N2787,N2788,
N2789,N2790,N2791,N2792,N2793,N2794,N2795,N2796,N2797,N2798,
N2799,N2800,N2801,N2802,N2803,N2804,N2805,N2806,N2807,N2808,
N2809,N2810,N2811,N2812,N2813,N2814,N2815,N2816,N2817,N2818,
N2819,N2820,N2821,N2822,N2823,N2824,N2825,N2826,N2827,N2828,
N2829,N2830,N2831,N2832,N2833,N2834,N2835,N2836,N2837,N2838,
N2839,N2840,N2841,N2842,N2843,N2844,N2845,N2846,N2847,N2848,
N2849,N2850,N2851,N2852,N2853,N2854,N2855,N2856,N2857,N2858,
N2859,N2860,N2861,N2862,N2863,N2864,N2865,N2866,N2867,N2868,
N2869,N2870,N2871,N2872,N2873,N2874,N2875,N2876,N2877,N2878,
N2879,N2880,N2881,N2882,N2883,N2884,N2885,N2886,N2887,N2888,
N2889,N2890,N2891,N2892,N2893,N2894,N2895,N2896,N2897,N2898,
N2899,N2900,N2901,N2902,N2903,N2904,N2905,N2906,N2907,N2908,
N2909,N2910,N2911,N2912,N2913,N2914,N2915,N2916,N2917,N2918,
N2919,N2920,N2921,N2922,N2923,N2924,N2925,N2926,N2927,N2928,
N2929,N2930,N2931,N2932,N2933,N2934,N2935,N2936,N2937,N2938,
N2939,N2940,N2941,N2942,N2943,N2944,N2945,N2946,N2947,N2948,
N2949,N2950,N2951,N2952,N2953,N2954,N2955,N2956,N2957,N2958,
N2959,N2960,N2961,N2962,N2963,N2964,N2965,N2966,N2967,N2968,
N2969,N2970,N2971,N2972,N2973,N2974,N2975,N2976,N2977,N2978,
N2979,N2980,N2981,N2982,N2983,N2984,N2985,N2986,N2987,N2988,
N2989,N2990,N2991,N2992,N2993,N2994,N2995,N2996,N2997,N2998,
N2999,N3000,N3001,N3002,N3003,N3004,N3005,N3006,N3007,N3008,
N3009,N3010,N3011,N3012,N3013,N3014,N3015,N3016,N3017,N3018,
N3019,N3020,N3021,N3022,N3023,N3024,N3025,N3026,N3027,N3028,
N3029,N3030,N3031,N3032,N3033,N3034,N3035,N3036,N3037,N3038,
N3039,N3040,N3041,N3042,N3043,N3044,N3045,N3046,N3047,N3048,
N3049,N3050,N3051,N3052,N3053,N3054,N3055,N3056,N3057,N3058,
N3059,N3060,N3061,N3062,N3063,N3064,N3065,N3066,N3067,N3068,
N3069,N3070,N3071,N3072,N3073,N3074,N3075,N3076,N3077,N3078,
N3079,N3080,N3081,N3082,N3083,N3084,N3085,N3086,N3087,N3088,
N3089,N3090,N3091,N3092,N3093,N3094,N3095,N3096,N3097,N3098,
N3099,N3100,N3101,N3102,N3103,N3104,N3105,N3106,N3107,N3108,
N3109,N3110,N3111,N3112,N3113,N3114,N3115,N3116,N3117,N3118,
N3119,N3120,N3121,N3122,N3123,N3124,N3125,N3126,N3127,N3128,
N3129,N3130,N3131,N3132,N3133,N3134,N3135,N3136,N3137,N3138,
N3139,N3140,N3141,N3142,N3143,N3144,N3145,N3146,N3147,N3148,
N3149,N3150,N3151,N3152,N3153,N3154,N3155,N3156,N3157,N3158,
N3159,N3160,N3161,N3162,N3163,N3164,N3165,N3166,N3167,N3168,
N3169,N3170,N3171,N3172,N3173,N3174,N3175,N3176,N3177,N3178,
N3179,N3180,N3181,N3182,N3183,N3184,N3185,N3186,N3187,N3188,
N3189,N3190,N3191,N3192,N3193,N3194,N3195,N3196,N3197,N3198,
N3199,N3200,N3201,N3202,N3203,N3204,N3205,N3206,N3207,N3208,
N3209,N3210,N3211,N3212,N3213,N3214,N3215,N3216,N3217,N3218,
N3219,N3220,N3221,N3222,N3223,N3224,N3225,N3226,N3227,N3228,
N3229,N3230,N3231,N3232,N3233,N3234,N3235,N3236,N3237,N3238,
N3239,N3240,N3241,N3242,N3243,N3244,N3245,N3246,N3247,N3248,
N3249,N3250,N3251,N3252,N3253,N3254,N3255,N3256,N3257,N3258,
N3259,N3260,N3261,N3262,N3263,N3264,N3265,N3266,N3267,N3268,
N3269,N3270,N3271,N3272,N3273,N3274,N3275,N3276,N3277,N3278,
N3279,N3280,N3281,N3282,N3283,N3284,N3285,N3286,N3287,N3288,
N3289,N3290,N3291,N3292,N3293,N3294,N3295,N3296,N3297,N3298,
N3299,N3300,N3301,N3302,N3303,N3304,N3305,N3306,N3307,N3308,
N3309,N3310,N3311,N3312,N3313,N3314,N3315,N3316,N3317,N3318,
N3319,N3320,N3321,N3322,N3323,N3324,N3325,N3326,N3327,N3328,
N3329,N3330,N3331,N3332,N3333,N3334,N3335,N3336,N3337,N3338,
N3339,N3340,N3341,N3342,N3343,N3344,N3345,N3346,N3347,N3348,
N3349,N3350,N3351,N3352,N3353,N3354,N3355,N3356,N3357,N3358,
N3359,N3360,N3361,N3362,N3363,N3364,N3365,N3366,N3367,N3368,
N3369,N3370,N3371,N3372,N3373,N3374,N3375,N3376,N3377,N3378,
N3379,N3380,N3381,N3382,N3383,N3384,N3385,N3386,N3387,N3388,
N3389,N3390,N3391,N3392,N3393,N3394,N3395,N3396,N3397,N3398,
N3399,N3400,N3401,N3402,N3403,N3404,N3405,N3406,N3407,N3408,
N3409,N3410,N3411,N3412,N3413,N3414,N3415,N3416,N3417,N3418,
N3419,N3420,N3421,N3422,N3423,N3424,N3425,N3426,N3427,N3428,
N3429,N3430,N3431,N3432,N3433,N3434,N3435,N3436,N3437,N3438,
N3439,N3440,N3441,N3442,N3443,N3444,N3445,N3446,N3447,N3448,
N3449,N3450,N3451,N3452,N3453,N3454,N3455,N3456,N3457,N3458,
N3459,N3460,N3461,N3462,N3463,N3464,N3465,N3466,N3467,N3468,
N3469,N3470,N3471,N3472,N3473,N3474,N3475,N3476,N3477,N3478,
N3479,N3480,N3481,N3482,N3483,N3484,N3485,N3486,N3487,N3488,
N3489,N3490,N3491,N3492,N3493,N3494,N3495,N3496,N3497,N3498,
N3499,N3500,N3501,N3502,N3503,N3504,N3505,N3506,N3507,N3508,
N3509,N3510,N3511,N3512,N3513,N3514,N3515,N3516,N3517,N3518,
N3519,N3520,N3521,N3522,N3523,N3524,N3525,N3526,N3527,N3528,
N3529,N3530,N3531,N3532,N3533,N3534,N3535,N3536,N3537,N3538,
N3539,N3540,N3541,N3542,N3543,N3544,N3545,N3546,N3547,N3548,
N3549,N3550,N3551,N3552,N3553,N3554,N3555,N3556,N3557,N3558,
N3559,N3560,N3561,N3562,N3563,N3564,N3565,N3566,N3567,N3568,
N3569,N3570,N3571,N3572,N3573,N3574,N3575,N3576,N3577,N3578,
N3579,N3580,N3581,N3582,N3583,N3584,N3585,N3586,N3587,N3588,
N3589,N3590,N3591,N3592,N3593,N3594,N3595,N3596,N3597,N3598,
N3599,N3600,N3601,N3602,N3603,N3604,N3605,N3606,N3607,N3608,
N3609,N3610,N3611,N3612,N3613,N3614,N3615,N3616,N3617,N3618,
N3619,N3620,N3621,N3622,N3623,N3624,N3625,N3626,N3627,N3628,
N3629,N3630,N3631,N3632,N3633,N3634,N3635,N3636,N3637,N3638,
N3639,N3640,N3641,N3642,N3643,N3644,N3645,N3646,N3647,N3648,
N3649,N3650,N3651,N3652,N3653,N3654,N3655,N3656,N3657,N3658,
N3659,N3660,N3661,N3662,N3663,N3664,N3665,N3666,N3667,N3668,
N3669,N3670,N3671,N3672,N3673,N3674,N3675,N3676,N3677,N3678,
N3679,N3680,N3681,N3682,N3683,N3684,N3685,N3686,N3687,N3688,
N3689,N3690,N3691,N3692,N3693,N3694,N3695,N3696,N3697,N3698,
N3699,N3700,N3701,N3702,N3703,N3704,N3705,N3706,N3707,N3708,
N3709,N3710,N3711,N3712,N3713,N3714,N3715,N3716,N3717,N3718,
N3719,N3720,N3721,N3722,N3723,N3724,N3725,N3726,N3727,N3728,
N3729,N3730,N3731,N3732,N3733,N3734,N3735,N3736,N3737,N3738,
N3739,N3740,N3741,N3742,N3743,N3744,N3745,N3746,N3747,N3748,
N3749,N3750,N3751,N3752,N3753,N3754,N3755,N3756,N3757,N3758,
N3759,N3760,N3761,N3762,N3763,N3764,N3765,N3766,N3767,N3768,
N3769,N3770,N3771,N3772,N3773,N3774,N3775,N3776,N3777,N3778,
N3779,N3780,N3781,N3782,N3783,N3784,N3785,N3786,N3787,N3788,
N3789,N3790,N3791,N3792,N3793,N3794,N3795,N3796,N3797,N3798,
N3799,N3800,N3801,N3802,N3803,N3804,N3805,N3806,N3807,N3808,
N3809,N3810,N3811,N3812,N3813,N3814,N3815,N3816,N3817,N3818,
N3819,N3820,N3821,N3822,N3823,N3824,N3825,N3826,N3827,N3828,
N3829,N3830,N3831,N3832,N3833,N3834,N3835,N3836,N3837,N3838,
N3839,N3840,N3841,N3842,N3843,N3844,N3845,N3846,N3847,N3848,
N3849,N3850,N3851,N3852,N3853,N3854,N3855,N3856,N3857,N3858,
N3859,N3860,N3861,N3862,N3863,N3864,N3865,N3866,N3867,N3868,
N3869,N3870,N3871,N3872,N3873,N3874,N3875,N3876,N3877,N3878,
N3879,N3880,N3881,N3882,N3883,N3884,N3885,N3886,N3887,N3888,
N3889,N3890,N3891,N3892,N3893,N3894,N3895,N3896,N3897,N3898,
N3899,N3900,N3901,N3902,N3903,N3904,N3905,N3906,N3907,N3908,
N3909,N3910,N3911,N3912,N3913,N3914,N3915,N3916,N3917,N3918,
N3919,N3920,N3921,N3922,N3923,N3924,N3925,N3926,N3927,N3928,
N3929,N3930,N3931,N3932,N3933,N3934,N3935,N3936,N3937,N3938,
N3939,N3940,N3941,N3942,N3943,N3944,N3945,N3946,N3947,N3948,
N3949,N3950,N3951,N3952,N3953,N3954,N3955,N3956,N3957,N3958,
N3959,N3960,N3961,N3962,N3963,N3964,N3965,N3966,N3967,N3968,
N3969,N3970,N3971,N3972,N3973,N3974,N3975,N3976,N3977,N3978,
N3979,N3980,N3981,N3982,N3983,N3984,N3985,N3986,N3987,N3988,
N3989,N3990,N3991,N3992,N3993,N3994,N3995,N3996,N3997,N3998,
N3999,N4000,N4001,N4002,N4003,N4004,N4005,N4006,N4007,N4008,
N4009,N4010,N4011,N4012,N4013,N4014,N4015,N4016,N4017,N4018,
N4019,N4020,N4021,N4022,N4023,N4024,N4025,N4026,N4027,N4028,
N4029,N4030,N4031,N4032,N4033,N4034,N4035,N4036,N4037,N4038,
N4039,N4040,N4041,N4042,N4043,N4044,N4045,N4046,N4047,N4048,
N4049,N4050,N4051,N4052,N4053,N4054,N4055,N4056,N4057,N4058,
N4059,N4060,N4061,N4062,N4063,N4064,N4065,N4066,N4067,N4068,
N4069,N4070,N4071,N4072,N4073,N4074,N4075,N4076,N4077,N4078,
N4079,N4080,N4081,N4082,N4083,N4084,N4085,N4086,N4087,N4088,
N4089,N4090,N4091,N4092,N4093,N4094,N4095,N4096,N4097,N4098,
N4099,N4100,N4101,N4102,N4103,N4104,N4105,N4106,N4107,N4108,
N4109,N4110,N4111,N4112,N4113,N4114,N4115,N4116,N4117,N4118,
N4119,N4120,N4121,N4122,N4123,N4124,N4125,N4126,N4127,N4128,
N4129,N4130,N4131,N4132,N4133,N4134,N4135,N4136,N4137,N4138,
N4139,N4140,N4141,N4142,N4143,N4144,N4145,N4146,N4147,N4148,
N4149,N4150,N4151,N4152,N4153,N4154,N4155,N4156,N4157,N4158,
N4159,N4160,N4161,N4162,N4163,N4164,N4165,N4166,N4167,N4168,
N4169,N4170,N4171,N4172,N4173,N4174,N4175,N4176,N4177,N4178,
N4179,N4180,N4181,N4182,N4183,N4184,N4185,N4186,N4187,N4188,
N4189,N4190,N4191,N4192,N4193,N4194,N4195,N4196,N4197,N4198,
N4199,N4200,N4201,N4202,N4203,N4204,N4205,N4206,N4207,N4208,
N4209,N4210,N4211,N4212,N4213,N4214,N4215,N4216,N4217,N4218,
N4219,N4220,N4221,N4222,N4223,N4224,N4225,N4226,N4227,N4228,
N4229,N4230,N4231,N4232,N4233,N4234,N4235,N4236,N4237,N4238,
N4239,N4240,N4241,N4242,N4243,N4244,N4245,N4246,N4247,N4248,
N4249,N4250,N4251,N4252,N4253,N4254,N4255,N4256,N4257,N4258,
N4259,N4260,N4261,N4262,N4263,N4264,N4265,N4266,N4267,N4268,
N4269,N4270,N4271,N4272,N4273,N4274,N4275,N4276,N4277,N4278,
N4279,N4280,N4281,N4282,N4283,N4284,N4285,N4286,N4287,N4288,
N4289,N4290,N4291,N4292,N4293,N4294,N4295,N4296,N4297,N4298,
N4299,N4300,N4301,N4302,N4303,N4304,N4305,N4306,N4307,N4308,
N4309,N4310,N4311,N4312,N4313,N4314,N4315,N4316,N4317,N4318,
N4319,N4320,N4321,N4322,N4323,N4324,N4325,N4326,N4327,N4328,
N4329,N4330,N4331,N4332,N4333,N4334,N4335,N4336,N4337,N4338,
N4339,N4340,N4341,N4342,N4343,N4344,N4345,N4346,N4347,N4348,
N4349,N4350,N4351,N4352,N4353,N4354,N4355,N4356,N4357,N4358,
N4359,N4360,N4361,N4362,N4363,N4364,N4365,N4366,N4367,N4368,
N4369,N4370,N4371,N4372,N4373,N4374,N4375,N4376,N4377,N4378,
N4379,N4380,N4381,N4382,N4383,N4384,N4385,N4386,N4387,N4388,
N4389,N4390,N4391,N4392,N4393,N4394,N4395,N4396,N4397,N4398,
N4399,N4400,N4401,N4402,N4403,N4404,N4405,N4406,N4407,N4408,
N4409,N4410,N4411,N4412,N4413,N4414,N4415,N4416,N4417,N4418,
N4419,N4420,N4421,N4422,N4423,N4424,N4425,N4426,N4427,N4428,
N4429,N4430,N4431,N4432,N4433,N4434,N4435,N4436,N4437,N4438,
N4439,N4440,N4441,N4442,N4443,N4444,N4445,N4446,N4447,N4448,
N4449,N4450,N4451,N4452,N4453,N4454,N4455,N4456,N4457,N4458,
N4459,N4460,N4461,N4462,N4463,N4464,N4465,N4466,N4467,N4468,
N4469,N4470,N4471,N4472,N4473,N4474,N4475,N4476,N4477,N4478,
N4479,N4480,N4481,N4482,N4483,N4484,N4485,N4486,N4487,N4488,
N4489,N4490,N4491,N4492,N4493,N4494,N4495,N4496,N4497,N4498,
N4499,N4500,N4501,N4502,N4503,N4504,N4505,N4506,N4507,N4508,
N4509,N4510,N4511,N4512,N4513,N4514,N4515,N4516,N4517,N4518,
N4519,N4520,N4521,N4522,N4523,N4524,N4525,N4526,N4527,N4528,
N4529,N4530,N4531,N4532,N4533,N4534,N4535,N4536,N4537,N4538,
N4539,N4540,N4541,N4542,N4543,N4544,N4545,N4546,N4547,N4548,
N4549,N4550,N4551,N4552,N4553,N4554,N4555,N4556,N4557,N4558,
N4559,N4560,N4561,N4562,N4563,N4564,N4565,N4566,N4567,N4568,
N4569,N4570,N4571,N4572,N4573,N4574,N4575,N4576,N4577,N4578,
N4579,N4580,N4581,N4582,N4583,N4584,N4585,N4586,N4587,N4588,
N4589,N4590,N4591,N4592,N4593,N4594,N4595,N4596,N4597,N4598,
N4599,N4600,N4601,N4602,N4603,N4604,N4605,N4606,N4607,N4608,
N4609,N4610,N4611,N4612,N4613,N4614,N4615,N4616,N4617,N4618,
N4619,N4620,N4621,N4622,N4623,N4624,N4625,N4626,N4627,N4628,
N4629,N4630,N4631,N4632,N4633,N4634,N4635,N4636,N4637,N4638,
N4639,N4640,N4641,N4642,N4643,N4644,N4645,N4646,N4647,N4648,
N4649,N4650,N4651,N4652,N4653,N4654,N4655,N4656,N4657,N4658,
N4659,N4660,N4661,N4662,N4663,N4664,N4665,N4666,N4667,N4668,
N4669,N4670,N4671,N4672,N4673,N4674,N4675,N4676,N4677,N4678,
N4679,N4680,N4681,N4682,N4683,N4684,N4685,N4686,N4687,N4688,
N4689,N4690,N4691,N4692,N4693,N4694,N4695,N4696,N4697,N4698,
N4699,N4700,N4701,N4702,N4703,N4704,N4705,N4706,N4707,N4708,
N4709,N4710,N4711,N4712,N4713,N4714,N4715,N4716,N4717,N4718,
N4719,N4720,N4721,N4722,N4723,N4724,N4725,N4726,N4727,N4728,
N4729,N4730,N4731,N4732,N4733,N4734,N4735,N4736,N4737,N4738,
N4739,N4740,N4741,N4742,N4743,N4744,N4745,N4746,N4747,N4748,
N4749,N4750,N4751,N4752,N4753,N4754,N4755,N4756,N4757,N4758,
N4759,N4760,N4761,N4762,N4763,N4764,N4765,N4766,N4767,N4768,
N4769,N4770,N4771,N4772,N4773,N4774,N4775,N4776,N4777,N4778,
N4779,N4780,N4781,N4782,N4783,N4784,N4785,N4786,N4787,N4788,
N4789,N4790,N4791,N4792,N4793,N4794,N4795,N4796,N4797,N4798,
N4799,N4800,N4801,N4802,N4803,N4804,N4805,N4806,N4807,N4808,
N4809,N4810,N4811,N4812,N4813,N4814,N4815,N4816,N4817,N4818,
N4819,N4820,N4821,N4822,N4823,N4824,N4825,N4826,N4827,N4828,
N4829,N4830,N4831,N4832,N4833,N4834,N4835,N4836,N4837,N4838,
N4839,N4840,N4841,N4842,N4843,N4844,N4845,N4846,N4847,N4848,
N4849,N4850,N4851,N4852,N4853,N4854,N4855,N4856,N4857,N4858,
N4859,N4860,N4861,N4862,N4863,N4864,N4865,N4866,N4867,N4868,
N4869,N4870,N4871,N4872,N4873,N4874,N4875,N4876,N4877,N4878,
N4879,N4880,N4881,N4882,N4883,N4884,N4885,N4886,N4887,N4888,
N4889,N4890,N4891,N4892,N4893,N4894,N4895,N4896,N4897,N4898,
N4899,N4900,N4901,N4902,N4903,N4904,N4905,N4906,N4907,N4908,
N4909,N4910,N4911,N4912,N4913,N4914,N4915,N4916,N4917,N4918,
N4919,N4920,N4921,N4922,N4923,N4924,N4925,N4926,N4927,N4928,
N4929,N4930,N4931,N4932,N4933,N4934,N4935,N4936,N4937,N4938,
N4939,N4940,N4941,N4942,N4943,N4944,N4945,N4946,N4947,N4948,
N4949,N4950,N4951,N4952,N4953,N4954,N4955,N4956,N4957,N4958,
N4959,N4960,N4961,N4962,N4963,N4964,N4965,N4966,N4967,N4968,
N4969,N4970,N4971,N4972,N4973,N4974,N4975,N4976,N4977,N4978,
N4979,N4980,N4981,N4982,N4983,N4984,N4985,N4986,N4987,N4988,
N4989,N4990,N4991,N4992,N4993,N4994,N4995,N4996,N4997,N4998,
N4999,N5000,N5001,N5002,N5003,N5004,N5005,N5006,N5007,N5008,
N5009,N5010,N5011,N5012,N5013,N5014,N5015,N5016,N5017,N5018,
N5019,N5020,N5021,N5022,N5023,N5024,N5025,N5026,N5027,N5028,
N5029,N5030,N5031,N5032,N5033,N5034,N5035,N5036,N5037,N5038,
N5039,N5040,N5041,N5042,N5043,N5044,N5045,N5046,N5047,N5048,
N5049,N5050,N5051,N5052,N5053,N5054,N5055,N5056,N5057,N5058,
N5059,N5060,N5061,N5062,N5063,N5064,N5065,N5066,N5067,N5068,
N5069,N5070,N5071,N5072,N5073,N5074,N5075,N5076,N5077,N5078,
N5079,N5080,N5081,N5082,N5083,N5084,N5085,N5086,N5087,N5088,
N5089,N5090,N5091,N5092,N5093,N5094,N5095,N5096,N5097,N5098,
N5099,N5100,N5101,N5102,N5103,N5104,N5105,N5106,N5107,N5108,
N5109,N5110,N5111,N5112,N5113,N5114,N5115,N5116,N5117,N5118,
N5119,N5120,N5121,N5122,N5123,N5124,N5125,N5126,N5127,N5128,
N5129,N5130,N5131,N5132,N5133,N5134,N5135,N5136,N5137,N5138,
N5139,N5140,N5141,N5142,N5143,N5144,N5145,N5146,N5147,N5148,
N5149,N5150,N5151,N5152,N5153,N5154,N5155,N5156,N5157,N5158,
N5159,N5160,N5161,N5162,N5163,N5164,N5165,N5166,N5167,N5168,
N5169,N5170,N5171,N5172,N5173,N5174,N5175,N5176,N5177,N5178,
N5179,N5180,N5181,N5182,N5183,N5184,N5185,N5186,N5187,N5188,
N5189,N5190,N5191,N5192,N5193,N5194,N5195,N5196,N5197,N5198,
N5199,N5200,N5201,N5202,N5203,N5204,N5205,N5206,N5207,N5208,
N5209,N5210,N5211,N5212,N5213,N5214,N5215,N5216,N5217,N5218,
N5219,N5220,N5221,N5222,N5223,N5224,N5225,N5226,N5227,N5228,
N5229,N5230,N5231,N5232,N5233,N5234,N5235,N5236,N5237,N5238,
N5239,N5240,N5241,N5242,N5243,N5244,N5245,N5246,N5247,N5248,
N5249,N5250,N5251,N5252,N5253,N5254,N5255,N5256,N5257,N5258,
N5259,N5260,N5261,N5262,N5263,N5264,N5265,N5266,N5267,N5268,
N5269,N5270,N5271,N5272,N5273,N5274,N5275,N5276,N5277,N5278,
N5279,N5280,N5281,N5282,N5283,N5284,N5285,N5286,N5287,N5288,
N5289,N5290,N5291,N5292,N5293,N5294,N5295,N5296,N5297,N5298,
N5299,N5300,N5301,N5302,N5303,N5304,N5305,N5306,N5307,N5308,
N5309,N5310,N5311,N5312,N5313,N5314,N5315,N5316,N5317,N5318,
N5319,N5320,N5321,N5322,N5323,N5324,N5325,N5326,N5327,N5328,
N5329,N5330,N5331,N5332,N5333,N5334,N5335,N5336,N5337,N5338,
N5339,N5340,N5341,N5342,N5343,N5344,N5345,N5346,N5347,N5348,
N5349,N5350,N5351,N5352,N5353,N5354,N5355,N5356,N5357,N5358,
N5359,N5360,N5361,N5362,N5363,N5364,N5365,N5366,N5367,N5368,
N5369,N5370,N5371,N5372,N5373,N5374,N5375,N5376,N5377,N5378,
N5379,N5380,N5381,N5382,N5383,N5384,N5385,N5386,N5387,N5388,
N5389,N5390,N5391,N5392,N5393,N5394,N5395,N5396,N5397,N5398,
N5399,N5400,N5401,N5402,N5403,N5404,N5405,N5406,N5407,N5408,
N5409,N5410,N5411,N5412,N5413,N5414,N5415,N5416,N5417,N5418,
N5419,N5420,N5421,N5422,N5423,N5424,N5425,N5426,N5427,N5428,
N5429,N5430,N5431,N5432,N5433,N5434,N5435,N5436,N5437,N5438,
N5439,N5440,N5441,N5442,N5443,N5444,N5445,N5446,N5447,N5448,
N5449,N5450,N5451,N5452,N5453,N5454,N5455,N5456,N5457,N5458,
N5459,N5460,N5461,N5462,N5463,N5464,N5465,N5466,N5467,N5468,
N5469,N5470,N5471,N5472,N5473,N5474,N5475,N5476,N5477,N5478,
N5479,N5480,N5481,N5482,N5483,N5484,N5485,N5486,N5487,N5488,
N5489,N5490,N5491,N5492,N5493,N5494,N5495,N5496,N5497,N5498,
N5499,N5500,N5501,N5502,N5503,N5504,N5505,N5506,N5507,N5508,
N5509,N5510,N5511,N5512,N5513,N5514,N5515,N5516,N5517,N5518,
N5519,N5520,N5521,N5522,N5523,N5524,N5525,N5526,N5527,N5528,
N5529,N5530,N5531,N5532,N5533,N5534,N5535,N5536,N5537,N5538,
N5539,N5540,N5541,N5542,N5543,N5544,N5545,N5546,N5547,N5548,
N5549,N5550,N5551,N5552,N5553,N5554,N5555,N5556,N5557,N5558,
N5559,N5560,N5561,N5562,N5563,N5564,N5565,N5566,N5567,N5568,
N5569,N5570,N5571,N5572,N5573,N5574,N5575,N5576,N5577,N5578,
N5579,N5580,N5581,N5582,N5583,N5584,N5585,N5586,N5587,N5588,
N5589,N5590,N5591,N5592,N5593,N5594,N5595,N5596,N5597,N5598,
N5599,N5600,N5601,N5602,N5603,N5604,N5605,N5606,N5607,N5608,
N5609,N5610,N5611,N5612,N5613,N5614,N5615,N5616,N5617,N5618,
N5619,N5620,N5621,N5622,N5623,N5624,N5625,N5626,N5627,N5628,
N5629,N5630,N5631,N5632,N5633,N5634,N5635,N5636,N5637,N5638,
N5639,N5640,N5641,N5642,N5643,N5644,N5645,N5646,N5647,N5648,
N5649,N5650,N5651,N5652,N5653,N5654,N5655,N5656,N5657,N5658,
N5659,N5660,N5661,N5662,N5663,N5664,N5665,N5666,N5667,N5668,
N5669,N5670,N5671,N5672,N5673,N5674,N5675,N5676,N5677,N5678,
N5679,N5680,N5681,N5682,N5683,N5684,N5685,N5686,N5687,N5688,
N5689,N5690,N5691,N5692,N5693,N5694,N5695,N5696,N5697,N5698,
N5699,N5700,N5701,N5702,N5703,N5704,N5705,N5706,N5707,N5708,
N5709,N5710,N5711,N5712,N5713,N5714,N5715,N5716,N5717,N5718,
N5719,N5720,N5721,N5722,N5723,N5724,N5725,N5726,N5727,N5728,
N5729,N5730,N5731,N5732,N5733,N5734,N5735,N5736,N5737,N5738,
N5739,N5740,N5741,N5742,N5743,N5744,N5745,N5746,N5747,N5748,
N5749,N5750,N5751,N5752,N5753,N5754,N5755,N5756,N5757,N5758,
N5759,N5760,N5761,N5762,N5763,N5764,N5765,N5766,N5767,N5768,
N5769,N5770,N5771,N5772,N5773,N5774,N5775,N5776,N5777,N5778,
N5779,N5780,N5781,N5782,N5783,N5784,N5785,N5786,N5787,N5788,
N5789,N5790,N5791,N5792,N5793,N5794,N5795,N5796,N5797,N5798,
N5799,N5800,N5801,N5802,N5803,N5804,N5805,N5806,N5807,N5808,
N5809,N5810,N5811,N5812,N5813,N5814,N5815,N5816,N5817,N5818,
N5819,N5820,N5821,N5822,N5823,N5824,N5825,N5826,N5827,N5828,
N5829,N5830,N5831,N5832,N5833,N5834,N5835,N5836,N5837,N5838,
N5839,N5840,N5841,N5842,N5843,N5844,N5845,N5846,N5847,N5848,
N5849,N5850,N5851,N5852,N5853,N5854,N5855,N5856,N5857,N5858,
N5859,N5860,N5861,N5862,N5863,N5864,N5865,N5866,N5867,N5868,
N5869,N5870,N5871,N5872,N5873,N5874,N5875,N5876,N5877,N5878,
N5879,N5880,N5881,N5882,N5883,N5884,N5885,N5886,N5887,N5888,
N5889,N5890,N5891,N5892,N5893,N5894,N5895,N5896,N5897,N5898,
N5899,N5900,N5901,N5902,N5903,N5904,N5905,N5906,N5907,N5908,
N5909,N5910,N5911,N5912,N5913,N5914,N5915,N5916,N5917,N5918,
N5919,N5920,N5921,N5922,N5923,N5924,N5925,N5926,N5927,N5928,
N5929,N5930,N5931,N5932,N5933,N5934,N5935,N5936,N5937,N5938,
N5939,N5940,N5941,N5942,N5943,N5944,N5945,N5946,N5947,N5948,
N5949,N5950,N5951,N5952,N5953,N5954,N5955,N5956,N5957,N5958,
N5959,N5960,N5961,N5962,N5963,N5964,N5965,N5966,N5967,N5968,
N5969,N5970,N5971,N5972,N5973,N5974,N5975,N5976,N5977,N5978,
N5979,N5980,N5981,N5982,N5983,N5984,N5985,N5986,N5987,N5988,
N5989,N5990,N5991,N5992,N5993,N5994,N5995,N5996,N5997,N5998,
N5999,N6000,N6001,N6002,N6003,N6004,N6005,N6006,N6007,N6008,
N6009,N6010,N6011,N6012,N6013,N6014,N6015,N6016,N6017,N6018,
N6019,N6020,N6021,N6022,N6023,N6024,N6025,N6026,N6027,N6028,
N6029,N6030,N6031,N6032,N6033,N6034,N6035,N6036,N6037,N6038,
N6039,N6040,N6041,N6042,N6043,N6044,N6045,N6046,N6047,N6048,
N6049,N6050,N6051,N6052,N6053,N6054,N6055,N6056,N6057,N6058,
N6059,N6060,N6061,N6062,N6063,N6064,N6065,N6066,N6067,N6068,
N6069,N6070,N6071,N6072,N6073,N6074,N6075,N6076,N6077,N6078,
N6079,N6080,N6081,N6082,N6083,N6084,N6085,N6086,N6087,N6088,
N6089,N6090,N6091,N6092,N6093,N6094,N6095,N6096,N6097,N6098,
N6099,N6100,N6101,N6102,N6103,N6104,N6105,N6106,N6107,N6108,
N6109,N6110,N6111,N6112,N6113,N6114,N6115,N6116,N6117,N6118,
N6119,N6120,N6121,N6122,N6123,N6124,N6125,N6126,N6127,N6128,
N6129,N6130,N6131,N6132,N6133,N6134,N6135,N6136,N6137,N6138,
N6139,N6140,N6141,N6142,N6143,N6144,N6145,N6146,N6147,N6148,
N6149,N6150,N6151,N6152,N6153,N6154,N6155,N6156,N6157,N6158,
N6159,N6160,N6161,N6162,N6163,N6164,N6165,N6166,N6167,N6168,
N6169,N6170,N6171,N6172,N6173,N6174,N6175,N6176,N6177,N6178,
N6179,N6180,N6181,N6182,N6183,N6184,N6185,N6186,N6187,N6188,
N6189,N6190,N6191,N6192,N6193,N6194,N6195,N6196,N6197,N6198,
N6199,N6200,N6201,N6202,N6203,N6204,N6205,N6206,N6207,N6208,
N6209,N6210,N6211,N6212,N6213,N6214,N6215,N6216,N6217,N6218,
N6219,N6220,N6221,N6222,N6223,N6224,N6225,N6226,N6227,N6228,
N6229,N6230,N6231,N6232,N6233,N6234,N6235,N6236,N6237,N6238,
N6239,N6240,N6241,N6242,N6243,N6244,N6245,N6246,N6247,N6248,
N6249,N6250,N6251,N6252,N6253,N6254,N6255,N6256,N6257,N6258,
N6259,N6260,N6261,N6262,N6263,N6264,N6265,N6266,N6267,N6268,
N6269,N6270,N6271,N6272,N6273,N6274,N6275,N6276,N6277,N6278,
N6279,N6280,N6281,N6282,N6283,N6284,N6285,N6286,N6287,N6288,
N6289,N6290,N6291,N6292,N6293,N6294,N6295,N6296,N6297,N6298,
N6299,N6300,N6301,N6302,N6303,N6304,N6305,N6306,N6307,N6308,
N6309,N6310,N6311,N6312,N6313,N6314,N6315,N6316,N6317,N6318,
N6319,N6320,N6321,N6322,N6323,N6324,N6325,N6326,N6327,N6328,
N6329,N6330,N6331,N6332,N6333,N6334,N6335,N6336,N6337,N6338,
N6339,N6340,N6341,N6342,N6343,N6344,N6345,N6346,N6347,N6348,
N6349,N6350,N6351,N6352,N6353,N6354,N6355,N6356,N6357,N6358,
N6359,N6360,N6361,N6362,N6363,N6364,N6365,N6366,N6367,N6368,
N6369,N6370,N6371,N6372,N6373,N6374,N6375,N6376,N6377,N6378,
N6379,N6380,N6381,N6382,N6383,N6384,N6385,N6386,N6387,N6388,
N6389,N6390,N6391,N6392,N6393,N6394,N6395,N6396,N6397,N6398,
N6399,N6400,N6401,N6402,N6403,N6404,N6405,N6406,N6407,N6408,
N6409,N6410,N6411,N6412,N6413,N6414,N6415,N6416,N6417,N6418,
N6419,N6420,N6421,N6422,N6423,N6424,N6425,N6426,N6427,N6428,
N6429,N6430,N6431,N6432,N6433,N6434,N6435,N6436,N6437,N6438,
N6439,N6440,N6441,N6442,N6443,N6444,N6445,N6446,N6447,N6448,
N6449,N6450,N6451,N6452,N6453,N6454,N6455,N6456,N6457,N6458,
N6459,N6460,N6461,N6462,N6463,N6464,N6465,N6466,N6467,N6468,
N6469,N6470,N6471,N6472,N6473,N6474,N6475,N6476,N6477,N6478,
N6479,N6480,N6481,N6482,N6483,N6484,N6485,N6486,N6487,N6488,
N6489,N6490,N6491,N6492,N6493,N6494,N6495,N6496,N6497,N6498,
N6499,N6500,N6501,N6502,N6503,N6504,N6505,N6506,N6507,N6508,
N6509,N6510,N6511,N6512,N6513,N6514,N6515,N6516,N6517,N6518,
N6519,N6520,N6521,N6522,N6523,N6524,N6525,N6526,N6527,N6528,
N6529,N6530,N6531,N6532,N6533,N6534,N6535,N6536,N6537,N6538,
N6539,N6540,N6541,N6542,N6543,N6544,N6545,N6546,N6547,N6548,
N6549,N6550,N6551,N6552,N6553,N6554,N6555,N6556,N6557,N6558,
N6559,N6560,N6561,N6562,N6563,N6564,N6565,N6566,N6567,N6568,
N6569,N6570,N6571,N6572,N6573,N6574,N6575,N6576,N6577,N6578,
N6579,N6580,N6581,N6582,N6583,N6584,N6585,N6586,N6587,N6588,
N6589,N6590,N6591,N6592,N6593,N6594,N6595,N6596,N6597,N6598,
N6599,N6600,N6601,N6602,N6603,N6604,N6605,N6606,N6607,N6608,
N6609,N6610,N6611,N6612,N6613,N6614,N6615,N6616,N6617,N6618,
N6619,N6620,N6621,N6622,N6623,N6624,N6625,N6626,N6627,N6628,
N6629,N6630,N6631,N6632,N6633,N6634,N6635,N6636,N6637,N6638,
N6639,N6640,N6641,N6642,N6643,N6644,N6645,N6646,N6647,N6648,
N6649,N6650,N6651,N6652,N6653,N6654,N6655,N6656,N6657,N6658,
N6659,N6660,N6661,N6662,N6663,N6664,N6665,N6666,N6667,N6668,
N6669,N6670,N6671,N6672,N6673,N6674,N6675,N6676,N6677,N6678,
N6679,N6680,N6681,N6682,N6683,N6684,N6685,N6686,N6687,N6688,
N6689,N6690,N6691,N6692,N6693,N6694,N6695,N6696,N6697,N6698,
N6699,N6700,N6701,N6702,N6703,N6704,N6705,N6706,N6707,N6708,
N6709,N6710,N6711,N6712,N6713,N6714,N6715,N6716,N6717,N6718,
N6719,N6720,N6721,N6722,N6723,N6724,N6725,N6726,N6727,N6728,
N6729,N6730,N6731,N6732,N6733,N6734,N6735,N6736,N6737,N6738,
N6739,N6740,N6741,N6742,N6743,N6744,N6745,N6746,N6747,N6748,
N6749,N6750,N6751,N6752,N6753,N6754,N6755,N6756,N6757,N6758,
N6759,N6760,N6761,N6762,N6763,N6764,N6765,N6766,N6767,N6768,
N6769,N6770,N6771,N6772,N6773,N6774,N6775,N6776,N6777,N6778,
N6779,N6780,N6781,N6782,N6783,N6784,N6785,N6786,N6787,N6788,
N6789,N6790,N6791,N6792,N6793,N6794,N6795,N6796,N6797,N6798,
N6799,N6800,N6801,N6802,N6803,N6804,N6805,N6806,N6807,N6808,
N6809,N6810,N6811,N6812,N6813,N6814,N6815,N6816,N6817,N6818,
N6819,N6820,N6821,N6822,N6823,N6824,N6825,N6826,N6827,N6828,
N6829,N6830,N6831,N6832,N6833,N6834,N6835,N6836,N6837,N6838,
N6839,N6840,N6841,N6842,N6843,N6844,N6845,N6846,N6847,N6848,
N6849,N6850,N6851,N6852,N6853,N6854,N6855,N6856,N6857,N6858,
N6859,N6860,N6861,N6862,N6863,N6864,N6865,N6866,N6867,N6868,
N6869,N6870,N6871,N6872,N6873,N6874,N6875,N6876,N6877,N6878,
N6879,N6880,N6881,N6882,N6883,N6884,N6885,N6886,N6887,N6888,
N6889,N6890,N6891,N6892,N6893,N6894,N6895,N6896,N6897,N6898,
N6899,N6900,N6901,N6902,N6903,N6904,N6905,N6906,N6907,N6908,
N6909,N6910,N6911,N6912,N6913,N6914,N6915,N6916,N6917,N6918,
N6919,N6920,N6921,N6922,N6923,N6924,N6925,N6926,N6927,N6928,
N6929,N6930,N6931,N6932,N6933,N6934,N6935,N6936,N6937,N6938,
N6939,N6940,N6941,N6942,N6943,N6944,N6945,N6946,N6947,N6948,
N6949,N6950,N6951,N6952,N6953,N6954,N6955,N6956,N6957,N6958,
N6959,N6960,N6961,N6962,N6963,N6964,N6965,N6966,N6967,N6968,
N6969,N6970,N6971,N6972,N6973,N6974,N6975,N6976,N6977,N6978,
N6979,N6980,N6981,N6982,N6983,N6984,N6985,N6986,N6987,N6988,
N6989,N6990,N6991,N6992,N6993,N6994,N6995,N6996,N6997,N6998,
N6999,N7000,N7001,N7002,N7003,N7004,N7005,N7006,N7007,N7008,
N7009,N7010,N7011,N7012,N7013,N7014,N7015,N7016,N7017,N7018,
N7019,N7020,N7021,N7022,N7023,N7024,N7025,N7026,N7027,N7028,
N7029,N7030,N7031,N7032,N7033,N7034,N7035,N7036,N7037,N7038,
N7039,N7040,N7041,N7042,N7043,N7044,N7045,N7046,N7047,N7048,
N7049,N7050,N7051,N7052,N7053,N7054,N7055,N7056,N7057,N7058,
N7059,N7060,N7061,N7062,N7063,N7064,N7065,N7066,N7067,N7068,
N7069,N7070,N7071,N7072,N7073,N7074,N7075,N7076,N7077,N7078,
N7079,N7080,N7081,N7082,N7083,N7084,N7085,N7086,N7087,N7088,
N7089,N7090,N7091,N7092,N7093,N7094,N7095,N7096,N7097,N7098,
N7099,N7100,N7101,N7102,N7103,N7104,N7105,N7106,N7107,N7108,
N7109,N7110,N7111,N7112,N7113,N7114,N7115,N7116,N7117,N7118,
N7119,N7120,N7121,N7122,N7123,N7124,N7125,N7126,N7127,N7128,
N7129,N7130,N7131,N7132,N7133,N7134,N7135,N7136,N7137,N7138,
N7139,N7140,N7141,N7142,N7143,N7144,N7145,N7146,N7147,N7148,
N7149,N7150,N7151,N7152,N7153,N7154,N7155,N7156,N7157,N7158,
N7159,N7160,N7161,N7162,N7163,N7164,N7165,N7166,N7167,N7168,
N7169,N7170,N7171,N7172,N7173,N7174,N7175,N7176,N7177,N7178,
N7179,N7180,N7181,N7182,N7183,N7184,N7185,N7186,N7187,N7188,
N7189,N7190,N7191,N7192,N7193,N7194,N7195,N7196,N7197,N7198,
N7199,N7200,N7201,N7202,N7203,N7204,N7205,N7206,N7207,N7208,
N7209,N7210,N7211,N7212,N7213,N7214,N7215,N7216,N7217,N7218,
N7219,N7220,N7221,N7222,N7223,N7224,N7225,N7226,N7227,N7228,
N7229,N7230,N7231,N7232,N7233,N7234,N7235,N7236,N7237,N7238,
N7239,N7240,N7241,N7242,N7243,N7244,N7245,N7246,N7247,N7248,
N7249,N7250,N7251,N7252,N7253,N7254,N7255,N7256,N7257,N7258,
N7259,N7260,N7261,N7262,N7263,N7264,N7265,N7266,N7267,N7268,
N7269,N7270,N7271,N7272,N7273,N7274,N7275,N7276,N7277,N7278,
N7279,N7280,N7281,N7282,N7283,N7284,N7285,N7286,N7287,N7288,
N7289,N7290,N7291,N7292,N7293,N7294,N7295,N7296,N7297,N7298,
N7299,N7300,N7301,N7302,N7303,N7304,N7305,N7306,N7307,N7308,
N7309,N7310,N7311,N7312,N7313,N7314,N7315,N7316,N7317,N7318,
N7319,N7320,N7321,N7322,N7323,N7324,N7325,N7326,N7327,N7328,
N7329,N7330,N7331,N7332,N7333,N7334,N7335,N7336,N7337,N7338,
N7339,N7340,N7341,N7342,N7343,N7344,N7345,N7346,N7347,N7348,
N7349,N7350,N7351,N7352,N7353,N7354,N7355,N7356,N7357,N7358,
N7359,N7360,N7361,N7362,N7363,N7364,N7365,N7366,N7367,N7368,
N7369,N7370,N7371,N7372,N7373,N7374,N7375,N7376,N7377,N7378,
N7379,N7380,N7381,N7382,N7383,N7384,N7385,N7386,N7387,N7388,
N7389,N7390,N7391,N7392,N7393,N7394,N7395,N7396,N7397,N7398,
N7399,N7400,N7401,N7402,N7403,N7404,N7405,N7406,N7407,N7408,
N7409,N7410,N7411,N7412,N7413,N7414,N7415,N7416,N7417,N7418,
N7419,N7420,N7421,N7422,N7423,N7424,N7425,N7426,N7427,N7428,
N7429,N7430,N7431,N7432,N7433,N7434,N7435,N7436,N7437,N7438,
N7439,N7440,N7441,N7442,N7443,N7444,N7445,N7446,N7447,N7448,
N7449,N7450,N7451,N7452,N7453,N7454,N7455,N7456,N7457,N7458,
N7459,N7460,N7461,N7462,N7463,N7464,N7465,N7466,N7467,N7468,
N7469,N7470,N7471,N7472,N7473,N7474,N7475,N7476,N7477,N7478,
N7479,N7480,N7481,N7482,N7483,N7484,N7485,N7486,N7487,N7488,
N7489,N7490,N7491,N7492,N7493,N7494,N7495,N7496,N7497,N7498,
N7499,N7500,N7501,N7502,N7503,N7504,N7505,N7506,N7507,N7508,
N7509,N7510,N7511,N7512,N7513,N7514,N7515,N7516,N7517,N7518,
N7519,N7520,N7521,N7522,N7523,N7524,N7525,N7526,N7527,N7528,
N7529,N7530,N7531,N7532,N7533,N7534,N7535,N7536,N7537,N7538,
N7539,N7540,N7541,N7542,N7543,N7544,N7545,N7546,N7547,N7548,
N7549,N7550,N7551,N7552,N7553,N7554,N7555,N7556,N7557,N7558,
N7559,N7560,N7561,N7562,N7563,N7564,N7565,N7566,N7567,N7568,
N7569,N7570,N7571,N7572,N7573,N7574,N7575,N7576,N7577,N7578,
N7579,N7580,N7581,N7582,N7583,N7584,N7585,N7586,N7587,N7588,
N7589,N7590,N7591,N7592,N7593,N7594,N7595,N7596,N7597,N7598,
N7599,N7600,N7601,N7602,N7603,N7604,N7605,N7606,N7607,N7608,
N7609,N7610,N7611,N7612,N7613,N7614,N7615,N7616,N7617,N7618,
N7619,N7620,N7621,N7622,N7623,N7624,N7625,N7626,N7627,N7628,
N7629,N7630,N7631,N7632,N7633,N7634,N7635,N7636,N7637,N7638,
N7639,N7640,N7641,N7642,N7643,N7644,N7645,N7646,N7647,N7648,
N7649,N7650,N7651,N7652,N7653,N7654,N7655,N7656,N7657,N7658,
N7659,N7660,N7661,N7662,N7663,N7664,N7665,N7666,N7667,N7668,
N7669,N7670,N7671,N7672,N7673,N7674,N7675,N7676,N7677,N7678,
N7679,N7680,N7681,N7682,N7683,N7684,N7685,N7686,N7687,N7688,
N7689,N7690,N7691,N7692,N7693,N7694,N7695,N7696,N7697,N7698,
N7699,N7700,N7701,N7702,N7703,N7704,N7705,N7706,N7707,N7708,
N7709,N7710,N7711,N7712,N7713,N7714,N7715,N7716,N7717,N7718,
N7719,N7720,N7721,N7722,N7723,N7724,N7725,N7726,N7727,N7728,
N7729,N7730,N7731,N7732,N7733,N7734,N7735,N7736,N7737,N7738,
N7739,N7740,N7741,N7742,N7743,N7744,N7745,N7746,N7747,N7748,
N7749,N7750,N7751,N7752,N7753,N7754,N7755,N7756,N7757,N7758,
N7759,N7760,N7761,N7762,N7763,N7764,N7765,N7766,N7767,N7768,
N7769,N7770,N7771,N7772,N7773,N7774,N7775,N7776,N7777,N7778,
N7779,N7780,N7781,N7782,N7783,N7784,N7785,N7786,N7787,N7788,
N7789,N7790,N7791,N7792,N7793,N7794,N7795,N7796,N7797,N7798,
N7799,N7800,N7801,N7802,N7803,N7804,N7805,N7806,N7807,N7808,
N7809,N7810,N7811,N7812,N7813,N7814,N7815,N7816,N7817,N7818,
N7819,N7820,N7821,N7822,N7823,N7824,N7825,N7826,N7827,N7828,
N7829,N7830,N7831,N7832,N7833,N7834,N7835,N7836,N7837,N7838,
N7839,N7840,N7841,N7842,N7843,N7844,N7845,N7846,N7847,N7848,
N7849,N7850,N7851,N7852,N7853,N7854,N7855,N7856,N7857,N7858,
N7859,N7860,N7861,N7862,N7863,N7864,N7865,N7866,N7867,N7868,
N7869,N7870,N7871,N7872,N7873,N7874,N7875,N7876,N7877,N7878,
N7879,N7880,N7881,N7882,N7883,N7884,N7885,N7886,N7887,N7888,
N7889,N7890,N7891,N7892,N7893,N7894,N7895,N7896,N7897,N7898,
N7899,N7900,N7901,N7902,N7903,N7904,N7905,N7906,N7907,N7908,
N7909,N7910,N7911,N7912,N7913,N7914,N7915,N7916,N7917,N7918,
N7919,N7920,N7921,N7922,N7923,N7924,N7925,N7926,N7927,N7928,
N7929,N7930,N7931,N7932,N7933,N7934,N7935,N7936,N7937,N7938,
N7939,N7940,N7941,N7942,N7943,N7944,N7945,N7946,N7947,N7948,
N7949,N7950,N7951,N7952,N7953,N7954,N7955,N7956,N7957,N7958,
N7959,N7960,N7961,N7962,N7963,N7964,N7965,N7966,N7967,N7968,
N7969,N7970,N7971,N7972,N7973,N7974,N7975,N7976,N7977,N7978,
N7979,N7980,N7981,N7982,N7983,N7984,N7985,N7986,N7987,N7988,
N7989,N7990,N7991,N7992,N7993,N7994,N7995,N7996,N7997,N7998,
N7999,N8000,N8001,N8002,N8003,N8004,N8005,N8006,N8007,N8008,
N8009,N8010,N8011,N8012,N8013,N8014,N8015,N8016,N8017,N8018,
N8019,N8020,N8021,N8022,N8023,N8024,N8025,N8026,N8027,N8028,
N8029,N8030,N8031,N8032,N8033,N8034,N8035,N8036,N8037,N8038,
N8039,N8040,N8041,N8042,N8043,N8044,N8045,N8046,N8047,N8048,
N8049,N8050,N8051,N8052,N8053,N8054,N8055,N8056,N8057,N8058,
N8059,N8060,N8061,N8062,N8063,N8064,N8065,N8066,N8067,N8068,
N8069,N8070,N8071,N8072,N8073,N8074,N8075,N8076,N8077,N8078,
N8079,N8080,N8081,N8082,N8083,N8084,N8085,N8086,N8087,N8088,
N8089,N8090,N8091,N8092,N8093,N8094,N8095,N8096,N8097,N8098,
N8099,N8100,N8101,N8102,N8103,N8104,N8105,N8106,N8107,N8108,
N8109,N8110,N8111,N8112,N8113,N8114,N8115,N8116,N8117,N8118,
N8119,N8120,N8121,N8122,N8123,N8124,N8125,N8126,N8127,N8128,
N8129,N8130,N8131,N8132,N8133,N8134,N8135,N8136,N8137,N8138,
N8139,N8140,N8141,N8142,N8143,N8144,N8145,N8146,N8147,N8148,
N8149,N8150,N8151,N8152,N8153,N8154,N8155,N8156,N8157,N8158,
N8159,N8160,N8161,N8162,N8163,N8164,N8165,N8166,N8167,N8168,
N8169,N8170,N8171,N8172,N8173,N8174,N8175,N8176,N8177,N8178,
N8179,N8180,N8181,N8182,N8183,N8184,N8185,N8186,N8187,N8188,
N8189,N8190,N8191,N8192,N8193,N8194,N8195,N8196,N8197,N8198,
N8199,N8200,N8201,N8202,N8203,N8204,N8205,N8206,N8207,N8208,
N8209,N8210,N8211,N8212,N8213,N8214,N8215,N8216,N8217,N8218,
N8219,N8220,N8221,N8222,N8223,N8224,N8225,N8226,N8227,N8228,
N8229,N8230,N8231,N8232,N8233,N8234,N8235,N8236,N8237,N8238,
N8239,N8240,N8241,N8242,N8243,N8244,N8245,N8246,N8247,N8248,
N8249,N8250,N8251,N8252,N8253,N8254,N8255,N8256,N8257,N8258,
N8259,N8260,N8261,N8262,N8263,N8264,N8265,N8266,N8267,N8268,
N8269,N8270,N8271,N8272,N8273,N8274,N8275,N8276,N8277,N8278,
N8279,N8280,N8281,N8282,N8283,N8284,N8285,N8286,N8287,N8288,
N8289,N8290,N8291,N8292,N8293,N8294,N8295,N8296,N8297,N8298,
N8299,N8300,N8301,N8302,N8303,N8304,N8305,N8306,N8307,N8308,
N8309,N8310,N8311,N8312,N8313,N8314,N8315,N8316,N8317,N8318,
N8319,N8320,N8321,N8322,N8323,N8324,N8325,N8326,N8327,N8328,
N8329,N8330,N8331,N8332,N8333,N8334,N8335,N8336,N8337,N8338,
N8339,N8340,N8341,N8342,N8343,N8344,N8345,N8346,N8347,N8348,
N8349,N8350,N8351,N8352,N8353,N8354,N8355,N8356,N8357,N8358,
N8359,N8360,N8361,N8362,N8363,N8364,N8365,N8366,N8367,N8368,
N8369,N8370,N8371,N8372,N8373,N8374,N8375,N8376,N8377,N8378,
N8379,N8380,N8381,N8382,N8383,N8384,N8385,N8386,N8387,N8388,
N8389,N8390,N8391,N8392,N8393,N8394,N8395,N8396,N8397,N8398,
N8399,N8400,N8401,N8402,N8403,N8404,N8405,N8406,N8407,N8408,
N8409,N8410,N8411,N8412,N8413,N8414,N8415,N8416,N8417,N8418,
N8419,N8420,N8421,N8422,N8423,N8424,N8425,N8426,N8427,N8428,
N8429,N8430,N8431,N8432,N8433,N8434,N8435,N8436,N8437,N8438,
N8439,N8440,N8441,N8442,N8443,N8444,N8445,N8446,N8447,N8448,
N8449,N8450,N8451,N8452,N8453,N8454,N8455,N8456,N8457,N8458,
N8459,N8460,N8461,N8462,N8463,N8464,N8465,N8466,N8467,N8468,
N8469,N8470,N8471,N8472,N8473,N8474,N8475,N8476,N8477,N8478,
N8479,N8480,N8481,N8482,N8483,N8484,N8485,N8486,N8487,N8488,
N8489,N8490,N8491,N8492,N8493,N8494,N8495,N8496,N8497,N8498,
N8499,N8500,N8501,N8502,N8503,N8504,N8505,N8506,N8507,N8508,
N8509,N8510,N8511,N8512,N8513,N8514,N8515,N8516,N8517,N8518,
N8519,N8520,N8521,N8522,N8523,N8524,N8525,N8526,N8527,N8528,
N8529,N8530,N8531,N8532,N8533,N8534,N8535,N8536,N8537,N8538,
N8539,N8540,N8541,N8542,N8543,N8544,N8545,N8546,N8547,N8548,
N8549,N8550,N8551,N8552,N8553,N8554,N8555,N8556,N8557,N8558,
N8559,N8560,N8561,N8562,N8563,N8564,N8565,N8566,N8567,N8568,
N8569,N8570,N8571,N8572,N8573,N8574,N8575,N8576,N8577,N8578,
N8579,N8580,N8581,N8582,N8583,N8584,N8585,N8586,N8587,N8588,
N8589,N8590,N8591,N8592,N8593,N8594,N8595,N8596,N8597,N8598,
N8599,N8600,N8601,N8602,N8603,N8604,N8605,N8606,N8607,N8608,
N8609,N8610,N8611,N8612,N8613,N8614,N8615,N8616,N8617,N8618,
N8619,N8620,N8621,N8622,N8623,N8624,N8625,N8626,N8627,N8628,
N8629,N8630,N8631,N8632,N8633,N8634,N8635,N8636,N8637,N8638,
N8639,N8640,N8641,N8642,N8643,N8644,N8645,N8646,N8647,N8648,
N8649,N8650,N8651,N8652,N8653,N8654,N8655,N8656,N8657,N8658,
N8659,N8660,N8661,N8662,N8663,N8664,N8665,N8666,N8667,N8668,
N8669,N8670,N8671,N8672,N8673,N8674,N8675,N8676,N8677,N8678,
N8679,N8680,N8681,N8682,N8683,N8684,N8685,N8686,N8687,N8688,
N8689,N8690,N8691,N8692,N8693,N8694,N8695,N8696,N8697,N8698,
N8699,N8700,N8701,N8702,N8703,N8704,N8705,N8706,N8707,N8708,
N8709,N8710,N8711,N8712,N8713,N8714,N8715,N8716,N8717,N8718,
N8719,N8720,N8721,N8722,N8723,N8724,N8725,N8726,N8727,N8728,
N8729,N8730,N8731,N8732,N8733,N8734,N8735,N8736,N8737,N8738,
N8739,N8740,N8741,N8742,N8743,N8744,N8745,N8746,N8747,N8748,
N8749,N8750,N8751,N8752,N8753,N8754,N8755,N8756,N8757,N8758,
N8759,N8760,N8761,N8762,N8763,N8764,N8765,N8766,N8767,N8768,
N8769,N8770,N8771,N8772,N8773,N8774,N8775,N8776,N8777,N8778,
N8779,N8780,N8781,N8782,N8783,N8784,N8785,N8786,N8787,N8788,
N8789,N8790,N8791,N8792,N8793,N8794,N8795,N8796,N8797,N8798,
N8799,N8800,N8801,N8802,N8803,N8804,N8805,N8806,N8807,N8808,
N8809,N8810,N8811,N8812,N8813,N8814,N8815,N8816,N8817,N8818,
N8819,N8820,N8821,N8822,N8823,N8824,N8825,N8826,N8827,N8828,
N8829,N8830,N8831,N8832,N8833,N8834,N8835,N8836,N8837,N8838,
N8839,N8840,N8841,N8842,N8843,N8844,N8845,N8846,N8847,N8848,
N8849,N8850,N8851,N8852,N8853,N8854,N8855,N8856,N8857,N8858,
N8859,N8860,N8861,N8862,N8863,N8864,N8865,N8866,N8867,N8868,
N8869,N8870,N8871,N8872,N8873,N8874,N8875,N8876,N8877,N8878,
N8879,N8880,N8881,N8882,N8883,N8884,N8885,N8886,N8887,N8888,
N8889,N8890,N8891,N8892,N8893,N8894,N8895,N8896,N8897,N8898,
N8899,N8900,N8901,N8902,N8903,N8904,N8905,N8906,N8907,N8908,
N8909,N8910,N8911,N8912,N8913,N8914,N8915,N8916,N8917,N8918,
N8919,N8920,N8921,N8922,N8923,N8924,N8925,N8926,N8927,N8928,
N8929,N8930,N8931,N8932,N8933,N8934,N8935,N8936,N8937,N8938,
N8939,N8940,N8941,N8942,N8943,N8944,N8945,N8946,N8947,N8948,
N8949,N8950,N8951,N8952,N8953,N8954,N8955,N8956,N8957,N8958,
N8959,N8960,N8961,N8962,N8963,N8964,N8965,N8966,N8967,N8968,
N8969,N8970,N8971,N8972,N8973,N8974,N8975,N8976,N8977,N8978,
N8979,N8980,N8981,N8982,N8983,N8984,N8985,N8986,N8987,N8988,
N8989,N8990,N8991,N8992,N8993,N8994,N8995,N8996,N8997,N8998,
N8999,N9000,N9001,N9002,N9003,N9004,N9005,N9006,N9007,N9008,
N9009,N9010,N9011,N9012,N9013,N9014,N9015,N9016,N9017,N9018,
N9019,N9020,N9021,N9022,N9023,N9024,N9025,N9026,N9027,N9028,
N9029,N9030,N9031,N9032,N9033,N9034,N9035,N9036,N9037,N9038,
N9039,N9040,N9041,N9042,N9043,N9044,N9045,N9046,N9047,N9048,
N9049,N9050,N9051,N9052,N9053,N9054,N9055,N9056,N9057,N9058,
N9059,N9060,N9061,N9062,N9063,N9064,N9065,N9066,N9067,N9068,
N9069,N9070,N9071,N9072,N9073,N9074,N9075,N9076,N9077,N9078,
N9079,N9080,N9081,N9082,N9083,N9084,N9085,N9086,N9087,N9088,
N9089,N9090,N9091,N9092,N9093,N9094,N9095,N9096,N9097,N9098,
N9099,N9100,N9101,N9102,N9103,N9104,N9105,N9106,N9107,N9108,
N9109,N9110,N9111,N9112,N9113,N9114,N9115,N9116,N9117,N9118,
N9119,N9120,N9121,N9122,N9123,N9124,N9125,N9126,N9127,N9128,
N9129,N9130,N9131,N9132,N9133,N9134,N9135,N9136,N9137,N9138,
N9139,N9140,N9141,N9142,N9143,N9144,N9145,N9146,N9147,N9148,
N9149,N9150,N9151,N9152,N9153,N9154,N9155,N9156,N9157,N9158,
N9159,N9160,N9161,N9162,N9163,N9164,N9165,N9166,N9167,N9168,
N9169,N9170,N9171,N9172,N9173,N9174,N9175,N9176,N9177,N9178,
N9179,N9180,N9181,N9182,N9183,N9184,N9185,N9186,N9187,N9188,
N9189,N9190,N9191,N9192,N9193,N9194,N9195,N9196,N9197,N9198,
N9199,N9200,N9201,N9202,N9203,N9204,N9205,N9206,N9207,N9208,
N9209,N9210,N9211,N9212,N9213,N9214,N9215,N9216,N9217,N9218,
N9219,N9220,N9221,N9222,N9223,N9224,N9225,N9226,N9227,N9228,
N9229,N9230,N9231,N9232,N9233,N9234,N9235,N9236,N9237,N9238,
N9239,N9240,N9241,N9242,N9243,N9244,N9245,N9246,N9247,N9248,
N9249,N9250,N9251,N9252,N9253,N9254,N9255,N9256,N9257,N9258,
N9259,N9260,N9261,N9262,N9263,N9264,N9265,N9266,N9267,N9268,
N9269,N9270,N9271,N9272,N9273,N9274,N9275,N9276,N9277,N9278,
N9279,N9280,N9281,N9282,N9283,N9284,N9285,N9286,N9287,N9288,
N9289,N9290,N9291,N9292,N9293,N9294,N9295,N9296,N9297,N9298,
N9299,N9300,N9301,N9302,N9303,N9304,N9305,N9306,N9307,N9308,
N9309,N9310,N9311,N9312,N9313,N9314,N9315,N9316,N9317,N9318,
N9319,N9320,N9321,N9322,N9323,N9324,N9325,N9326,N9327,N9328,
N9329,N9330,N9331,N9332,N9333,N9334,N9335,N9336,N9337,N9338,
N9339,N9340,N9341,N9342,N9343,N9344,N9345,N9346,N9347,N9348,
N9349,N9350,N9351,N9352,N9353,N9354,N9355,N9356,N9357,N9358,
N9359,N9360,N9361,N9362,N9363,N9364,N9365,N9366,N9367,N9368,
N9369,N9370,N9371,N9372,N9373,N9374,N9375,N9376,N9377,N9378,
N9379,N9380,N9381,N9382,N9383,N9384,N9385,N9386,N9387,N9388,
N9389,N9390,N9391,N9392,N9393,N9394,N9395,N9396,N9397,N9398,
N9399,N9400,N9401,N9402,N9403,N9404,N9405,N9406,N9407,N9408,
N9409,N9410,N9411,N9412,N9413,N9414,N9415,N9416,N9417,N9418,
N9419,N9420,N9421,N9422,N9423,N9424,N9425,N9426,N9427,N9428,
N9429,N9430,N9431,N9432,N9433,N9434,N9435,N9436,N9437,N9438,
N9439,N9440,N9441,N9442,N9443,N9444,N9445,N9446,N9447,N9448,
N9449,N9450,N9451,N9452,N9453,N9454,N9455,N9456,N9457,N9458,
N9459,N9460,N9461,N9462,N9463,N9464,N9465,N9466,N9467,N9468,
N9469,N9470,N9471,N9472,N9473,N9474,N9475,N9476,N9477,N9478,
N9479,N9480,N9481,N9482,N9483,N9484,N9485,N9486,N9487,N9488,
N9489,N9490,N9491,N9492,N9493,N9494,N9495,N9496,N9497,N9498,
N9499,N9500,N9501,N9502,N9503,N9504,N9505,N9506,N9507,N9508,
N9509,N9510,N9511,N9512,N9513,N9514,N9515,N9516,N9517,N9518,
N9519,N9520,N9521,N9522,N9523,N9524,N9525,N9526,N9527,N9528,
N9529,N9530,N9531,N9532,N9533,N9534,N9535,N9536,N9537,N9538,
N9539,N9540,N9541,N9542,N9543,N9544,N9545,N9546,N9547,N9548,
N9549,N9550,N9551,N9552,N9553,N9554,N9555,N9556,N9557,N9558,
N9559,N9560,N9561,N9562,N9563,N9564,N9565,N9566,N9567,N9568,
N9569,N9570,N9571,N9572,N9573,N9574,N9575,N9576,N9577,N9578,
N9579,N9580,N9581,N9582,N9583,N9584,N9585,N9586,N9587,N9588,
N9589,N9590,N9591,N9592,N9593,N9594,N9595,N9596,N9597,N9598,
N9599,N9600,N9601,N9602,N9603,N9604,N9605,N9606,N9607,N9608,
N9609,N9610,N9611,N9612,N9613,N9614,N9615,N9616,N9617,N9618,
N9619,N9620,N9621,N9622,N9623,N9624,N9625,N9626,N9627,N9628,
N9629,N9630,N9631,N9632,N9633,N9634,N9635,N9636,N9637,N9638,
N9639,N9640,N9641,N9642,N9643,N9644,N9645,N9646,N9647,N9648,
N9649,N9650,N9651,N9652,N9653,N9654,N9655,N9656,N9657,N9658,
N9659,N9660,N9661,N9662,N9663,N9664,N9665,N9666,N9667,N9668,
N9669,N9670,N9671,N9672,N9673,N9674,N9675,N9676,N9677,N9678,
N9679,N9680,N9681,N9682,N9683,N9684,N9685,N9686,N9687,N9688,
N9689,N9690,N9691,N9692,N9693,N9694,N9695,N9696,N9697,N9698,
N9699,N9700,N9701,N9702,N9703,N9704,N9705,N9706,N9707,N9708,
N9709,N9710,N9711,N9712,N9713,N9714,N9715,N9716,N9717,N9718,
N9719,N9720,N9721,N9722,N9723,N9724,N9725,N9726,N9727,N9728,
N9729,N9730,N9731,N9732,N9733,N9734,N9735,N9736,N9737,N9738,
N9739,N9740,N9741,N9742,N9743,N9744,N9745,N9746,N9747,N9748,
N9749,N9750,N9751,N9752,N9753,N9754,N9755,N9756,N9757,N9758,
N9759,N9760,N9761,N9762,N9763,N9764,N9765,N9766,N9767,N9768,
N9769,N9770,N9771,N9772,N9773,N9774,N9775,N9776,N9777,N9778,
N9779,N9780,N9781,N9782,N9783,N9784,N9785,N9786,N9787,N9788,
N9789,N9790,N9791,N9792,N9793,N9794,N9795,N9796,N9797,N9798,
N9799,N9800,N9801,N9802,N9803,N9804,N9805,N9806,N9807,N9808,
N9809,N9810,N9811,N9812,N9813,N9814,N9815,N9816,N9817,N9818,
N9819,N9820,N9821,N9822,N9823,N9824,N9825,N9826,N9827,N9828,
N9829,N9830,N9831,N9832,N9833,N9834,N9835,N9836,N9837,N9838,
N9839,N9840,N9841,N9842,N9843,N9844,N9845,N9846,N9847,N9848,
N9849,N9850,N9851,N9852,N9853,N9854,N9855,N9856,N9857,N9858,
N9859,N9860,N9861,N9862,N9863,N9864,N9865,N9866,N9867,N9868,
N9869,N9870,N9871,N9872,N9873,N9874,N9875,N9876,N9877,N9878,
N9879,N9880,N9881,N9882,N9883,N9884,N9885,N9886,N9887,N9888,
N9889,N9890,N9891,N9892,N9893,N9894,N9895,N9896,N9897,N9898,
N9899,N9900,N9901,N9902,N9903,N9904,N9905,N9906,N9907,N9908,
N9909,N9910,N9911,N9912,N9913,N9914,N9915,N9916,N9917,N9918,
N9919,N9920,N9921,N9922,N9923,N9924,N9925,N9926,N9927,N9928,
N9929,N9930,N9931,N9932,N9933,N9934,N9935,N9936,N9937,N9938,
N9939,N9940,N9941,N9942,N9943,N9944,N9945,N9946,N9947,N9948,
N9949,N9950,N9951,N9952,N9953,N9954,N9955,N9956,N9957,N9958,
N9959,N9960,N9961,N9962,N9963,N9964,N9965,N9966,N9967,N9968,
N9969,N9970,N9971,N9972,N9973,N9974,N9975,N9976,N9977,N9978,
N9979,N9980,N9981,N9982,N9983,N9984,N9985,N9986,N9987,N9988,
N9989,N9990,N9991,N9992,N9993,N9994,N9995,N9996,N9997,N9998,
N9999,N10000,N10001,N10002,N10003,N10004,N10005,N10006,N10007,N10008,
N10009,N10010,N10011,N10012,N10013,N10014,N10015,N10016,N10017,N10018,
N10019,N10020,N10021,N10022,N10023,N10024,N10025,N10026,N10027,N10028,
N10029,N10030,N10031,N10032,N10033,N10034,N10035,N10036,N10037,N10038,
N10039,N10040,N10041,N10042,N10043,N10044,N10045,N10046,N10047,N10048,
N10049,N10050,N10051,N10052,N10053,N10054,N10055,N10056,N10057,N10058,
N10059,N10060,N10061,N10062,N10063,N10064,N10065,N10066,N10067,N10068,
N10069,N10070,N10071,N10072,N10073,N10074,N10075,N10076,N10077,N10078,
N10079,N10080,N10081,N10082,N10083,N10084,N10085,N10086,N10087,N10088,
N10089,N10090,N10091,N10092,N10093,N10094,N10095,N10096,N10097,N10098,
N10099,N10100,N10101,N10102,N10103,N10104,N10105,N10106,N10107,N10108,
N10109,N10110,N10111,N10112,N10113,N10114,N10115,N10116,N10117,N10118,
N10119,N10120,N10121,N10122,N10123,N10124,N10125,N10126,N10127,N10128,
N10129,N10130,N10131,N10132,N10133,N10134,N10135,N10136,N10137,N10138,
N10139,N10140,N10141,N10142,N10143,N10144,N10145,N10146,N10147,N10148,
N10149,N10150,N10151,N10152,N10153,N10154,N10155,N10156,N10157,N10158,
N10159,N10160,N10161,N10162,N10163,N10164,N10165,N10166,N10167,N10168,
N10169,N10170,N10171,N10172,N10173,N10174,N10175,N10176,N10177,N10178,
N10179,N10180,N10181,N10182,N10183,N10184,N10185,N10186,N10187,N10188,
N10189,N10190,N10191,N10192,N10193,N10194,N10195,N10196,N10197,N10198,
N10199,N10200,N10201,N10202,N10203,N10204,N10205,N10206,N10207,N10208,
N10209,N10210,N10211,N10212,N10213,N10214,N10215,N10216,N10217,N10218,
N10219,N10220,N10221,N10222,N10223,N10224,N10225,N10226,N10227,N10228,
N10229,N10230,N10231,N10232,N10233,N10234,N10235,N10236,N10237,N10238,
N10239,N10240,N10241,N10242,N10243,N10244,N10245,N10246,N10247,N10248,
N10249,N10250,N10251,N10252,N10253,N10254,N10255,N10256,N10257,N10258,
N10259,N10260,N10261,N10262,N10263,N10264,N10265,N10266,N10267,N10268,
N10269,N10270,N10271,N10272,N10273,N10274,N10275,N10276,N10277,N10278,
N10279,N10280,N10281,N10282,N10283,N10284,N10285,N10286,N10287,N10288,
N10289,N10290,N10291,N10292,N10293,N10294,N10295,N10296,N10297,N10298,
N10299,N10300,N10301,N10302,N10303,N10304,N10305,N10306,N10307,N10308,
N10309,N10310,N10311,N10312,N10313,N10314,N10315,N10316,N10317,N10318,
N10319,N10320,N10321,N10322,N10323,N10324,N10325,N10326,N10327,N10328,
N10329,N10330,N10331,N10332,N10333,N10334,N10335,N10336,N10337,N10338,
N10339,N10340,N10341,N10342,N10343,N10344,N10345,N10346,N10347,N10348,
N10349,N10350,N10351,N10352,N10353,N10354,N10355,N10356,N10357,N10358,
N10359,N10360,N10361,N10362,N10363,N10364,N10365,N10366,N10367,N10368,
N10369,N10370,N10371,N10372,N10373,N10374,N10375,N10376,N10377,N10378,
N10379,N10380,N10381,N10382,N10383,N10384,N10385,N10386,N10387,N10388,
N10389,N10390,N10391,N10392,N10393,N10394,N10395,N10396,N10397,N10398,
N10399,N10400,N10401,N10402,N10403,N10404,N10405,N10406,N10407,N10408,
N10409,N10410,N10411,N10412,N10413,N10414,N10415,N10416,N10417,N10418,
N10419,N10420,N10421,N10422,N10423,N10424,N10425,N10426,N10427,N10428,
N10429,N10430,N10431,N10432,N10433,N10434,N10435,N10436,N10437,N10438,
N10439,N10440,N10441,N10442,N10443,N10444,N10445,N10446,N10447,N10448,
N10449,N10450,N10451,N10452,N10453,N10454,N10455,N10456,N10457,N10458,
N10459,N10460,N10461,N10462,N10463,N10464,N10465,N10466,N10467,N10468,
N10469,N10470,N10471,N10472,N10473,N10474,N10475,N10476,N10477,N10478,
N10479,N10480,N10481,N10482,N10483,N10484,N10485,N10486,N10487,N10488,
N10489,N10490,N10491,N10492,N10493,N10494,N10495,N10496,N10497,N10498,
N10499,N10500,N10501,N10502,N10503,N10504,N10505,N10506,N10507,N10508,
N10509,N10510,N10511,N10512,N10513,N10514,N10515,N10516,N10517,N10518,
N10519,N10520,N10521,N10522,N10523,N10524,N10525,N10526,N10527,N10528,
N10529,N10530,N10531,N10532,N10533,N10534,N10535,N10536,N10537,N10538,
N10539,N10540,N10541,N10542,N10543,N10544,N10545,N10546,N10547,N10548,
N10549,N10550,N10551,N10552,N10553,N10554,N10555,N10556,N10557,N10558,
N10559,N10560,N10561,N10562,N10563,N10564,N10565,N10566,N10567,N10568,
N10569,N10570,N10571,N10572,N10573,N10574,N10575,N10576,N10577,N10578,
N10579,N10580,N10581,N10582,N10583,N10584,N10585,N10586,N10587,N10588,
N10589,N10590,N10591,N10592,N10593,N10594,N10595,N10596,N10597,N10598,
N10599,N10600,N10601,N10602,N10603,N10604,N10605,N10606,N10607,N10608,
N10609,N10610,N10611,N10612,N10613,N10614,N10615,N10616,N10617,N10618,
N10619,N10620,N10621,N10622,N10623,N10624,N10625,N10626,N10627,N10628,
N10629,N10630,N10631,N10632,N10633,N10634,N10635,N10636,N10637,N10638,
N10639,N10640,N10641,N10642,N10643,N10644,N10645,N10646,N10647,N10648,
N10649,N10650,N10651,N10652,N10653,N10654,N10655,N10656,N10657,N10658,
N10659,N10660,N10661,N10662,N10663,N10664,N10665,N10666,N10667,N10668,
N10669,N10670,N10671,N10672,N10673,N10674,N10675,N10676,N10677,N10678,
N10679,N10680,N10681,N10682,N10683,N10684,N10685,N10686,N10687,N10688,
N10689,N10690,N10691,N10692,N10693,N10694,N10695,N10696,N10697,N10698,
N10699,N10700,N10701,N10702,N10703,N10704,N10705,N10706,N10707,N10708,
N10709,N10710,N10711,N10712,N10713,N10714,N10715,N10716,N10717,N10718,
N10719,N10720,N10721,N10722,N10723,N10724,N10725,N10726,N10727,N10728,
N10729,N10730,N10731,N10732,N10733,N10734,N10735,N10736,N10737,N10738,
N10739,N10740,N10741,N10742,N10743,N10744,N10745,N10746,N10747,N10748,
N10749,N10750,N10751,N10752,N10753,N10754,N10755,N10756,N10757,N10758,
N10759,N10760,N10761,N10762,N10763,N10764,N10765,N10766,N10767,N10768,
N10769,N10770,N10771,N10772,N10773,N10774,N10775,N10776,N10777,N10778,
N10779,N10780,N10781,N10782,N10783,N10784,N10785,N10786,N10787,N10788,
N10789,N10790,N10791,N10792,N10793,N10794,N10795,N10796,N10797,N10798,
N10799,N10800,N10801,N10802,N10803,N10804,N10805,N10806,N10807,N10808,
N10809,N10810,N10811,N10812,N10813,N10814,N10815,N10816,N10817,N10818,
N10819,N10820,N10821,N10822,N10823,N10824,N10825,N10826,N10827,N10828,
N10829,N10830,N10831,N10832,N10833,N10834,N10835,N10836,N10837,N10838,
N10839,N10840,N10841,N10842,N10843,N10844,N10845,N10846,N10847,N10848,
N10849,N10850,N10851,N10852,N10853,N10854,N10855,N10856,N10857,N10858,
N10859,N10860,N10861,N10862,N10863,N10864,N10865,N10866,N10867,N10868,
N10869,N10870,N10871,N10872,N10873,N10874,N10875,N10876,N10877,N10878,
N10879,N10880,N10881,N10882,N10883,N10884,N10885,N10886,N10887,N10888,
N10889,N10890,N10891,N10892,N10893,N10894,N10895,N10896,N10897,N10898,
N10899,N10900,N10901,N10902,N10903,N10904,N10905,N10906,N10907,N10908,
N10909,N10910,N10911,N10912,N10913,N10914,N10915,N10916,N10917,N10918,
N10919,N10920,N10921,N10922,N10923,N10924,N10925,N10926,N10927,N10928,
N10929,N10930,N10931,N10932,N10933,N10934,N10935,N10936,N10937,N10938,
N10939,N10940,N10941,N10942,N10943,N10944,N10945,N10946,N10947,N10948,
N10949,N10950,N10951,N10952,N10953,N10954,N10955,N10956,N10957,N10958,
N10959,N10960,N10961,N10962,N10963,N10964,N10965,N10966,N10967,N10968,
N10969,N10970,N10971,N10972,N10973,N10974,N10975,N10976,N10977,N10978,
N10979,N10980,N10981,N10982,N10983,N10984,N10985,N10986,N10987,N10988,
N10989,N10990,N10991,N10992,N10993,N10994,N10995,N10996,N10997,N10998,
N10999,N11000,N11001,N11002,N11003,N11004,N11005,N11006,N11007,N11008,
N11009,N11010,N11011,N11012,N11013,N11014,N11015,N11016,N11017,N11018,
N11019,N11020,N11021,N11022,N11023,N11024,N11025,N11026,N11027,N11028,
N11029,N11030,N11031,N11032,N11033,N11034,N11035,N11036,N11037,N11038,
N11039,N11040,N11041,N11042,N11043,N11044,N11045,N11046,N11047,N11048,
N11049,N11050,N11051,N11052,N11053,N11054,N11055,N11056,N11057,N11058,
N11059,N11060,N11061,N11062,N11063,N11064,N11065,N11066,N11067,N11068,
N11069,N11070,N11071,N11072,N11073,N11074,N11075,N11076,N11077,N11078,
N11079,N11080,N11081,N11082,N11083,N11084,N11085,N11086,N11087,N11088,
N11089,N11090,N11091,N11092,N11093,N11094,N11095,N11096,N11097,N11098,
N11099,N11100,N11101,N11102,N11103,N11104,N11105,N11106,N11107,N11108,
N11109,N11110,N11111,N11112,N11113,N11114,N11115,N11116,N11117,N11118,
N11119,N11120,N11121,N11122,N11123,N11124,N11125,N11126,N11127,N11128,
N11129,N11130,N11131,N11132,N11133,N11134,N11135,N11136,N11137,N11138,
N11139,N11140,N11141,N11142,N11143,N11144,N11145,N11146,N11147,N11148,
N11149,N11150,N11151,N11152,N11153,N11154,N11155,N11156,N11157,N11158,
N11159,N11160,N11161,N11162,N11163,N11164,N11165,N11166,N11167,N11168,
N11169,N11170,N11171,N11172,N11173,N11174,N11175,N11176,N11177,N11178,
N11179,N11180,N11181,N11182,N11183,N11184,N11185,N11186,N11187,N11188,
N11189,N11190,N11191,N11192,N11193,N11194,N11195,N11196,N11197,N11198,
N11199,N11200,N11201,N11202,N11203,N11204,N11205,N11206,N11207,N11208,
N11209,N11210,N11211,N11212,N11213,N11214,N11215,N11216,N11217,N11218,
N11219,N11220,N11221,N11222,N11223,N11224,N11225,N11226,N11227,N11228,
N11229,N11230,N11231,N11232,N11233,N11234,N11235,N11236,N11237,N11238,
N11239,N11240,N11241,N11242,N11243,N11244,N11245,N11246,N11247,N11248,
N11249,N11250,N11251,N11252,N11253,N11254,N11255,N11256,N11257,N11258,
N11259,N11260,N11261,N11262,N11263,N11264,N11265,N11266,N11267,N11268,
N11269,N11270,N11271,N11272,N11273,N11274,N11275,N11276,N11277,N11278,
N11279,N11280,N11281,N11282,N11283,N11284,N11285,N11286,N11287,N11288,
N11289,N11290,N11291,N11292,N11293,N11294,N11295,N11296,N11297,N11298,
N11299,N11300,N11301,N11302,N11303,N11304,N11305,N11306,N11307,N11308,
N11309,N11310,N11311,N11312,N11313,N11314,N11315,N11316,N11317,N11318,
N11319,N11320,N11321,N11322,N11323,N11324,N11325,N11326,N11327,N11328,
N11329,N11330,N11331,N11332,N11333,N11334,N11335,N11336,N11337,N11338,
N11339,N11340,N11341,N11342,N11343,N11344,N11345,N11346,N11347,N11348,
N11349,N11350,N11351,N11352,N11353,N11354,N11355,N11356,N11357,N11358,
N11359,N11360,N11361,N11362,N11363,N11364,N11365,N11366,N11367,N11368,
N11369,N11370,N11371,N11372,N11373,N11374,N11375,N11376,N11377,N11378,
N11379,N11380,N11381,N11382,N11383,N11384,N11385,N11386,N11387,N11388,
N11389,N11390,N11391,N11392,N11393,N11394,N11395,N11396,N11397,N11398,
N11399,N11400,N11401,N11402,N11403,N11404,N11405,N11406,N11407,N11408,
N11409,N11410,N11411,N11412,N11413,N11414,N11415,N11416,N11417,N11418,
N11419,N11420,N11421,N11422,N11423,N11424,N11425,N11426,N11427,N11428,
N11429,N11430,N11431,N11432,N11433,N11434,N11435,N11436,N11437,N11438,
N11439,N11440,N11441,N11442,N11443,N11444,N11445,N11446,N11447,N11448,
N11449,N11450,N11451,N11452,N11453,N11454,N11455,N11456,N11457,N11458,
N11459,N11460,N11461,N11462,N11463,N11464,N11465,N11466,N11467,N11468,
N11469,N11470,N11471,N11472,N11473,N11474,N11475,N11476,N11477,N11478,
N11479,N11480,N11481,N11482,N11483,N11484,N11485,N11486,N11487,N11488,
N11489,N11490,N11491,N11492,N11493,N11494,N11495,N11496,N11497,N11498,
N11499,N11500,N11501,N11502,N11503,N11504,N11505,N11506,N11507,N11508,
N11509,N11510,N11511,N11512,N11513,N11514,N11515,N11516,N11517,N11518,
N11519,N11520,N11521,N11522,N11523,N11524,N11525,N11526,N11527,N11528,
N11529,N11530,N11531,N11532,N11533,N11534,N11535,N11536,N11537,N11538,
N11539,N11540,N11541,N11542,N11543,N11544,N11545,N11546,N11547,N11548,
N11549,N11550,N11551,N11552,N11553,N11554,N11555,N11556,N11557,N11558,
N11559,N11560,N11561,N11562,N11563,N11564,N11565,N11566,N11567,N11568,
N11569,N11570,N11571,N11572,N11573,N11574,N11575,N11576,N11577,N11578,
N11579,N11580,N11581,N11582,N11583,N11584,N11585,N11586,N11587,N11588,
N11589,N11590,N11591,N11592,N11593,N11594,N11595,N11596,N11597,N11598,
N11599,N11600,N11601,N11602,N11603,N11604,N11605,N11606,N11607,N11608,
N11609,N11610,N11611,N11612,N11613,N11614,N11615,N11616,N11617,N11618,
N11619,N11620,N11621,N11622,N11623,N11624,N11625,N11626,N11627,N11628,
N11629,N11630,N11631,N11632,N11633,N11634,N11635,N11636,N11637,N11638,
N11639,N11640,N11641,N11642,N11643,N11644,N11645,N11646,N11647,N11648,
N11649,N11650,N11651,N11652,N11653,N11654,N11655,N11656,N11657,N11658,
N11659,N11660,N11661,N11662,N11663,N11664,N11665,N11666,N11667,N11668,
N11669,N11670,N11671,N11672,N11673,N11674,N11675,N11676,N11677,N11678,
N11679,N11680,N11681,N11682,N11683,N11684,N11685,N11686,N11687,N11688,
N11689,N11690,N11691,N11692,N11693,N11694,N11695,N11696,N11697,N11698,
N11699,N11700,N11701,N11702,N11703,N11704,N11705,N11706,N11707,N11708,
N11709,N11710,N11711,N11712,N11713,N11714,N11715,N11716,N11717,N11718,
N11719,N11720,N11721,N11722,N11723,N11724,N11725,N11726,N11727,N11728,
N11729,N11730,N11731,N11732,N11733,N11734,N11735,N11736,N11737,N11738,
N11739,N11740,N11741,N11742,N11743,N11744,N11745,N11746,N11747,N11748,
N11749,N11750,N11751,N11752,N11753,N11754,N11755,N11756,N11757,N11758,
N11759,N11760,N11761,N11762,N11763,N11764,N11765,N11766,N11767,N11768,
N11769,N11770,N11771,N11772,N11773,N11774,N11775,N11776,N11777,N11778,
N11779,N11780,N11781,N11782,N11783,N11784,N11785,N11786,N11787,N11788,
N11789,N11790,N11791,N11792,N11793,N11794,N11795,N11796,N11797,N11798,
N11799,N11800,N11801,N11802,N11803,N11804,N11805,N11806,N11807,N11808,
N11809,N11810,N11811,N11812,N11813,N11814,N11815,N11816,N11817,N11818,
N11819,N11820,N11821,N11822,N11823,N11824,N11825,N11826,N11827,N11828,
N11829,N11830,N11831,N11832,N11833,N11834,N11835,N11836,N11837,N11838,
N11839,N11840,N11841,N11842,N11843,N11844,N11845,N11846,N11847,N11848,
N11849,N11850,N11851,N11852,N11853,N11854,N11855,N11856,N11857,N11858,
N11859,N11860,N11861,N11862,N11863,N11864,N11865,N11866,N11867,N11868,
N11869,N11870,N11871,N11872,N11873,N11874,N11875,N11876,N11877,N11878,
N11879,N11880,N11881,N11882,N11883,N11884,N11885,N11886,N11887,N11888,
N11889,N11890,N11891,N11892,N11893,N11894,N11895,N11896,N11897,N11898,
N11899,N11900,N11901,N11902,N11903,N11904,N11905,N11906,N11907,N11908,
N11909,N11910,N11911,N11912,N11913,N11914,N11915,N11916,N11917,N11918,
N11919,N11920,N11921,N11922,N11923,N11924,N11925,N11926,N11927,N11928,
N11929,N11930,N11931,N11932,N11933,N11934,N11935,N11936,N11937,N11938,
N11939,N11940,N11941,N11942,N11943,N11944,N11945,N11946,N11947,N11948,
N11949,N11950,N11951,N11952,N11953,N11954,N11955,N11956,N11957,N11958,
N11959,N11960,N11961,N11962,N11963,N11964,N11965,N11966,N11967,N11968,
N11969,N11970,N11971,N11972,N11973,N11974,N11975,N11976,N11977,N11978,
N11979,N11980,N11981,N11982,N11983,N11984,N11985,N11986,N11987,N11988,
N11989,N11990,N11991,N11992,N11993,N11994,N11995,N11996,N11997,N11998,
N11999,N12000,N12001,N12002,N12003,N12004,N12005,N12006,N12007,N12008,
N12009,N12010,N12011,N12012,N12013,N12014,N12015,N12016,N12017,N12018,
N12019,N12020,N12021,N12022,N12023,N12024,N12025,N12026,N12027,N12028,
N12029,N12030,N12031,N12032,N12033,N12034,N12035,N12036,N12037,N12038,
N12039,N12040,N12041,N12042,N12043,N12044,N12045,N12046,N12047,N12048,
N12049,N12050,N12051,N12052,N12053,N12054,N12055,N12056,N12057,N12058,
N12059,N12060,N12061,N12062,N12063,N12064,N12065,N12066,N12067,N12068,
N12069,N12070,N12071,N12072,N12073,N12074,N12075,N12076,N12077,N12078,
N12079,N12080,N12081,N12082,N12083,N12084,N12085,N12086,N12087,N12088,
N12089,N12090,N12091,N12092,N12093,N12094,N12095,N12096,N12097,N12098,
N12099,N12100,N12101,N12102,N12103,N12104,N12105,N12106,N12107,N12108,
N12109,N12110,N12111,N12112,N12113,N12114,N12115,N12116,N12117,N12118,
N12119,N12120,N12121,N12122,N12123,N12124,N12125,N12126,N12127,N12128,
N12129,N12130,N12131,N12132,N12133,N12134,N12135,N12136,N12137,N12138,
N12139,N12140,N12141,N12142,N12143,N12144,N12145,N12146,N12147,N12148,
N12149,N12150,N12151,N12152,N12153,N12154,N12155,N12156,N12157,N12158,
N12159,N12160,N12161,N12162,N12163,N12164,N12165,N12166,N12167,N12168,
N12169,N12170,N12171,N12172,N12173,N12174,N12175,N12176,N12177,N12178,
N12179,N12180,N12181,N12182,N12183,N12184,N12185,N12186,N12187,N12188,
N12189,N12190,N12191,N12192,N12193,N12194,N12195,N12196,N12197,N12198,
N12199,N12200,N12201,N12202,N12203,N12204,N12205,N12206,N12207,N12208,
N12209,N12210,N12211,N12212,N12213,N12214,N12215,N12216,N12217,N12218,
N12219,N12220,N12221,N12222,N12223,N12224,N12225,N12226,N12227,N12228,
N12229,N12230,N12231,N12232,N12233,N12234,N12235,N12236,N12237,N12238,
N12239,N12240,N12241,N12242,N12243,N12244,N12245,N12246,N12247,N12248,
N12249,N12250,N12251,N12252,N12253,N12254,N12255,N12256,N12257,N12258,
N12259,N12260,N12261,N12262,N12263,N12264,N12265,N12266,N12267,N12268,
N12269,N12270,N12271,N12272,N12273,N12274,N12275,N12276,N12277,N12278,
N12279,N12280,N12281,N12282,N12283,N12284,N12285,N12286,N12287,N12288,
N12289,N12290,N12291,N12292,N12293,N12294,N12295,N12296,N12297,N12298,
N12299,N12300,N12301,N12302,N12303,N12304,N12305,N12306,N12307,N12308,
N12309,N12310,N12311,N12312,N12313,N12314,N12315,N12316,N12317,N12318,
N12319,N12320,N12321,N12322,N12323,N12324,N12325,N12326,N12327,N12328,
N12329,N12330,N12331,N12332,N12333,N12334,N12335,N12336,N12337,N12338,
N12339,N12340,N12341,N12342,N12343,N12344,N12345,N12346,N12347,N12348,
N12349,N12350,N12351,N12352,N12353,N12354,N12355,N12356,N12357,N12358,
N12359,N12360,N12361,N12362,N12363,N12364,N12365,N12366,N12367,N12368,
N12369,N12370,N12371,N12372,N12373,N12374,N12375,N12376,N12377,N12378,
N12379,N12380,N12381,N12382,N12383,N12384,N12385,N12386,N12387,N12388,
N12389,N12390,N12391,N12392,N12393,N12394,N12395,N12396,N12397,N12398,
N12399,N12400,N12401,N12402,N12403,N12404,N12405,N12406,N12407,N12408,
N12409,N12410,N12411,N12412,N12413,N12414,N12415,N12416,N12417,N12418,
N12419,N12420,N12421,N12422,N12423,N12424,N12425,N12426,N12427,N12428,
N12429,N12430,N12431,N12432,N12433,N12434,N12435,N12436,N12437,N12438,
N12439,N12440,N12441,N12442,N12443,N12444,N12445,N12446,N12447,N12448,
N12449,N12450,N12451,N12452,N12453,N12454,N12455,N12456,N12457,N12458,
N12459,N12460,N12461,N12462,N12463,N12464,N12465,N12466,N12467,N12468,
N12469,N12470,N12471,N12472,N12473,N12474,N12475,N12476,N12477,N12478,
N12479,N12480,N12481,N12482,N12483,N12484,N12485,N12486,N12487,N12488,
N12489,N12490,N12491,N12492,N12493,N12494,N12495,N12496,N12497,N12498,
N12499,N12500,N12501,N12502,N12503,N12504,N12505,N12506,N12507,N12508,
N12509,N12510,N12511,N12512,N12513,N12514,N12515,N12516,N12517,N12518,
N12519,N12520,N12521,N12522,N12523,N12524,N12525,N12526,N12527,N12528,
N12529,N12530,N12531,N12532,N12533,N12534,N12535,N12536,N12537,N12538,
N12539,N12540,N12541,N12542,N12543,N12544,N12545,N12546,N12547,N12548,
N12549,N12550,N12551,N12552,N12553,N12554,N12555,N12556,N12557,N12558,
N12559,N12560,N12561,N12562,N12563,N12564,N12565,N12566,N12567,N12568,
N12569,N12570,N12571,N12572,N12573,N12574,N12575,N12576,N12577,N12578,
N12579,N12580,N12581,N12582,N12583,N12584,N12585,N12586,N12587,N12588,
N12589,N12590,N12591,N12592,N12593,N12594,N12595,N12596,N12597,N12598,
N12599,N12600,N12601,N12602,N12603,N12604,N12605,N12606,N12607,N12608,
N12609,N12610,N12611,N12612,N12613,N12614,N12615,N12616,N12617,N12618,
N12619,N12620,N12621,N12622,N12623,N12624,N12625,N12626,N12627,N12628,
N12629,N12630,N12631,N12632,N12633,N12634,N12635,N12636,N12637,N12638,
N12639,N12640,N12641,N12642,N12643,N12644,N12645,N12646,N12647,N12648,
N12649,N12650,N12651,N12652,N12653,N12654,N12655,N12656,N12657,N12658,
N12659,N12660,N12661,N12662,N12663,N12664,N12665,N12666,N12667,N12668,
N12669,N12670,N12671,N12672,N12673,N12674,N12675,N12676,N12677,N12678,
N12679,N12680,N12681,N12682,N12683,N12684,N12685,N12686,N12687,N12688,
N12689,N12690,N12691,N12692,N12693,N12694,N12695,N12696,N12697,N12698,
N12699,N12700,N12701,N12702,N12703,N12704,N12705,N12706,N12707,N12708,
N12709,N12710,N12711,N12712,N12713,N12714,N12715,N12716,N12717,N12718,
N12719,N12720,N12721,N12722,N12723,N12724,N12725,N12726,N12727,N12728,
N12729,N12730,N12731,N12732,N12733,N12734,N12735,N12736,N12737,N12738,
N12739,N12740,N12741,N12742,N12743,N12744,N12745,N12746,N12747,N12748,
N12749,N12750,N12751,N12752,N12753,N12754,N12755,N12756,N12757,N12758,
N12759,N12760,N12761,N12762,N12763,N12764,N12765,N12766,N12767,N12768,
N12769,N12770,N12771,N12772,N12773,N12774,N12775,N12776,N12777,N12778,
N12779,N12780,N12781,N12782,N12783,N12784,N12785,N12786,N12787,N12788,
N12789,N12790,N12791,N12792,N12793,N12794,N12795,N12796,N12797,N12798,
N12799,N12800,N12801,N12802,N12803,N12804,N12805,N12806,N12807,N12808,
N12809,N12810,N12811,N12812,N12813,N12814,N12815,N12816,N12817,N12818,
N12819,N12820,N12821,N12822,N12823,N12824,N12825,N12826,N12827,N12828,
N12829,N12830,N12831,N12832,N12833,N12834,N12835,N12836,N12837,N12838,
N12839,N12840,N12841,N12842,N12843,N12844,N12845,N12846,N12847,N12848,
N12849,N12850,N12851,N12852,N12853,N12854,N12855,N12856,N12857,N12858,
N12859,N12860,N12861,N12862,N12863,N12864,N12865,N12866,N12867,N12868,
N12869,N12870,N12871,N12872,N12873,N12874,N12875,N12876,N12877,N12878,
N12879,N12880,N12881,N12882,N12883,N12884,N12885,N12886,N12887,N12888,
N12889,N12890,N12891,N12892,N12893,N12894,N12895,N12896,N12897,N12898,
N12899,N12900,N12901,N12902,N12903,N12904,N12905,N12906,N12907,N12908,
N12909,N12910,N12911,N12912,N12913,N12914,N12915,N12916,N12917,N12918,
N12919,N12920,N12921,N12922,N12923,N12924,N12925,N12926,N12927,N12928,
N12929,N12930,N12931,N12932,N12933,N12934,N12935,N12936,N12937,N12938,
N12939,N12940,N12941,N12942,N12943,N12944,N12945,N12946,N12947,N12948,
N12949,N12950,N12951,N12952,N12953,N12954,N12955,N12956,N12957,N12958,
N12959,N12960,N12961,N12962,N12963,N12964,N12965,N12966,N12967,N12968,
N12969,N12970,N12971,N12972,N12973,N12974,N12975,N12976,N12977,N12978,
N12979,N12980,N12981,N12982,N12983,N12984,N12985,N12986,N12987,N12988,
N12989,N12990,N12991,N12992,N12993,N12994,N12995,N12996,N12997,N12998,
N12999,N13000,N13001,N13002,N13003,N13004,N13005,N13006,N13007,N13008,
N13009,N13010,N13011,N13012,N13013,N13014,N13015,N13016,N13017,N13018,
N13019,N13020,N13021,N13022,N13023,N13024,N13025,N13026,N13027,N13028,
N13029,N13030,N13031,N13032,N13033,N13034,N13035,N13036,N13037,N13038,
N13039,N13040,N13041,N13042,N13043,N13044,N13045,N13046,N13047,N13048,
N13049,N13050,N13051,N13052,N13053,N13054,N13055,N13056,N13057,N13058,
N13059,N13060,N13061,N13062,N13063,N13064,N13065,N13066,N13067,N13068,
N13069,N13070,N13071,N13072,N13073,N13074,N13075,N13076,N13077,N13078,
N13079,N13080,N13081,N13082,N13083,N13084,N13085,N13086,N13087,N13088,
N13089,N13090,N13091,N13092,N13093,N13094,N13095,N13096,N13097,N13098,
N13099,N13100,N13101,N13102,N13103,N13104,N13105,N13106,N13107,N13108,
N13109,N13110,N13111,N13112,N13113,N13114,N13115,N13116,N13117,N13118,
N13119,N13120,N13121,N13122,N13123,N13124,N13125,N13126,N13127,N13128,
N13129,N13130,N13131,N13132,N13133,N13134,N13135,N13136,N13137,N13138,
N13139,N13140,N13141,N13142,N13143,N13144,N13145,N13146,N13147,N13148,
N13149,N13150,N13151,N13152,N13153,N13154,N13155,N13156,N13157,N13158,
N13159,N13160,N13161,N13162,N13163,N13164,N13165,N13166,N13167,N13168,
N13169,N13170,N13171,N13172,N13173,N13174,N13175,N13176,N13177,N13178,
N13179,N13180,N13181,N13182,N13183,N13184,N13185,N13186,N13187,N13188,
N13189,N13190,N13191,N13192,N13193,N13194,N13195,N13196,N13197,N13198,
N13199,N13200,N13201,N13202,N13203,N13204,N13205,N13206,N13207,N13208,
N13209,N13210,N13211,N13212,N13213,N13214,N13215,N13216,N13217,N13218,
N13219,N13220,N13221,N13222,N13223,N13224,N13225,N13226,N13227,N13228,
N13229,N13230,N13231,N13232,N13233,N13234,N13235,N13236,N13237,N13238,
N13239,N13240,N13241,N13242,N13243,N13244,N13245,N13246,N13247,N13248,
N13249,N13250,N13251,N13252,N13253,N13254,N13255,N13256,N13257,N13258,
N13259,N13260,N13261,N13262,N13263,N13264,N13265,N13266,N13267,N13268,
N13269,N13270,N13271,N13272,N13273,N13274,N13275,N13276,N13277,N13278,
N13279,N13280,N13281,N13282,N13283,N13284,N13285,N13286,N13287,N13288,
N13289,N13290,N13291,N13292,N13293,N13294,N13295,N13296,N13297,N13298,
N13299,N13300,N13301,N13302,N13303,N13304,N13305,N13306,N13307,N13308,
N13309,N13310,N13311,N13312,N13313,N13314,N13315,N13316,N13317,N13318,
N13319,N13320,N13321,N13322,N13323,N13324,N13325,N13326,N13327,N13328,
N13329,N13330,N13331,N13332,N13333,N13334,N13335,N13336,N13337,N13338,
N13339,N13340,N13341,N13342,N13343,N13344,N13345,N13346,N13347,N13348,
N13349,N13350,N13351,N13352,N13353,N13354,N13355,N13356,N13357,N13358,
N13359,N13360,N13361,N13362,N13363,N13364,N13365,N13366,N13367,N13368,
N13369,N13370,N13371,N13372,N13373,N13374,N13375,N13376,N13377,N13378,
N13379,N13380,N13381,N13382,N13383,N13384,N13385,N13386,N13387,N13388,
N13389,N13390,N13391,N13392,N13393,N13394,N13395,N13396,N13397,N13398,
N13399,N13400,N13401,N13402,N13403,N13404,N13405,N13406,N13407,N13408,
N13409,N13410,N13411,N13412,N13413,N13414,N13415,N13416,N13417,N13418,
N13419,N13420,N13421,N13422,N13423,N13424,N13425,N13426,N13427,N13428,
N13429,N13430,N13431,N13432,N13433,N13434,N13435,N13436,N13437,N13438,
N13439,N13440,N13441,N13442,N13443,N13444,N13445,N13446,N13447,N13448,
N13449,N13450,N13451,N13452,N13453,N13454,N13455,N13456,N13457,N13458,
N13459,N13460,N13461,N13462,N13463,N13464,N13465,N13466,N13467,N13468,
N13469,N13470,N13471,N13472,N13473,N13474,N13475,N13476,N13477,N13478,
N13479,N13480,N13481,N13482,N13483,N13484,N13485,N13486,N13487,N13488,
N13489,N13490,N13491,N13492,N13493,N13494,N13495,N13496,N13497,N13498,
N13499,N13500,N13501,N13502,N13503,N13504,N13505,N13506,N13507,N13508,
N13509,N13510,N13511,N13512,N13513,N13514,N13515,N13516,N13517,N13518,
N13519,N13520,N13521,N13522,N13523,N13524,N13525,N13526,N13527,N13528,
N13529,N13530,N13531,N13532,N13533,N13534,N13535,N13536,N13537,N13538,
N13539,N13540,N13541,N13542,N13543,N13544,N13545,N13546,N13547,N13548,
N13549,N13550,N13551,N13552,N13553,N13554,N13555,N13556,N13557,N13558,
N13559,N13560,N13561,N13562,N13563,N13564,N13565,N13566,N13567,N13568,
N13569,N13570,N13571,N13572,N13573,N13574,N13575,N13576,N13577,N13578,
N13579,N13580,N13581,N13582,N13583,N13584,N13585,N13586,N13587,N13588,
N13589,N13590,N13591,N13592,N13593,N13594,N13595,N13596,N13597,N13598,
N13599,N13600,N13601,N13602,N13603,N13604,N13605,N13606,N13607,N13608,
N13609,N13610,N13611,N13612,N13613,N13614,N13615,N13616,N13617,N13618,
N13619,N13620,N13621,N13622,N13623,N13624,N13625,N13626,N13627,N13628,
N13629,N13630,N13631,N13632,N13633,N13634,N13635,N13636,N13637,N13638,
N13639,N13640,N13641,N13642,N13643,N13644,N13645,N13646,N13647,N13648,
N13649,N13650,N13651,N13652,N13653,N13654,N13655,N13656,N13657,N13658,
N13659,N13660,N13661,N13662,N13663,N13664,N13665,N13666,N13667,N13668,
N13669,N13670,N13671,N13672,N13673,N13674,N13675,N13676,N13677,N13678,
N13679,N13680,N13681,N13682,N13683,N13684,N13685,N13686,N13687,N13688,
N13689,N13690,N13691,N13692,N13693,N13694,N13695,N13696,N13697,N13698,
N13699,N13700,N13701,N13702,N13703,N13704,N13705,N13706,N13707,N13708,
N13709,N13710,N13711,N13712,N13713,N13714,N13715,N13716,N13717,N13718,
N13719,N13720,N13721,N13722,N13723,N13724,N13725,N13726,N13727,N13728,
N13729,N13730,N13731,N13732,N13733,N13734,N13735,N13736,N13737,N13738,
N13739,N13740,N13741,N13742,N13743,N13744,N13745,N13746,N13747,N13748,
N13749,N13750,N13751,N13752,N13753,N13754,N13755,N13756,N13757,N13758,
N13759,N13760,N13761,N13762,N13763,N13764,N13765,N13766,N13767,N13768,
N13769,N13770,N13771,N13772,N13773,N13774,N13775,N13776,N13777,N13778,
N13779,N13780,N13781,N13782,N13783,N13784,N13785,N13786,N13787,N13788,
N13789,N13790,N13791,N13792,N13793,N13794,N13795,N13796,N13797,N13798,
N13799,N13800,N13801,N13802,N13803,N13804,N13805,N13806,N13807,N13808,
N13809,N13810,N13811,N13812,N13813,N13814,N13815,N13816,N13817,N13818,
N13819,N13820,N13821,N13822,N13823,N13824,N13825,N13826,N13827,N13828,
N13829,N13830,N13831,N13832,N13833,N13834,N13835,N13836,N13837,N13838,
N13839,N13840,N13841,N13842,N13843,N13844,N13845,N13846,N13847,N13848,
N13849,N13850,N13851,N13852,N13853,N13854,N13855,N13856,N13857,N13858,
N13859,N13860,N13861,N13862,N13863,N13864,N13865,N13866,N13867,N13868,
N13869,N13870,N13871,N13872,N13873,N13874,N13875,N13876,N13877,N13878,
N13879,N13880,N13881,N13882,N13883,N13884,N13885,N13886,N13887,N13888,
N13889,N13890,N13891,N13892,N13893,N13894,N13895,N13896,N13897,N13898,
N13899,N13900,N13901,N13902,N13903,N13904,N13905,N13906,N13907,N13908,
N13909,N13910,N13911,N13912,N13913,N13914,N13915,N13916,N13917,N13918,
N13919,N13920,N13921,N13922,N13923,N13924,N13925,N13926,N13927,N13928,
N13929,N13930,N13931,N13932,N13933,N13934,N13935,N13936,N13937,N13938,
N13939,N13940,N13941,N13942,N13943,N13944,N13945,N13946,N13947,N13948,
N13949,N13950,N13951,N13952,N13953,N13954,N13955,N13956,N13957,N13958,
N13959,N13960,N13961,N13962,N13963,N13964,N13965,N13966,N13967,N13968,
N13969,N13970,N13971,N13972,N13973,N13974,N13975,N13976,N13977,N13978,
N13979,N13980,N13981,N13982,N13983,N13984,N13985,N13986,N13987,N13988,
N13989,N13990,N13991,N13992,N13993,N13994,N13995,N13996,N13997,N13998,
N13999,N14000,N14001,N14002,N14003,N14004,N14005,N14006,N14007,N14008,
N14009,N14010,N14011,N14012,N14013,N14014,N14015,N14016,N14017,N14018,
N14019,N14020,N14021,N14022,N14023,N14024,N14025,N14026,N14027,N14028,
N14029,N14030,N14031,N14032,N14033,N14034,N14035,N14036,N14037,N14038,
N14039,N14040,N14041,N14042,N14043,N14044,N14045,N14046,N14047,N14048,
N14049,N14050,N14051,N14052,N14053,N14054,N14055,N14056,N14057,N14058,
N14059,N14060,N14061,N14062,N14063,N14064,N14065,N14066,N14067,N14068,
N14069,N14070,N14071,N14072,N14073,N14074,N14075,N14076,N14077,N14078,
N14079,N14080,N14081,N14082,N14083,N14084,N14085,N14086,N14087,N14088,
N14089,N14090,N14091,N14092,N14093,N14094,N14095,N14096,N14097,N14098,
N14099,N14100,N14101,N14102,N14103,N14104,N14105,N14106,N14107,N14108,
N14109,N14110,N14111,N14112,N14113,N14114,N14115,N14116,N14117,N14118,
N14119,N14120,N14121,N14122,N14123,N14124,N14125,N14126,N14127,N14128,
N14129,N14130,N14131,N14132,N14133,N14134,N14135,N14136,N14137,N14138,
N14139,N14140,N14141,N14142,N14143,N14144,N14145,N14146,N14147,N14148,
N14149,N14150,N14151,N14152,N14153,N14154,N14155,N14156,N14157,N14158,
N14159,N14160,N14161,N14162,N14163,N14164,N14165,N14166,N14167,N14168,
N14169,N14170,N14171,N14172,N14173,N14174,N14175,N14176,N14177,N14178,
N14179,N14180,N14181,N14182,N14183,N14184,N14185,N14186,N14187,N14188,
N14189,N14190,N14191,N14192,N14193,N14194,N14195,N14196,N14197,N14198,
N14199,N14200,N14201,N14202,N14203,N14204,N14205,N14206,N14207,N14208,
N14209,N14210,N14211,N14212,N14213,N14214,N14215,N14216,N14217,N14218,
N14219,N14220,N14221,N14222,N14223,N14224,N14225,N14226,N14227,N14228,
N14229,N14230,N14231,N14232,N14233,N14234,N14235,N14236,N14237,N14238,
N14239,N14240,N14241,N14242,N14243,N14244,N14245,N14246,N14247,N14248,
N14249,N14250,N14251,N14252,N14253,N14254,N14255,N14256,N14257,N14258,
N14259,N14260,N14261,N14262,N14263,N14264,N14265,N14266,N14267,N14268,
N14269,N14270,N14271,N14272,N14273,N14274,N14275,N14276,N14277,N14278,
N14279,N14280,N14281,N14282,N14283,N14284,N14285,N14286,N14287,N14288,
N14289,N14290,N14291,N14292,N14293,N14294,N14295,N14296,N14297,N14298,
N14299,N14300,N14301,N14302,N14303,N14304,N14305,N14306,N14307,N14308,
N14309,N14310,N14311,N14312,N14313,N14314,N14315,N14316,N14317,N14318,
N14319,N14320,N14321,N14322,N14323,N14324,N14325,N14326,N14327,N14328,
N14329,N14330,N14331,N14332,N14333,N14334,N14335,N14336,N14337,N14338,
N14339,N14340,N14341,N14342,N14343,N14344,N14345,N14346,N14347,N14348,
N14349,N14350,N14351,N14352,N14353,N14354,N14355,N14356,N14357,N14358,
N14359,N14360,N14361,N14362,N14363,N14364,N14365,N14366,N14367,N14368,
N14369,N14370,N14371,N14372,N14373,N14374,N14375,N14376,N14377,N14378,
N14379,N14380,N14381,N14382,N14383,N14384,N14385,N14386,N14387,N14388,
N14389,N14390,N14391,N14392,N14393,N14394,N14395,N14396,N14397,N14398,
N14399,N14400,N14401,N14402,N14403,N14404,N14405,N14406,N14407,N14408,
N14409,N14410,N14411,N14412,N14413,N14414,N14415,N14416,N14417,N14418,
N14419,N14420,N14421,N14422,N14423,N14424,N14425,N14426,N14427,N14428,
N14429,N14430,N14431,N14432,N14433,N14434,N14435,N14436,N14437,N14438,
N14439,N14440,N14441,N14442,N14443,N14444,N14445,N14446,N14447,N14448,
N14449,N14450,N14451,N14452,N14453,N14454,N14455,N14456,N14457,N14458,
N14459,N14460,N14461,N14462,N14463,N14464,N14465,N14466,N14467,N14468,
N14469,N14470,N14471,N14472,N14473,N14474,N14475,N14476,N14477,N14478,
N14479,N14480,N14481,N14482,N14483,N14484,N14485,N14486,N14487,N14488,
N14489,N14490,N14491,N14492,N14493,N14494,N14495,N14496,N14497,N14498,
N14499,N14500,N14501,N14502,N14503,N14504,N14505,N14506,N14507,N14508,
N14509,N14510,N14511,N14512,N14513,N14514,N14515,N14516,N14517,N14518,
N14519,N14520,N14521,N14522,N14523,N14524,N14525,N14526,N14527,N14528,
N14529,N14530,N14531,N14532,N14533,N14534,N14535,N14536,N14537,N14538,
N14539,N14540,N14541,N14542,N14543,N14544,N14545,N14546,N14547,N14548,
N14549,N14550,N14551,N14552,N14553,N14554,N14555,N14556,N14557,N14558,
N14559,N14560,N14561,N14562,N14563,N14564,N14565,N14566,N14567,N14568,
N14569,N14570,N14571,N14572,N14573,N14574,N14575,N14576,N14577,N14578,
N14579,N14580,N14581,N14582,N14583,N14584,N14585,N14586,N14587,N14588,
N14589,N14590,N14591,N14592,N14593,N14594,N14595,N14596,N14597,N14598,
N14599,N14600,N14601,N14602,N14603,N14604,N14605,N14606,N14607,N14608,
N14609,N14610,N14611,N14612,N14613,N14614,N14615,N14616,N14617,N14618,
N14619,N14620,N14621,N14622,N14623,N14624,N14625,N14626,N14627,N14628,
N14629,N14630,N14631,N14632,N14633,N14634,N14635,N14636,N14637,N14638,
N14639,N14640,N14641,N14642,N14643,N14644,N14645,N14646,N14647,N14648,
N14649,N14650,N14651,N14652,N14653,N14654,N14655,N14656,N14657,N14658,
N14659,N14660,N14661,N14662,N14663,N14664,N14665,N14666,N14667,N14668,
N14669,N14670,N14671,N14672,N14673,N14674,N14675,N14676,N14677,N14678,
N14679,N14680,N14681,N14682,N14683,N14684,N14685,N14686,N14687,N14688,
N14689,N14690,N14691,N14692,N14693,N14694,N14695,N14696,N14697,N14698,
N14699,N14700,N14701,N14702,N14703,N14704,N14705,N14706,N14707,N14708,
N14709,N14710,N14711,N14712,N14713,N14714,N14715,N14716,N14717,N14718,
N14719,N14720,N14721,N14722,N14723,N14724,N14725,N14726,N14727,N14728,
N14729,N14730,N14731,N14732,N14733,N14734,N14735,N14736,N14737,N14738,
N14739,N14740,N14741,N14742,N14743,N14744,N14745,N14746,N14747,N14748,
N14749,N14750,N14751,N14752,N14753,N14754,N14755,N14756,N14757,N14758,
N14759,N14760,N14761,N14762,N14763,N14764,N14765,N14766,N14767,N14768,
N14769,N14770,N14771,N14772,N14773,N14774,N14775,N14776,N14777,N14778,
N14779,N14780,N14781,N14782,N14783,N14784,N14785,N14786,N14787,N14788,
N14789,N14790,N14791,N14792,N14793,N14794,N14795,N14796,N14797,N14798,
N14799,N14800,N14801,N14802,N14803,N14804,N14805,N14806,N14807,N14808,
N14809,N14810,N14811,N14812,N14813,N14814,N14815,N14816,N14817,N14818,
N14819,N14820,N14821,N14822,N14823,N14824,N14825,N14826,N14827,N14828,
N14829,N14830,N14831,N14832,N14833,N14834,N14835,N14836,N14837,N14838,
N14839,N14840,N14841,N14842,N14843,N14844,N14845,N14846,N14847,N14848,
N14849,N14850,N14851,N14852,N14853,N14854,N14855,N14856,N14857,N14858,
N14859,N14860,N14861,N14862,N14863,N14864,N14865,N14866,N14867,N14868,
N14869,N14870,N14871,N14872,N14873,N14874,N14875,N14876,N14877,N14878,
N14879,N14880,N14881,N14882,N14883,N14884,N14885,N14886,N14887,N14888,
N14889,N14890,N14891,N14892,N14893,N14894,N14895,N14896,N14897,N14898,
N14899,N14900,N14901,N14902,N14903,N14904,N14905,N14906,N14907,N14908,
N14909,N14910,N14911,N14912,N14913,N14914,N14915,N14916,N14917,N14918,
N14919,N14920,N14921,N14922,N14923,N14924,N14925,N14926,N14927,N14928,
N14929,N14930,N14931,N14932,N14933,N14934,N14935,N14936,N14937,N14938,
N14939,N14940,N14941,N14942,N14943,N14944,N14945,N14946,N14947,N14948,
N14949,N14950,N14951,N14952,N14953,N14954,N14955,N14956,N14957,N14958,
N14959,N14960,N14961,N14962,N14963,N14964,N14965,N14966,N14967,N14968,
N14969,N14970,N14971,N14972,N14973,N14974,N14975,N14976,N14977,N14978,
N14979,N14980,N14981,N14982,N14983,N14984,N14985,N14986,N14987,N14988,
N14989,N14990,N14991,N14992,N14993,N14994,N14995,N14996,N14997,N14998,
N14999,N15000,N15001,N15002,N15003,N15004,N15005,N15006,N15007,N15008,
N15009,N15010,N15011,N15012,N15013,N15014,N15015,N15016,N15017,N15018,
N15019,N15020,N15021,N15022,N15023,N15024,N15025,N15026,N15027,N15028,
N15029,N15030,N15031,N15032,N15033,N15034,N15035,N15036,N15037,N15038,
N15039,N15040,N15041,N15042,N15043,N15044,N15045,N15046,N15047,N15048,
N15049,N15050,N15051,N15052,N15053,N15054,N15055,N15056,N15057,N15058,
N15059,N15060,N15061,N15062,N15063,N15064,N15065,N15066,N15067,N15068,
N15069,N15070,N15071,N15072,N15073,N15074,N15075,N15076,N15077,N15078,
N15079,N15080,N15081,N15082,N15083,N15084,N15085,N15086,N15087,N15088,
N15089,N15090,N15091,N15092,N15093,N15094,N15095,N15096,N15097,N15098,
N15099,N15100,N15101,N15102,N15103,N15104,N15105,N15106,N15107,N15108,
N15109,N15110,N15111,N15112,N15113,N15114,N15115,N15116,N15117,N15118,
N15119,N15120,N15121,N15122,N15123,N15124,N15125,N15126,N15127,N15128,
N15129,N15130,N15131,N15132,N15133,N15134,N15135,N15136,N15137,N15138,
N15139,N15140,N15141,N15142,N15143,N15144,N15145,N15146,N15147,N15148,
N15149,N15150,N15151,N15152,N15153,N15154,N15155,N15156,N15157,N15158,
N15159,N15160,N15161,N15162,N15163,N15164,N15165,N15166,N15167,N15168,
N15169,N15170,N15171,N15172,N15173,N15174,N15175,N15176,N15177,N15178,
N15179,N15180,N15181,N15182,N15183,N15184,N15185,N15186,N15187,N15188,
N15189,N15190,N15191,N15192,N15193,N15194,N15195,N15196,N15197,N15198,
N15199,N15200,N15201,N15202,N15203,N15204,N15205,N15206,N15207,N15208,
N15209,N15210,N15211,N15212,N15213,N15214,N15215,N15216,N15217,N15218,
N15219,N15220,N15221,N15222,N15223,N15224,N15225,N15226,N15227,N15228,
N15229,N15230,N15231,N15232,N15233,N15234,N15235,N15236,N15237,N15238,
N15239,N15240,N15241,N15242,N15243,N15244,N15245,N15246,N15247,N15248,
N15249,N15250,N15251,N15252,N15253,N15254,N15255,N15256,N15257,N15258,
N15259,N15260,N15261,N15262,N15263,N15264,N15265,N15266,N15267,N15268,
N15269,N15270,N15271,N15272,N15273,N15274,N15275,N15276,N15277,N15278,
N15279,N15280,N15281,N15282,N15283,N15284,N15285,N15286,N15287,N15288,
N15289,N15290,N15291,N15292,N15293,N15294,N15295,N15296,N15297,N15298,
N15299,N15300,N15301,N15302,N15303,N15304,N15305,N15306,N15307,N15308,
N15309,N15310,N15311,N15312,N15313,N15314,N15315,N15316,N15317,N15318,
N15319,N15320,N15321,N15322,N15323,N15324,N15325,N15326,N15327,N15328,
N15329,N15330,N15331,N15332,N15333,N15334,N15335,N15336,N15337,N15338,
N15339,N15340,N15341,N15342,N15343,N15344,N15345,N15346,N15347,N15348,
N15349,N15350,N15351,N15352,N15353,N15354,N15355,N15356,N15357,N15358,
N15359,N15360,N15361,N15362,N15363,N15364,N15365,N15366,N15367,N15368,
N15369,N15370,N15371,N15372,N15373,N15374,N15375,N15376,N15377,N15378,
N15379,N15380,N15381,N15382,N15383,N15384,N15385,N15386,N15387,N15388,
N15389,N15390,N15391,N15392,N15393,N15394,N15395,N15396,N15397,N15398,
N15399,N15400,N15401,N15402,N15403,N15404,N15405,N15406,N15407,N15408,
N15409,N15410,N15411,N15412,N15413,N15414,N15415,N15416,N15417,N15418,
N15419,N15420,N15421,N15422,N15423,N15424,N15425,N15426,N15427,N15428,
N15429,N15430,N15431,N15432,N15433,N15434,N15435,N15436,N15437,N15438,
N15439,N15440,N15441,N15442,N15443,N15444,N15445,N15446,N15447,N15448,
N15449,N15450,N15451,N15452,N15453,N15454,N15455,N15456,N15457,N15458,
N15459,N15460,N15461,N15462,N15463,N15464,N15465,N15466,N15467,N15468,
N15469,N15470,N15471,N15472,N15473,N15474,N15475,N15476,N15477,N15478,
N15479,N15480,N15481,N15482,N15483,N15484,N15485,N15486,N15487,N15488,
N15489,N15490,N15491,N15492,N15493,N15494,N15495,N15496,N15497,N15498,
N15499,N15500,N15501,N15502,N15503,N15504,N15505,N15506,N15507,N15508,
N15509,N15510,N15511,N15512,N15513,N15514,N15515,N15516,N15517,N15518,
N15519,N15520,N15521,N15522,N15523,N15524,N15525,N15526,N15527,N15528,
N15529,N15530,N15531,N15532,N15533,N15534,N15535,N15536,N15537,N15538,
N15539,N15540,N15541,N15542,N15543,N15544,N15545,N15546,N15547,N15548,
N15549,N15550,N15551,N15552,N15553,N15554,N15555,N15556,N15557,N15558,
N15559,N15560,N15561,N15562,N15563,N15564,N15565,N15566,N15567,N15568,
N15569,N15570,N15571,N15572,N15573,N15574,N15575,N15576,N15577,N15578,
N15579,N15580,N15581,N15582,N15583,N15584,N15585,N15586,N15587,N15588,
N15589,N15590,N15591,N15592,N15593,N15594,N15595,N15596,N15597,N15598,
N15599,N15600,N15601,N15602,N15603,N15604,N15605,N15606,N15607,N15608,
N15609,N15610,N15611,N15612,N15613,N15614,N15615,N15616,N15617,N15618,
N15619,N15620,N15621,N15622,N15623,N15624,N15625,N15626,N15627,N15628,
N15629,N15630,N15631,N15632,N15633,N15634,N15635,N15636,N15637,N15638,
N15639,N15640,N15641,N15642,N15643,N15644,N15645,N15646,N15647,N15648,
N15649,N15650,N15651,N15652,N15653,N15654,N15655,N15656,N15657,N15658,
N15659,N15660,N15661,N15662,N15663,N15664,N15665,N15666,N15667,N15668,
N15669,N15670,N15671,N15672,N15673,N15674,N15675,N15676,N15677,N15678,
N15679,N15680,N15681,N15682,N15683,N15684,N15685,N15686,N15687,N15688,
N15689,N15690,N15691,N15692,N15693,N15694,N15695,N15696,N15697,N15698,
N15699,N15700,N15701,N15702,N15703,N15704,N15705,N15706,N15707,N15708,
N15709,N15710,N15711,N15712,N15713,N15714,N15715,N15716,N15717,N15718,
N15719,N15720,N15721,N15722,N15723,N15724,N15725,N15726,N15727,N15728,
N15729,N15730,N15731,N15732,N15733,N15734,N15735,N15736,N15737,N15738,
N15739,N15740,N15741,N15742,N15743,N15744,N15745,N15746,N15747,N15748,
N15749,N15750,N15751,N15752,N15753,N15754,N15755,N15756,N15757,N15758,
N15759,N15760,N15761,N15762,N15763,N15764,N15765,N15766,N15767,N15768,
N15769,N15770,N15771,N15772,N15773,N15774,N15775,N15776,N15777,N15778,
N15779,N15780,N15781,N15782,N15783,N15784,N15785,N15786,N15787,N15788,
N15789,N15790,N15791,N15792,N15793,N15794,N15795,N15796,N15797,N15798,
N15799,N15800,N15801,N15802,N15803,N15804,N15805,N15806,N15807,N15808,
N15809,N15810,N15811,N15812,N15813,N15814,N15815,N15816,N15817,N15818,
N15819,N15820,N15821,N15822,N15823,N15824,N15825,N15826,N15827,N15828,
N15829,N15830,N15831,N15832,N15833,N15834,N15835,N15836,N15837,N15838,
N15839,N15840,N15841,N15842,N15843,N15844,N15845,N15846,N15847,N15848,
N15849,N15850,N15851,N15852,N15853,N15854,N15855,N15856,N15857,N15858,
N15859,N15860,N15861,N15862,N15863,N15864,N15865,N15866,N15867,N15868,
N15869,N15870,N15871,N15872,N15873,N15874,N15875,N15876,N15877,N15878,
N15879,N15880,N15881,N15882,N15883,N15884,N15885,N15886,N15887,N15888,
N15889,N15890,N15891,N15892,N15893,N15894,N15895,N15896,N15897,N15898,
N15899,N15900,N15901,N15902,N15903,N15904,N15905,N15906,N15907,N15908,
N15909,N15910,N15911,N15912,N15913,N15914,N15915,N15916,N15917,N15918,
N15919,N15920,N15921,N15922,N15923,N15924,N15925,N15926,N15927,N15928,
N15929,N15930,N15931,N15932,N15933,N15934,N15935,N15936,N15937,N15938,
N15939,N15940,N15941,N15942,N15943,N15944,N15945,N15946,N15947,N15948,
N15949,N15950,N15951,N15952,N15953,N15954,N15955,N15956,N15957,N15958,
N15959,N15960,N15961,N15962,N15963,N15964,N15965,N15966,N15967,N15968,
N15969,N15970,N15971,N15972,N15973,N15974,N15975,N15976,N15977,N15978,
N15979,N15980,N15981,N15982,N15983,N15984,N15985,N15986,N15987,N15988,
N15989,N15990,N15991,N15992,N15993,N15994,N15995,N15996,N15997,N15998,
N15999,N16000,N16001,N16002,N16003,N16004,N16005,N16006,N16007,N16008,
N16009,N16010,N16011,N16012,N16013,N16014,N16015,N16016,N16017,N16018,
N16019,N16020,N16021,N16022,N16023,N16024,N16025,N16026,N16027,N16028,
N16029,N16030,N16031,N16032,N16033,N16034,N16035,N16036,N16037,N16038,
N16039,N16040,N16041,N16042,N16043,N16044,N16045,N16046,N16047,N16048,
N16049,N16050,N16051,N16052,N16053,N16054,N16055,N16056,N16057,N16058,
N16059,N16060,N16061,N16062,N16063,N16064,N16065,N16066,N16067,N16068,
N16069,N16070,N16071,N16072,N16073,N16074,N16075,N16076,N16077,N16078,
N16079,N16080,N16081,N16082,N16083,N16084,N16085,N16086,N16087,N16088,
N16089,N16090,N16091,N16092,N16093,N16094,N16095,N16096,N16097,N16098,
N16099,N16100,N16101,N16102,N16103,N16104,N16105,N16106,N16107,N16108,
N16109,N16110,N16111,N16112,N16113,N16114,N16115,N16116,N16117,N16118,
N16119,N16120,N16121,N16122,N16123,N16124,N16125,N16126,N16127,N16128,
N16129,N16130,N16131,N16132,N16133,N16134,N16135,N16136,N16137,N16138,
N16139,N16140,N16141,N16142,N16143,N16144,N16145,N16146,N16147,N16148,
N16149,N16150,N16151,N16152,N16153,N16154,N16155,N16156,N16157,N16158,
N16159,N16160,N16161,N16162,N16163,N16164,N16165,N16166,N16167,N16168,
N16169,N16170,N16171,N16172,N16173,N16174,N16175,N16176,N16177,N16178,
N16179,N16180,N16181,N16182,N16183,N16184,N16185,N16186,N16187,N16188,
N16189,N16190,N16191,N16192,N16193,N16194,N16195,N16196,N16197,N16198,
N16199,N16200,N16201,N16202,N16203,N16204,N16205,N16206,N16207,N16208,
N16209,N16210,N16211,N16212,N16213,N16214,N16215,N16216,N16217,N16218,
N16219,N16220,N16221,N16222,N16223,N16224,N16225,N16226,N16227,N16228,
N16229,N16230,N16231,N16232,N16233,N16234,N16235,N16236,N16237,N16238,
N16239,N16240,N16241,N16242,N16243,N16244,N16245,N16246,N16247,N16248,
N16249,N16250,N16251,N16252,N16253,N16254,N16255,N16256,N16257,N16258,
N16259,N16260,N16261,N16262,N16263,N16264,N16265,N16266,N16267,N16268,
N16269,N16270,N16271,N16272,N16273,N16274,N16275,N16276,N16277,N16278,
N16279,N16280,N16281,N16282,N16283,N16284,N16285,N16286,N16287,N16288,
N16289,N16290,N16291,N16292,N16293,N16294,N16295,N16296,N16297,N16298,
N16299,N16300,N16301,N16302,N16303,N16304,N16305,N16306,N16307,N16308,
N16309,N16310,N16311,N16312,N16313,N16314,N16315,N16316,N16317,N16318,
N16319,N16320,N16321,N16322,N16323,N16324,N16325,N16326,N16327,N16328,
N16329,N16330,N16331,N16332,N16333,N16334,N16335,N16336,N16337,N16338,
N16339,N16340,N16341,N16342,N16343,N16344,N16345,N16346,N16347,N16348,
N16349,N16350,N16351,N16352,N16353,N16354,N16355,N16356,N16357,N16358,
N16359,N16360,N16361,N16362,N16363,N16364,N16365,N16366,N16367,N16368,
N16369,N16370,N16371,N16372,N16373,N16374,N16375,N16376,N16377,N16378,
N16379,N16380,N16381,N16382,N16383,N16384,N16385,N16386,N16387,N16388,
N16389,N16390,N16391,N16392,N16393,N16394,N16395,N16396,N16397,N16398,
N16399,N16400,N16401,N16402,N16403,N16404,N16405,N16406,N16407,N16408,
N16409,N16410,N16411,N16412,N16413,N16414,N16415,N16416,N16417,N16418,
N16419,N16420,N16421,N16422,N16423,N16424,N16425,N16426,N16427,N16428,
N16429,N16430,N16431,N16432,N16433,N16434,N16435,N16436,N16437,N16438,
N16439,N16440,N16441,N16442,N16443,N16444,N16445,N16446,N16447,N16448,
N16449,N16450,N16451,N16452,N16453,N16454,N16455,N16456,N16457,N16458,
N16459,N16460,N16461,N16462,N16463,N16464,N16465,N16466,N16467,N16468,
N16469,N16470,N16471,N16472,N16473,N16474,N16475,N16476,N16477,N16478,
N16479,N16480,N16481,N16482,N16483,N16484,N16485,N16486,N16487,N16488,
N16489,N16490,N16491,N16492,N16493,N16494,N16495,N16496,N16497,N16498,
N16499,N16500,N16501,N16502,N16503,N16504,N16505,N16506,N16507,N16508,
N16509,N16510,N16511,N16512,N16513,N16514,N16515,N16516,N16517,N16518,
N16519,N16520,N16521,N16522,N16523,N16524,N16525,N16526,N16527,N16528,
N16529,N16530,N16531,N16532,N16533,N16534,N16535,N16536,N16537,N16538,
N16539,N16540,N16541,N16542,N16543,N16544,N16545,N16546,N16547,N16548,
N16549,N16550,N16551,N16552,N16553,N16554,N16555,N16556,N16557,N16558,
N16559,N16560,N16561,N16562,N16563,N16564,N16565,N16566,N16567,N16568,
N16569,N16570,N16571,N16572,N16573,N16574,N16575,N16576,N16577,N16578,
N16579,N16580,N16581,N16582,N16583,N16584,N16585,N16586,N16587,N16588,
N16589,N16590,N16591,N16592,N16593,N16594,N16595,N16596,N16597,N16598,
N16599,N16600,N16601,N16602,N16603,N16604,N16605,N16606,N16607,N16608,
N16609,N16610,N16611,N16612,N16613,N16614,N16615,N16616,N16617,N16618,
N16619,N16620,N16621,N16622,N16623,N16624,N16625,N16626,N16627,N16628,
N16629,N16630,N16631,N16632,N16633,N16634,N16635,N16636,N16637,N16638,
N16639,N16640,N16641,N16642,N16643,N16644,N16645,N16646,N16647,N16648,
N16649,N16650,N16651,N16652,N16653,N16654,N16655,N16656,N16657,N16658,
N16659,N16660,N16661,N16662,N16663,N16664,N16665,N16666,N16667,N16668,
N16669,N16670,N16671,N16672,N16673,N16674,N16675,N16676,N16677,N16678,
N16679,N16680,N16681,N16682,N16683,N16684,N16685,N16686,N16687,N16688,
N16689,N16690,N16691,N16692,N16693,N16694,N16695,N16696,N16697,N16698,
N16699,N16700,N16701,N16702,N16703,N16704,N16705,N16706,N16707,N16708,
N16709,N16710,N16711,N16712,N16713,N16714,N16715,N16716,N16717,N16718,
N16719,N16720,N16721,N16722,N16723,N16724,N16725,N16726,N16727,N16728,
N16729,N16730,N16731,N16732,N16733,N16734,N16735,N16736,N16737,N16738,
N16739,N16740,N16741,N16742,N16743,N16744,N16745,N16746,N16747,N16748,
N16749,N16750,N16751,N16752,N16753,N16754,N16755,N16756,N16757,N16758,
N16759,N16760,N16761,N16762,N16763,N16764,N16765,N16766,N16767,N16768,
N16769,N16770,N16771,N16772,N16773,N16774,N16775,N16776,N16777,N16778,
N16779,N16780,N16781,N16782,N16783,N16784,N16785,N16786,N16787,N16788,
N16789,N16790,N16791,N16792,N16793,N16794,N16795,N16796,N16797,N16798,
N16799,N16800,N16801,N16802,N16803,N16804,N16805,N16806,N16807,N16808,
N16809,N16810,N16811,N16812,N16813,N16814,N16815,N16816,N16817,N16818,
N16819,N16820,N16821,N16822,N16823,N16824,N16825,N16826,N16827,N16828,
N16829,N16830,N16831,N16832,N16833,N16834,N16835,N16836,N16837,N16838,
N16839,N16840,N16841,N16842,N16843,N16844,N16845,N16846,N16847,N16848,
N16849,N16850,N16851,N16852,N16853,N16854,N16855,N16856,N16857,N16858,
N16859,N16860,N16861,N16862,N16863,N16864,N16865,N16866,N16867,N16868,
N16869,N16870,N16871,N16872,N16873,N16874,N16875,N16876,N16877,N16878,
N16879,N16880,N16881,N16882,N16883,N16884,N16885,N16886,N16887,N16888,
N16889,N16890,N16891,N16892,N16893,N16894,N16895,N16896,N16897,N16898,
N16899,N16900,N16901,N16902,N16903,N16904,N16905,N16906,N16907,N16908,
N16909,N16910,N16911,N16912,N16913,N16914,N16915,N16916,N16917,N16918,
N16919,N16920,N16921,N16922,N16923,N16924,N16925,N16926,N16927,N16928,
N16929,N16930,N16931,N16932,N16933,N16934,N16935,N16936,N16937,N16938,
N16939,N16940,N16941,N16942,N16943,N16944,N16945,N16946,N16947,N16948,
N16949,N16950,N16951,N16952,N16953,N16954,N16955,N16956,N16957,N16958,
N16959,N16960,N16961,N16962,N16963,N16964,N16965,N16966,N16967,N16968,
N16969,N16970,N16971,N16972,N16973,N16974,N16975,N16976,N16977,N16978,
N16979,N16980,N16981,N16982,N16983,N16984,N16985,N16986,N16987,N16988,
N16989,N16990,N16991,N16992,N16993,N16994,N16995,N16996,N16997,N16998,
N16999,N17000,N17001,N17002,N17003,N17004,N17005,N17006,N17007,N17008,
N17009,N17010,N17011,N17012,N17013,N17014,N17015,N17016,N17017,N17018,
N17019,N17020,N17021,N17022,N17023,N17024,N17025,N17026,N17027,N17028,
N17029,N17030,N17031,N17032,N17033,N17034,N17035,N17036,N17037,N17038,
N17039,N17040,N17041,N17042,N17043,N17044,N17045,N17046,N17047,N17048,
N17049,N17050,N17051,N17052,N17053,N17054,N17055,N17056,N17057,N17058,
N17059,N17060,N17061,N17062,N17063,N17064,N17065,N17066,N17067,N17068,
N17069,N17070,N17071,N17072,N17073,N17074,N17075,N17076,N17077,N17078,
N17079,N17080,N17081,N17082,N17083,N17084,N17085,N17086,N17087,N17088,
N17089,N17090,N17091,N17092,N17093,N17094,N17095,N17096,N17097,N17098,
N17099,N17100,N17101,N17102,N17103,N17104,N17105,N17106,N17107,N17108,
N17109,N17110,N17111,N17112,N17113,N17114,N17115,N17116,N17117,N17118,
N17119,N17120,N17121,N17122,N17123,N17124,N17125,N17126,N17127,N17128,
N17129,N17130,N17131,N17132,N17133,N17134,N17135,N17136,N17137,N17138,
N17139,N17140,N17141,N17142,N17143,N17144,N17145,N17146,N17147,N17148,
N17149,N17150,N17151,N17152,N17153,N17154,N17155,N17156,N17157,N17158,
N17159,N17160,N17161,N17162,N17163,N17164,N17165,N17166,N17167,N17168,
N17169,N17170,N17171,N17172,N17173,N17174,N17175,N17176,N17177,N17178,
N17179,N17180,N17181,N17182,N17183,N17184,N17185,N17186,N17187,N17188,
N17189,N17190,N17191,N17192,N17193,N17194,N17195,N17196,N17197,N17198,
N17199,N17200,N17201,N17202,N17203,N17204,N17205,N17206,N17207,N17208,
N17209,N17210,N17211,N17212,N17213,N17214,N17215,N17216,N17217,N17218,
N17219,N17220,N17221,N17222,N17223,N17224,N17225,N17226,N17227,N17228,
N17229,N17230,N17231,N17232,N17233,N17234,N17235,N17236,N17237,N17238,
N17239,N17240,N17241,N17242,N17243,N17244,N17245,N17246,N17247,N17248,
N17249,N17250,N17251,N17252,N17253,N17254,N17255,N17256,N17257,N17258,
N17259,N17260,N17261,N17262,N17263,N17264,N17265,N17266,N17267,N17268,
N17269,N17270,N17271,N17272,N17273,N17274,N17275,N17276,N17277,N17278,
N17279,N17280,N17281,N17282,N17283,N17284,N17285,N17286,N17287,N17288,
N17289,N17290,N17291,N17292,N17293,N17294,N17295,N17296,N17297,N17298,
N17299,N17300,N17301,N17302,N17303,N17304,N17305,N17306,N17307,N17308,
N17309,N17310,N17311,N17312,N17313,N17314,N17315,N17316,N17317,N17318,
N17319,N17320,N17321,N17322,N17323,N17324,N17325,N17326,N17327,N17328,
N17329,N17330,N17331,N17332,N17333,N17334,N17335,N17336,N17337,N17338,
N17339,N17340,N17341,N17342,N17343,N17344,N17345,N17346,N17347,N17348,
N17349,N17350,N17351,N17352,N17353,N17354,N17355,N17356,N17357,N17358,
N17359,N17360,N17361,N17362,N17363,N17364,N17365,N17366,N17367,N17368,
N17369,N17370,N17371,N17372,N17373,N17374,N17375,N17376,N17377,N17378,
N17379,N17380,N17381,N17382,N17383,N17384,N17385,N17386,N17387,N17388,
N17389,N17390,N17391,N17392,N17393,N17394,N17395,N17396,N17397,N17398,
N17399,N17400,N17401,N17402,N17403,N17404,N17405,N17406,N17407,N17408,
N17409,N17410,N17411,N17412,N17413,N17414,N17415,N17416,N17417,N17418,
N17419,N17420,N17421,N17422,N17423,N17424,N17425,N17426,N17427,N17428,
N17429,N17430,N17431,N17432,N17433,N17434,N17435,N17436,N17437,N17438,
N17439,N17440,N17441,N17442,N17443,N17444,N17445,N17446,N17447,N17448,
N17449,N17450,N17451,N17452,N17453,N17454,N17455,N17456,N17457,N17458,
N17459,N17460,N17461,N17462,N17463,N17464,N17465,N17466,N17467,N17468,
N17469,N17470,N17471,N17472,N17473,N17474,N17475,N17476,N17477,N17478,
N17479,N17480,N17481,N17482,N17483,N17484,N17485,N17486,N17487,N17488,
N17489,N17490,N17491,N17492,N17493,N17494,N17495,N17496,N17497,N17498,
N17499,N17500,N17501,N17502,N17503,N17504,N17505,N17506,N17507,N17508,
N17509,N17510,N17511,N17512,N17513,N17514,N17515,N17516,N17517,N17518,
N17519,N17520,N17521,N17522,N17523,N17524,N17525,N17526,N17527,N17528,
N17529,N17530,N17531,N17532,N17533,N17534,N17535,N17536,N17537,N17538,
N17539,N17540,N17541,N17542,N17543,N17544,N17545,N17546,N17547,N17548,
N17549,N17550,N17551,N17552,N17553,N17554,N17555,N17556,N17557,N17558,
N17559,N17560,N17561,N17562,N17563,N17564,N17565,N17566,N17567,N17568,
N17569,N17570,N17571,N17572,N17573,N17574,N17575,N17576,N17577,N17578,
N17579,N17580,N17581,N17582,N17583,N17584,N17585,N17586,N17587,N17588,
N17589,N17590,N17591,N17592,N17593,N17594,N17595,N17596,N17597,N17598,
N17599,N17600,N17601,N17602,N17603,N17604,N17605,N17606,N17607,N17608,
N17609,N17610,N17611,N17612,N17613,N17614,N17615,N17616,N17617,N17618,
N17619,N17620,N17621,N17622,N17623,N17624,N17625,N17626,N17627,N17628,
N17629,N17630,N17631,N17632,N17633,N17634,N17635,N17636,N17637,N17638,
N17639,N17640,N17641,N17642,N17643,N17644,N17645,N17646,N17647,N17648,
N17649,N17650,N17651,N17652,N17653,N17654,N17655,N17656,N17657,N17658,
N17659,N17660,N17661,N17662,N17663,N17664,N17665,N17666,N17667,N17668,
N17669,N17670,N17671,N17672,N17673,N17674,N17675,N17676,N17677,N17678,
N17679,N17680,N17681,N17682,N17683,N17684,N17685,N17686,N17687,N17688,
N17689,N17690,N17691,N17692,N17693,N17694,N17695,N17696,N17697,N17698,
N17699,N17700,N17701,N17702,N17703,N17704,N17705,N17706,N17707,N17708,
N17709,N17710,N17711,N17712,N17713,N17714,N17715,N17716,N17717,N17718,
N17719,N17720,N17721,N17722,N17723,N17724,N17725,N17726,N17727,N17728,
N17729,N17730,N17731,N17732,N17733,N17734,N17735,N17736,N17737,N17738,
N17739,N17740,N17741,N17742,N17743,N17744,N17745,N17746,N17747,N17748,
N17749,N17750,N17751,N17752,N17753,N17754,N17755,N17756,N17757,N17758,
N17759,N17760,N17761,N17762,N17763,N17764,N17765,N17766,N17767,N17768,
N17769,N17770,N17771,N17772,N17773,N17774,N17775,N17776,N17777,N17778,
N17779,N17780,N17781,N17782,N17783,N17784,N17785,N17786,N17787,N17788,
N17789,N17790,N17791,N17792,N17793,N17794,N17795,N17796,N17797,N17798,
N17799,N17800,N17801,N17802,N17803,N17804,N17805,N17806,N17807,N17808,
N17809,N17810,N17811,N17812,N17813,N17814,N17815,N17816,N17817,N17818,
N17819,N17820,N17821,N17822,N17823,N17824,N17825,N17826,N17827,N17828,
N17829,N17830,N17831,N17832,N17833,N17834,N17835,N17836,N17837,N17838,
N17839,N17840,N17841,N17842,N17843,N17844,N17845,N17846,N17847,N17848,
N17849,N17850,N17851,N17852,N17853,N17854,N17855,N17856,N17857,N17858,
N17859,N17860,N17861,N17862,N17863,N17864,N17865,N17866,N17867,N17868,
N17869,N17870,N17871,N17872,N17873,N17874,N17875,N17876,N17877,N17878,
N17879,N17880,N17881,N17882,N17883,N17884,N17885,N17886,N17887,N17888,
N17889,N17890,N17891,N17892,N17893,N17894,N17895,N17896,N17897,N17898,
N17899,N17900,N17901,N17902,N17903,N17904,N17905,N17906,N17907,N17908,
N17909,N17910,N17911,N17912,N17913,N17914,N17915,N17916,N17917,N17918,
N17919,N17920,N17921,N17922,N17923,N17924,N17925,N17926,N17927,N17928,
N17929,N17930,N17931,N17932,N17933,N17934,N17935,N17936,N17937,N17938,
N17939,N17940,N17941,N17942,N17943,N17944,N17945,N17946,N17947,N17948,
N17949,N17950,N17951,N17952,N17953,N17954,N17955,N17956,N17957,N17958,
N17959,N17960,N17961,N17962,N17963,N17964,N17965,N17966,N17967,N17968,
N17969,N17970,N17971,N17972,N17973,N17974,N17975,N17976,N17977,N17978,
N17979,N17980,N17981,N17982,N17983,N17984,N17985,N17986,N17987,N17988,
N17989,N17990,N17991,N17992,N17993,N17994,N17995,N17996,N17997,N17998,
N17999,N18000,N18001,N18002,N18003,N18004,N18005,N18006,N18007,N18008,
N18009,N18010,N18011,N18012,N18013,N18014,N18015,N18016,N18017,N18018,
N18019,N18020,N18021,N18022,N18023,N18024,N18025,N18026,N18027,N18028,
N18029,N18030,N18031,N18032,N18033,N18034,N18035,N18036,N18037,N18038,
N18039,N18040,N18041,N18042,N18043,N18044,N18045,N18046,N18047,N18048,
N18049,N18050,N18051,N18052,N18053,N18054,N18055,N18056,N18057,N18058,
N18059,N18060,N18061,N18062,N18063,N18064,N18065,N18066,N18067,N18068,
N18069,N18070,N18071,N18072,N18073,N18074,N18075,N18076,N18077,N18078,
N18079,N18080,N18081,N18082,N18083,N18084,N18085,N18086,N18087,N18088,
N18089,N18090,N18091,N18092,N18093,N18094,N18095,N18096,N18097,N18098,
N18099,N18100,N18101,N18102,N18103,N18104,N18105,N18106,N18107,N18108,
N18109,N18110,N18111,N18112,N18113,N18114,N18115,N18116,N18117,N18118,
N18119,N18120,N18121,N18122,N18123,N18124,N18125,N18126,N18127,N18128,
N18129,N18130,N18131,N18132,N18133,N18134,N18135,N18136,N18137,N18138,
N18139,N18140,N18141,N18142,N18143,N18144,N18145,N18146,N18147,N18148,
N18149,N18150,N18151,N18152,N18153,N18154,N18155,N18156,N18157,N18158,
N18159,N18160,N18161,N18162,N18163,N18164,N18165,N18166,N18167,N18168,
N18169,N18170,N18171,N18172,N18173,N18174,N18175,N18176,N18177,N18178,
N18179,N18180,N18181,N18182,N18183,N18184,N18185,N18186,N18187,N18188,
N18189,N18190,N18191,N18192,N18193,N18194,N18195,N18196,N18197,N18198,
N18199,N18200,N18201,N18202,N18203,N18204,N18205,N18206,N18207,N18208,
N18209,N18210,N18211,N18212,N18213,N18214,N18215,N18216,N18217,N18218,
N18219,N18220,N18221,N18222,N18223,N18224,N18225,N18226,N18227,N18228,
N18229,N18230,N18231,N18232,N18233,N18234,N18235,N18236,N18237,N18238,
N18239,N18240,N18241,N18242,N18243,N18244,N18245,N18246,N18247,N18248,
N18249,N18250,N18251,N18252,N18253,N18254,N18255,N18256,N18257,N18258,
N18259,N18260,N18261,N18262,N18263,N18264,N18265,N18266,N18267,N18268,
N18269,N18270,N18271,N18272,N18273,N18274,N18275,N18276,N18277,N18278,
N18279,N18280,N18281,N18282,N18283,N18284,N18285,N18286,N18287,N18288,
N18289,N18290,N18291,N18292,N18293,N18294,N18295,N18296,N18297,N18298,
N18299,N18300,N18301,N18302,N18303,N18304,N18305,N18306,N18307,N18308,
N18309,N18310,N18311,N18312,N18313,N18314,N18315,N18316,N18317,N18318,
N18319,N18320,N18321,N18322,N18323,N18324,N18325,N18326,N18327,N18328,
N18329,N18330,N18331,N18332,N18333,N18334,N18335,N18336,N18337,N18338,
N18339,N18340,N18341,N18342,N18343,N18344,N18345,N18346,N18347,N18348,
N18349,N18350,N18351,N18352,N18353,N18354,N18355,N18356,N18357,N18358,
N18359,N18360,N18361,N18362,N18363,N18364,N18365,N18366,N18367,N18368,
N18369,N18370,N18371,N18372,N18373,N18374,N18375,N18376,N18377,N18378,
N18379,N18380,N18381,N18382,N18383,N18384,N18385,N18386,N18387,N18388,
N18389,N18390,N18391,N18392,N18393,N18394,N18395,N18396,N18397,N18398,
N18399,N18400,N18401,N18402,N18403,N18404,N18405,N18406,N18407,N18408,
N18409,N18410,N18411,N18412,N18413,N18414,N18415,N18416,N18417,N18418,
N18419,N18420,N18421,N18422,N18423,N18424,N18425,N18426,N18427,N18428,
N18429,N18430,N18431,N18432,N18433,N18434,N18435,N18436,N18437,N18438,
N18439,N18440,N18441,N18442,N18443,N18444,N18445,N18446,N18447,N18448,
N18449,N18450,N18451,N18452,N18453,N18454,N18455,N18456,N18457,N18458,
N18459,N18460,N18461,N18462,N18463,N18464,N18465,N18466,N18467,N18468,
N18469,N18470,N18471,N18472,N18473,N18474,N18475,N18476,N18477,N18478,
N18479,N18480,N18481,N18482,N18483,N18484,N18485,N18486,N18487,N18488,
N18489,N18490,N18491,N18492,N18493,N18494,N18495,N18496,N18497,N18498,
N18499,N18500,N18501,N18502,N18503,N18504,N18505,N18506,N18507,N18508,
N18509,N18510,N18511,N18512,N18513,N18514,N18515,N18516,N18517,N18518,
N18519,N18520,N18521,N18522,N18523,N18524,N18525,N18526,N18527,N18528,
N18529,N18530,N18531,N18532,N18533,N18534,N18535,N18536,N18537,N18538,
N18539,N18540,N18541,N18542,N18543,N18544,N18545,N18546,N18547,N18548,
N18549,N18550,N18551,N18552,N18553,N18554,N18555,N18556,N18557,N18558,
N18559,N18560,N18561,N18562,N18563,N18564,N18565,N18566,N18567,N18568,
N18569,N18570,N18571,N18572,N18573,N18574,N18575,N18576,N18577,N18578,
N18579,N18580,N18581,N18582,N18583,N18584,N18585,N18586,N18587,N18588,
N18589,N18590,N18591,N18592,N18593,N18594,N18595,N18596,N18597,N18598,
N18599,N18600,N18601,N18602,N18603,N18604,N18605,N18606,N18607,N18608,
N18609,N18610,N18611,N18612,N18613,N18614,N18615,N18616,N18617,N18618,
N18619,N18620,N18621,N18622,N18623,N18624,N18625,N18626,N18627,N18628,
N18629,N18630,N18631,N18632,N18633,N18634,N18635,N18636,N18637,N18638,
N18639,N18640,N18641,N18642,N18643,N18644,N18645,N18646,N18647,N18648,
N18649,N18650,N18651,N18652,N18653,N18654,N18655,N18656,N18657,N18658,
N18659,N18660,N18661,N18662,N18663,N18664,N18665,N18666,N18667,N18668,
N18669,N18670,N18671,N18672,N18673,N18674,N18675,N18676,N18677,N18678,
N18679,N18680,N18681,N18682,N18683,N18684,N18685,N18686,N18687,N18688,
N18689,N18690,N18691,N18692,N18693,N18694,N18695,N18696,N18697,N18698,
N18699,N18700,N18701,N18702,N18703,N18704,N18705,N18706,N18707,N18708,
N18709,N18710,N18711,N18712,N18713,N18714,N18715,N18716,N18717,N18718,
N18719,N18720,N18721,N18722,N18723,N18724,N18725,N18726,N18727,N18728,
N18729,N18730,N18731,N18732,N18733,N18734,N18735,N18736,N18737,N18738,
N18739,N18740,N18741,N18742,N18743,N18744,N18745,N18746,N18747,N18748,
N18749,N18750,N18751,N18752,N18753,N18754,N18755,N18756,N18757,N18758,
N18759,N18760,N18761,N18762,N18763,N18764,N18765,N18766,N18767,N18768,
N18769,N18770,N18771,N18772,N18773,N18774,N18775,N18776,N18777,N18778,
N18779,N18780,N18781,N18782,N18783,N18784,N18785,N18786,N18787,N18788,
N18789,N18790,N18791,N18792,N18793,N18794,N18795,N18796,N18797,N18798,
N18799,N18800,N18801,N18802,N18803,N18804,N18805,N18806,N18807,N18808,
N18809,N18810,N18811,N18812,N18813,N18814,N18815,N18816,N18817,N18818,
N18819,N18820,N18821,N18822,N18823,N18824,N18825,N18826,N18827,N18828,
N18829,N18830,N18831,N18832,N18833,N18834,N18835,N18836,N18837,N18838,
N18839,N18840,N18841,N18842,N18843,N18844,N18845,N18846,N18847,N18848,
N18849,N18850,N18851,N18852,N18853,N18854,N18855,N18856,N18857,N18858,
N18859,N18860,N18861,N18862,N18863,N18864,N18865,N18866,N18867,N18868,
N18869,N18870,N18871,N18872,N18873,N18874,N18875,N18876,N18877,N18878,
N18879,N18880,N18881,N18882,N18883,N18884,N18885,N18886,N18887,N18888,
N18889,N18890,N18891,N18892,N18893,N18894,N18895,N18896,N18897,N18898,
N18899,N18900,N18901,N18902,N18903,N18904,N18905,N18906,N18907,N18908,
N18909,N18910,N18911,N18912,N18913,N18914,N18915,N18916,N18917,N18918,
N18919,N18920,N18921,N18922,N18923,N18924,N18925,N18926,N18927,N18928,
N18929,N18930,N18931,N18932,N18933,N18934,N18935,N18936,N18937,N18938,
N18939,N18940,N18941,N18942,N18943,N18944,N18945,N18946,N18947,N18948,
N18949,N18950,N18951,N18952,N18953,N18954,N18955,N18956,N18957,N18958,
N18959,N18960,N18961,N18962,N18963,N18964,N18965,N18966,N18967,N18968,
N18969,N18970,N18971,N18972,N18973,N18974,N18975,N18976,N18977,N18978,
N18979,N18980,N18981,N18982,N18983,N18984,N18985,N18986,N18987,N18988,
N18989,N18990,N18991,N18992,N18993,N18994,N18995,N18996,N18997,N18998,
N18999,N19000,N19001,N19002,N19003,N19004,N19005,N19006,N19007,N19008,
N19009,N19010,N19011,N19012,N19013,N19014,N19015,N19016,N19017,N19018,
N19019,N19020,N19021,N19022,N19023,N19024,N19025,N19026,N19027,N19028,
N19029,N19030,N19031,N19032,N19033,N19034,N19035,N19036,N19037,N19038,
N19039,N19040,N19041,N19042,N19043,N19044,N19045,N19046,N19047,N19048,
N19049,N19050,N19051,N19052,N19053,N19054,N19055,N19056,N19057,N19058,
N19059,N19060,N19061,N19062,N19063,N19064,N19065,N19066,N19067,N19068,
N19069,N19070,N19071,N19072,N19073,N19074,N19075,N19076,N19077,N19078,
N19079,N19080,N19081,N19082,N19083,N19084,N19085,N19086,N19087,N19088,
N19089,N19090,N19091,N19092,N19093,N19094,N19095,N19096,N19097,N19098,
N19099,N19100,N19101,N19102,N19103,N19104,N19105,N19106,N19107,N19108,
N19109,N19110,N19111,N19112,N19113,N19114,N19115,N19116,N19117,N19118,
N19119,N19120,N19121,N19122,N19123,N19124,N19125,N19126,N19127,N19128,
N19129,N19130,N19131,N19132,N19133,N19134,N19135,N19136,N19137,N19138,
N19139,N19140,N19141,N19142,N19143,N19144,N19145,N19146,N19147,N19148,
N19149,N19150,N19151,N19152,N19153,N19154,N19155,N19156,N19157,N19158,
N19159,N19160,N19161,N19162,N19163,N19164,N19165,N19166,N19167,N19168,
N19169,N19170,N19171,N19172,N19173,N19174,N19175,N19176,N19177,N19178,
N19179,N19180,N19181,N19182,N19183,N19184,N19185,N19186,N19187,N19188,
N19189,N19190,N19191,N19192,N19193,N19194,N19195,N19196,N19197,N19198,
N19199,N19200,N19201,N19202,N19203,N19204,N19205,N19206,N19207,N19208,
N19209,N19210,N19211,N19212,N19213,N19214,N19215,N19216,N19217,N19218,
N19219,N19220,N19221,N19222,N19223,N19224,N19225,N19226,N19227,N19228,
N19229,N19230,N19231,N19232,N19233,N19234,N19235,N19236,N19237,N19238,
N19239,N19240,N19241,N19242,N19243,N19244,N19245,N19246,N19247,N19248,
N19249,N19250,N19251,N19252,N19253,N19254,N19255,N19256,N19257,N19258,
N19259,N19260,N19261,N19262,N19263,N19264,N19265,N19266,N19267,N19268,
N19269,N19270,N19271,N19272,N19273,N19274,N19275,N19276,N19277,N19278,
N19279,N19280,N19281,N19282,N19283,N19284,N19285,N19286,N19287,N19288,
N19289,N19290,N19291,N19292,N19293,N19294,N19295,N19296,N19297,N19298,
N19299,N19300,N19301,N19302,N19303,N19304,N19305,N19306,N19307,N19308,
N19309,N19310,N19311,N19312,N19313,N19314,N19315,N19316,N19317,N19318,
N19319,N19320,N19321,N19322,N19323,N19324,N19325,N19326,N19327,N19328,
N19329,N19330,N19331,N19332,N19333,N19334,N19335,N19336,N19337,N19338,
N19339,N19340,N19341,N19342,N19343,N19344,N19345,N19346,N19347,N19348,
N19349,N19350,N19351,N19352,N19353,N19354,N19355,N19356,N19357,N19358,
N19359,N19360,N19361,N19362,N19363,N19364,N19365,N19366,N19367,N19368,
N19369,N19370,N19371,N19372,N19373,N19374,N19375,N19376,N19377,N19378,
N19379,N19380,N19381,N19382,N19383,N19384,N19385,N19386,N19387,N19388,
N19389,N19390,N19391,N19392,N19393,N19394,N19395,N19396,N19397,N19398,
N19399,N19400,N19401,N19402,N19403,N19404,N19405,N19406,N19407,N19408,
N19409,N19410,N19411,N19412,N19413,N19414,N19415,N19416,N19417,N19418,
N19419,N19420,N19421,N19422,N19423,N19424,N19425,N19426,N19427,N19428,
N19429,N19430,N19431,N19432,N19433,N19434,N19435,N19436,N19437,N19438,
N19439,N19440,N19441,N19442,N19443,N19444,N19445,N19446,N19447,N19448,
N19449,N19450,N19451,N19452,N19453,N19454,N19455,N19456,N19457,N19458,
N19459,N19460,N19461,N19462,N19463,N19464,N19465,N19466,N19467,N19468,
N19469,N19470,N19471,N19472,N19473,N19474,N19475,N19476,N19477,N19478,
N19479,N19480,N19481,N19482,N19483,N19484,N19485,N19486,N19487,N19488,
N19489,N19490,N19491,N19492,N19493,N19494,N19495,N19496,N19497,N19498,
N19499,N19500,N19501,N19502,N19503,N19504,N19505,N19506,N19507,N19508,
N19509,N19510,N19511,N19512,N19513,N19514,N19515,N19516,N19517,N19518,
N19519,N19520,N19521,N19522,N19523,N19524,N19525,N19526,N19527,N19528,
N19529,N19530,N19531,N19532,N19533,N19534,N19535,N19536,N19537,N19538,
N19539,N19540,N19541,N19542,N19543,N19544,N19545,N19546,N19547,N19548,
N19549,N19550,N19551,N19552,N19553,N19554,N19555,N19556,N19557,N19558,
N19559,N19560,N19561,N19562,N19563,N19564,N19565,N19566,N19567,N19568,
N19569,N19570,N19571,N19572,N19573,N19574,N19575,N19576,N19577,N19578,
N19579,N19580,N19581,N19582,N19583,N19584,N19585,N19586,N19587,N19588,
N19589,N19590,N19591,N19592,N19593,N19594,N19595,N19596,N19597,N19598,
N19599,N19600,N19601,N19602,N19603,N19604,N19605,N19606,N19607,N19608,
N19609,N19610,N19611,N19612,N19613,N19614,N19615,N19616,N19617,N19618,
N19619,N19620,N19621,N19622,N19623,N19624,N19625,N19626,N19627,N19628,
N19629,N19630,N19631,N19632,N19633,N19634,N19635,N19636,N19637,N19638,
N19639,N19640,N19641,N19642,N19643,N19644,N19645,N19646,N19647,N19648,
N19649,N19650,N19651,N19652,N19653,N19654,N19655,N19656,N19657,N19658,
N19659,N19660,N19661,N19662,N19663,N19664,N19665,N19666,N19667,N19668,
N19669,N19670,N19671,N19672,N19673,N19674,N19675,N19676,N19677,N19678,
N19679,N19680,N19681,N19682,N19683,N19684,N19685,N19686,N19687,N19688,
N19689,N19690,N19691,N19692,N19693,N19694,N19695,N19696,N19697,N19698,
N19699,N19700,N19701,N19702,N19703,N19704,N19705,N19706,N19707,N19708,
N19709,N19710,N19711,N19712,N19713,N19714,N19715,N19716,N19717,N19718,
N19719,N19720,N19721,N19722,N19723,N19724,N19725,N19726,N19727,N19728,
N19729,N19730,N19731,N19732,N19733,N19734,N19735,N19736,N19737,N19738,
N19739,N19740,N19741,N19742,N19743,N19744,N19745,N19746,N19747,N19748,
N19749,N19750,N19751,N19752,N19753,N19754,N19755,N19756,N19757,N19758,
N19759,N19760,N19761,N19762,N19763,N19764,N19765,N19766,N19767,N19768,
N19769,N19770,N19771,N19772,N19773,N19774,N19775,N19776,N19777,N19778,
N19779,N19780,N19781,N19782,N19783,N19784,N19785,N19786,N19787,N19788,
N19789,N19790,N19791,N19792,N19793,N19794,N19795,N19796,N19797,N19798,
N19799,N19800,N19801,N19802,N19803,N19804,N19805,N19806,N19807,N19808,
N19809,N19810,N19811,N19812,N19813,N19814,N19815,N19816,N19817,N19818,
N19819,N19820,N19821,N19822,N19823,N19824,N19825,N19826,N19827,N19828,
N19829,N19830,N19831,N19832,N19833,N19834,N19835,N19836,N19837,N19838,
N19839,N19840,N19841,N19842,N19843,N19844,N19845,N19846,N19847,N19848,
N19849,N19850,N19851,N19852,N19853,N19854,N19855,N19856,N19857,N19858,
N19859,N19860,N19861,N19862,N19863,N19864,N19865,N19866,N19867,N19868,
N19869,N19870,N19871,N19872,N19873,N19874,N19875,N19876,N19877,N19878,
N19879,N19880,N19881,N19882,N19883,N19884,N19885,N19886,N19887,N19888,
N19889,N19890,N19891,N19892,N19893,N19894,N19895,N19896,N19897,N19898,
N19899,N19900,N19901,N19902,N19903,N19904,N19905,N19906,N19907,N19908,
N19909,N19910,N19911,N19912,N19913,N19914,N19915,N19916,N19917,N19918,
N19919,N19920,N19921,N19922,N19923,N19924,N19925,N19926,N19927,N19928,
N19929,N19930,N19931,N19932,N19933,N19934,N19935,N19936,N19937,N19938,
N19939,N19940,N19941,N19942,N19943,N19944,N19945,N19946,N19947,N19948,
N19949,N19950,N19951,N19952,N19953,N19954,N19955,N19956,N19957,N19958,
N19959,N19960,N19961,N19962,N19963,N19964,N19965,N19966,N19967,N19968,
N19969,N19970,N19971,N19972,N19973,N19974,N19975,N19976,N19977,N19978,
N19979,N19980,N19981,N19982,N19983,N19984,N19985,N19986,N19987,N19988,
N19989,N19990,N19991,N19992,N19993,N19994,N19995,N19996,N19997,N19998,
N19999,N20000,N20001,N20002,N20003,N20004,N20005,N20006,N20007,N20008,
N20009,N20010,N20011,N20012,N20013,N20014,N20015,N20016,N20017,N20018,
N20019,N20020,N20021,N20022,N20023,N20024,N20025,N20026,N20027,N20028,
N20029,N20030,N20031,N20032,N20033,N20034,N20035,N20036,N20037,N20038,
N20039,N20040,N20041,N20042,N20043,N20044,N20045,N20046,N20047,N20048,
N20049,N20050,N20051,N20052,N20053,N20054,N20055,N20056,N20057,N20058,
N20059,N20060,N20061,N20062,N20063,N20064,N20065,N20066,N20067,N20068,
N20069,N20070,N20071,N20072,N20073,N20074,N20075,N20076,N20077,N20078,
N20079,N20080,N20081,N20082,N20083,N20084,N20085,N20086,N20087,N20088,
N20089,N20090,N20091,N20092,N20093,N20094,N20095,N20096,N20097,N20098,
N20099,N20100,N20101,N20102,N20103,N20104,N20105,N20106,N20107,N20108,
N20109,N20110,N20111,N20112,N20113,N20114,N20115,N20116,N20117,N20118,
N20119,N20120,N20121,N20122,N20123,N20124,N20125,N20126,N20127,N20128,
N20129,N20130,N20131,N20132,N20133,N20134,N20135,N20136,N20137,N20138,
N20139,N20140,N20141,N20142,N20143,N20144,N20145,N20146,N20147,N20148,
N20149,N20150,N20151,N20152,N20153,N20154,N20155,N20156,N20157,N20158,
N20159,N20160,N20161,N20162,N20163,N20164,N20165,N20166,N20167,N20168,
N20169,N20170,N20171,N20172,N20173,N20174,N20175,N20176,N20177,N20178,
N20179,N20180,N20181,N20182,N20183,N20184,N20185,N20186,N20187,N20188,
N20189,N20190,N20191,N20192,N20193,N20194,N20195,N20196,N20197,N20198,
N20199,N20200,N20201,N20202,N20203,N20204,N20205,N20206,N20207,N20208,
N20209,N20210,N20211,N20212,N20213,N20214,N20215,N20216,N20217,N20218,
N20219,N20220,N20221,N20222,N20223,N20224,N20225,N20226,N20227,N20228,
N20229,N20230,N20231,N20232,N20233,N20234,N20235,N20236,N20237,N20238,
N20239,N20240,N20241,N20242,N20243,N20244,N20245,N20246,N20247,N20248,
N20249,N20250,N20251,N20252,N20253,N20254,N20255,N20256,N20257,N20258,
N20259,N20260,N20261,N20262,N20263,N20264,N20265,N20266,N20267,N20268,
N20269,N20270,N20271,N20272,N20273,N20274,N20275,N20276,N20277,N20278,
N20279,N20280,N20281,N20282,N20283,N20284,N20285,N20286,N20287,N20288,
N20289,N20290,N20291,N20292,N20293,N20294,N20295,N20296,N20297,N20298,
N20299,N20300,N20301,N20302,N20303,N20304,N20305,N20306,N20307,N20308,
N20309,N20310,N20311,N20312,N20313,N20314,N20315,N20316,N20317,N20318,
N20319,N20320,N20321,N20322,N20323,N20324,N20325,N20326,N20327,N20328,
N20329,N20330,N20331,N20332,N20333,N20334,N20335,N20336,N20337,N20338,
N20339,N20340,N20341,N20342,N20343,N20344,N20345,N20346,N20347,N20348,
N20349,N20350,N20351,N20352,N20353,N20354,N20355,N20356,N20357,N20358,
N20359,N20360,N20361,N20362,N20363,N20364,N20365,N20366,N20367,N20368,
N20369,N20370,N20371,N20372,N20373,N20374,N20375,N20376,N20377,N20378,
N20379,N20380,N20381,N20382,N20383,N20384,N20385,N20386,N20387,N20388,
N20389,N20390,N20391,N20392,N20393,N20394,N20395,N20396,N20397,N20398,
N20399,N20400,N20401,N20402,N20403,N20404,N20405,N20406,N20407,N20408,
N20409,N20410,N20411,N20412,N20413,N20414,N20415,N20416,N20417,N20418,
N20419,N20420,N20421,N20422,N20423,N20424,N20425,N20426,N20427,N20428,
N20429,N20430,N20431,N20432,N20433,N20434,N20435,N20436,N20437,N20438,
N20439,N20440,N20441,N20442,N20443,N20444,N20445,N20446,N20447,N20448,
N20449,N20450,N20451,N20452,N20453,N20454,N20455,N20456,N20457,N20458,
N20459,N20460,N20461,N20462,N20463,N20464,N20465,N20466,N20467,N20468,
N20469,N20470,N20471,N20472,N20473,N20474,N20475,N20476,N20477,N20478,
N20479,N20480,N20481,N20482,N20483,N20484,N20485,N20486,N20487,N20488,
N20489,N20490,N20491,N20492,N20493,N20494,N20495,N20496,N20497,N20498,
N20499,N20500,N20501,N20502,N20503,N20504,N20505,N20506,N20507,N20508,
N20509,N20510,N20511,N20512,N20513,N20514,N20515,N20516,N20517,N20518,
N20519,N20520,N20521,N20522,N20523,N20524,N20525,N20526,N20527,N20528,
N20529,N20530,N20531,N20532,N20533,N20534,N20535,N20536,N20537,N20538,
N20539,N20540,N20541,N20542,N20543,N20544,N20545,N20546,N20547,N20548,
N20549,N20550,N20551,N20552,N20553,N20554,N20555,N20556,N20557,N20558,
N20559,N20560,N20561,N20562,N20563,N20564,N20565,N20566,N20567,N20568,
N20569,N20570,N20571,N20572,N20573,N20574,N20575,N20576,N20577,N20578,
N20579,N20580,N20581,N20582,N20583,N20584,N20585,N20586,N20587,N20588,
N20589,N20590,N20591,N20592,N20593,N20594,N20595,N20596,N20597,N20598,
N20599,N20600,N20601,N20602,N20603,N20604,N20605,N20606,N20607,N20608,
N20609,N20610,N20611,N20612,N20613,N20614,N20615,N20616,N20617,N20618,
N20619,N20620,N20621,N20622,N20623,N20624,N20625,N20626,N20627,N20628,
N20629,N20630,N20631,N20632,N20633,N20634,N20635,N20636,N20637,N20638,
N20639,N20640,N20641,N20642,N20643,N20644,N20645,N20646,N20647,N20648,
N20649,N20650,N20651,N20652,N20653,N20654,N20655,N20656,N20657,N20658,
N20659,N20660,N20661,N20662,N20663,N20664,N20665,N20666,N20667,N20668,
N20669,N20670,N20671,N20672,N20673,N20674,N20675,N20676,N20677,N20678,
N20679,N20680,N20681,N20682,N20683,N20684,N20685,N20686,N20687,N20688,
N20689,N20690,N20691,N20692,N20693,N20694,N20695,N20696,N20697,N20698,
N20699,N20700,N20701,N20702,N20703,N20704,N20705,N20706,N20707,N20708,
N20709,N20710,N20711,N20712,N20713,N20714,N20715,N20716,N20717,N20718,
N20719,N20720,N20721,N20722,N20723,N20724,N20725,N20726,N20727,N20728,
N20729,N20730,N20731,N20732,N20733,N20734,N20735,N20736,N20737,N20738,
N20739,N20740,N20741,N20742,N20743,N20744,N20745,N20746,N20747,N20748,
N20749,N20750,N20751,N20752,N20753,N20754,N20755,N20756,N20757,N20758,
N20759,N20760,N20761,N20762,N20763,N20764,N20765,N20766,N20767,N20768,
N20769,N20770,N20771,N20772,N20773,N20774,N20775,N20776,N20777,N20778,
N20779,N20780,N20781,N20782,N20783,N20784,N20785,N20786,N20787,N20788,
N20789,N20790,N20791,N20792,N20793,N20794,N20795,N20796,N20797,N20798,
N20799,N20800,N20801,N20802,N20803,N20804,N20805,N20806,N20807,N20808,
N20809,N20810,N20811,N20812,N20813,N20814,N20815,N20816,N20817,N20818,
N20819,N20820,N20821,N20822,N20823,N20824,N20825,N20826,N20827,N20828,
N20829,N20830,N20831,N20832,N20833,N20834,N20835,N20836,N20837,N20838,
N20839,N20840,N20841,N20842,N20843,N20844,N20845,N20846,N20847,N20848,
N20849,N20850,N20851,N20852,N20853,N20854,N20855,N20856,N20857,N20858,
N20859,N20860,N20861,N20862,N20863,N20864,N20865,N20866,N20867,N20868,
N20869,N20870,N20871,N20872,N20873,N20874,N20875,N20876,N20877,N20878,
N20879,N20880,N20881,N20882,N20883,N20884,N20885,N20886,N20887,N20888,
N20889,N20890,N20891,N20892,N20893,N20894,N20895,N20896,N20897,N20898,
N20899,N20900,N20901,N20902,N20903,N20904,N20905,N20906,N20907,N20908,
N20909,N20910,N20911,N20912,N20913,N20914,N20915,N20916,N20917,N20918,
N20919,N20920,N20921,N20922,N20923,N20924,N20925,N20926,N20927,N20928,
N20929,N20930,N20931,N20932,N20933,N20934,N20935,N20936,N20937,N20938,
N20939,N20940,N20941,N20942,N20943,N20944,N20945,N20946,N20947,N20948,
N20949,N20950,N20951,N20952,N20953,N20954,N20955,N20956,N20957,N20958,
N20959,N20960,N20961,N20962,N20963,N20964,N20965,N20966,N20967,N20968,
N20969,N20970,N20971,N20972,N20973,N20974,N20975,N20976,N20977,N20978,
N20979,N20980,N20981,N20982,N20983,N20984,N20985,N20986,N20987,N20988,
N20989,N20990,N20991,N20992,N20993,N20994,N20995,N20996,N20997,N20998,
N20999,N21000,N21001,N21002,N21003,N21004,N21005,N21006,N21007,N21008,
N21009,N21010,N21011,N21012,N21013,N21014,N21015,N21016,N21017,N21018,
N21019,N21020,N21021,N21022,N21023,N21024,N21025,N21026,N21027,N21028,
N21029,N21030,N21031,N21032,N21033,N21034,N21035,N21036,N21037,N21038,
N21039,N21040,N21041,N21042,N21043,N21044,N21045,N21046,N21047,N21048,
N21049,N21050,N21051,N21052,N21053,N21054,N21055,N21056,N21057,N21058,
N21059,N21060,N21061,N21062,N21063,N21064,N21065,N21066,N21067,N21068,
N21069,N21070,N21071,N21072,N21073,N21074,N21075,N21076,N21077,N21078,
N21079,N21080,N21081,N21082,N21083,N21084,N21085,N21086,N21087,N21088,
N21089,N21090,N21091,N21092,N21093,N21094,N21095,N21096,N21097,N21098,
N21099,N21100,N21101,N21102,N21103,N21104,N21105,N21106,N21107,N21108,
N21109,N21110,N21111,N21112,N21113,N21114,N21115,N21116,N21117,N21118,
N21119,N21120,N21121,N21122,N21123,N21124,N21125,N21126,N21127,N21128,
N21129,N21130,N21131,N21132,N21133,N21134,N21135,N21136,N21137,N21138,
N21139,N21140,N21141,N21142,N21143,N21144,N21145,N21146,N21147,N21148,
N21149,N21150,N21151,N21152,N21153,N21154,N21155,N21156,N21157,N21158,
N21159,N21160,N21161,N21162,N21163,N21164,N21165,N21166,N21167,N21168,
N21169,N21170,N21171,N21172,N21173,N21174,N21175,N21176,N21177,N21178,
N21179,N21180,N21181,N21182,N21183,N21184,N21185,N21186,N21187,N21188,
N21189,N21190,N21191,N21192,N21193,N21194,N21195,N21196,N21197,N21198,
N21199,N21200,N21201,N21202,N21203,N21204,N21205,N21206,N21207,N21208,
N21209,N21210,N21211,N21212,N21213,N21214,N21215,N21216,N21217,N21218,
N21219,N21220,N21221,N21222,N21223,N21224,N21225,N21226,N21227,N21228,
N21229,N21230,N21231,N21232,N21233,N21234,N21235,N21236,N21237,N21238,
N21239,N21240,N21241,N21242,N21243,N21244,N21245,N21246,N21247,N21248,
N21249,N21250,N21251,N21252,N21253,N21254,N21255,N21256,N21257,N21258,
N21259,N21260,N21261,N21262,N21263,N21264,N21265,N21266,N21267,N21268,
N21269,N21270,N21271,N21272,N21273,N21274,N21275,N21276,N21277,N21278,
N21279,N21280,N21281,N21282,N21283,N21284,N21285,N21286,N21287,N21288,
N21289,N21290,N21291,N21292,N21293,N21294,N21295,N21296,N21297,N21298,
N21299,N21300,N21301,N21302,N21303,N21304,N21305,N21306,N21307,N21308,
N21309,N21310,N21311,N21312,N21313,N21314,N21315,N21316,N21317,N21318,
N21319,N21320,N21321,N21322,N21323,N21324,N21325,N21326,N21327,N21328,
N21329,N21330,N21331,N21332,N21333,N21334,N21335,N21336,N21337,N21338,
N21339,N21340,N21341,N21342,N21343,N21344,N21345,N21346,N21347,N21348,
N21349,N21350,N21351,N21352,N21353,N21354,N21355,N21356,N21357,N21358,
N21359,N21360,N21361,N21362,N21363,N21364,N21365,N21366,N21367,N21368,
N21369,N21370,N21371,N21372,N21373,N21374,N21375,N21376,N21377,N21378,
N21379,N21380,N21381,N21382,N21383,N21384,N21385,N21386,N21387,N21388,
N21389,N21390,N21391,N21392,N21393,N21394,N21395,N21396,N21397,N21398,
N21399,N21400,N21401,N21402,N21403,N21404,N21405,N21406,N21407,N21408,
N21409,N21410,N21411,N21412,N21413,N21414,N21415,N21416,N21417,N21418,
N21419,N21420,N21421,N21422,N21423,N21424,N21425,N21426,N21427,N21428,
N21429,N21430,N21431,N21432,N21433,N21434,N21435,N21436,N21437,N21438,
N21439,N21440,N21441,N21442,N21443,N21444,N21445,N21446,N21447,N21448,
N21449,N21450,N21451,N21452,N21453,N21454,N21455,N21456,N21457,N21458,
N21459,N21460,N21461,N21462,N21463,N21464,N21465,N21466,N21467,N21468,
N21469,N21470,N21471,N21472,N21473,N21474,N21475,N21476,N21477,N21478,
N21479,N21480,N21481,N21482,N21483,N21484,N21485,N21486,N21487,N21488,
N21489,N21490,N21491,N21492,N21493,N21494,N21495,N21496,N21497,N21498,
N21499,N21500,N21501,N21502,N21503,N21504,N21505,N21506,N21507,N21508,
N21509,N21510,N21511,N21512,N21513,N21514,N21515,N21516,N21517,N21518,
N21519,N21520,N21521,N21522,N21523,N21524,N21525,N21526,N21527,N21528,
N21529,N21530,N21531,N21532,N21533,N21534,N21535,N21536,N21537,N21538,
N21539,N21540,N21541,N21542,N21543,N21544,N21545,N21546,N21547,N21548,
N21549,N21550,N21551,N21552,N21553,N21554,N21555,N21556,N21557,N21558,
N21559,N21560,N21561,N21562,N21563,N21564,N21565,N21566,N21567,N21568,
N21569,N21570,N21571,N21572,N21573,N21574,N21575,N21576,N21577,N21578,
N21579,N21580,N21581,N21582,N21583,N21584,N21585,N21586,N21587,N21588,
N21589,N21590,N21591,N21592,N21593,N21594,N21595,N21596,N21597,N21598,
N21599,N21600,N21601,N21602,N21603,N21604,N21605,N21606,N21607,N21608,
N21609,N21610,N21611,N21612,N21613,N21614,N21615,N21616,N21617,N21618,
N21619,N21620,N21621,N21622,N21623,N21624,N21625,N21626,N21627,N21628,
N21629,N21630,N21631,N21632,N21633,N21634,N21635,N21636,N21637,N21638,
N21639,N21640,N21641,N21642,N21643,N21644,N21645,N21646,N21647,N21648,
N21649,N21650,N21651,N21652,N21653,N21654,N21655,N21656,N21657,N21658,
N21659,N21660,N21661,N21662,N21663,N21664,N21665,N21666,N21667,N21668,
N21669,N21670,N21671,N21672,N21673,N21674,N21675,N21676,N21677,N21678,
N21679,N21680,N21681,N21682,N21683,N21684,N21685,N21686,N21687,N21688,
N21689,N21690,N21691,N21692,N21693,N21694,N21695,N21696,N21697,N21698,
N21699,N21700,N21701,N21702,N21703,N21704,N21705,N21706,N21707,N21708,
N21709,N21710,N21711,N21712,N21713,N21714,N21715,N21716,N21717,N21718,
N21719,N21720,N21721,N21722,N21723,N21724,N21725,N21726,N21727,N21728,
N21729,N21730,N21731,N21732,N21733,N21734,N21735,N21736,N21737,N21738,
N21739,N21740,N21741,N21742,N21743,N21744,N21745,N21746,N21747,N21748,
N21749,N21750,N21751,N21752,N21753,N21754,N21755,N21756,N21757,N21758,
N21759,N21760,N21761,N21762,N21763,N21764,N21765,N21766,N21767,N21768,
N21769,N21770,N21771,N21772,N21773,N21774,N21775,N21776,N21777,N21778,
N21779,N21780,N21781,N21782,N21783,N21784,N21785,N21786,N21787,N21788,
N21789,N21790,N21791,N21792,N21793,N21794,N21795,N21796,N21797,N21798,
N21799,N21800,N21801,N21802,N21803,N21804,N21805,N21806,N21807,N21808,
N21809,N21810,N21811,N21812,N21813,N21814,N21815,N21816,N21817,N21818,
N21819,N21820,N21821,N21822,N21823,N21824,N21825,N21826,N21827,N21828,
N21829,N21830,N21831,N21832,N21833,N21834,N21835,N21836,N21837,N21838,
N21839,N21840,N21841,N21842,N21843,N21844,N21845,N21846,N21847,N21848,
N21849,N21850,N21851,N21852,N21853,N21854,N21855,N21856,N21857,N21858,
N21859,N21860,N21861,N21862,N21863,N21864,N21865,N21866,N21867,N21868,
N21869,N21870,N21871,N21872,N21873,N21874,N21875,N21876,N21877,N21878,
N21879,N21880,N21881,N21882,N21883,N21884,N21885,N21886,N21887,N21888,
N21889,N21890,N21891,N21892,N21893,N21894,N21895,N21896,N21897,N21898,
N21899,N21900,N21901,N21902,N21903,N21904,N21905,N21906,N21907,N21908,
N21909,N21910,N21911,N21912,N21913,N21914,N21915,N21916,N21917,N21918,
N21919,N21920,N21921,N21922,N21923,N21924,N21925,N21926,N21927,N21928,
N21929,N21930,N21931,N21932,N21933,N21934,N21935,N21936,N21937,N21938,
N21939,N21940,N21941,N21942,N21943,N21944,N21945,N21946,N21947,N21948,
N21949,N21950,N21951,N21952,N21953,N21954,N21955,N21956,N21957,N21958,
N21959,N21960,N21961,N21962,N21963,N21964,N21965,N21966,N21967,N21968,
N21969,N21970,N21971,N21972,N21973,N21974,N21975,N21976,N21977,N21978,
N21979,N21980,N21981,N21982,N21983,N21984,N21985,N21986,N21987,N21988,
N21989,N21990,N21991,N21992,N21993,N21994,N21995,N21996,N21997,N21998,
N21999,N22000,N22001,N22002,N22003,N22004,N22005,N22006,N22007,N22008,
N22009,N22010,N22011,N22012,N22013,N22014,N22015,N22016,N22017,N22018,
N22019,N22020,N22021,N22022,N22023,N22024,N22025,N22026,N22027,N22028,
N22029,N22030,N22031,N22032,N22033,N22034,N22035,N22036,N22037,N22038,
N22039,N22040,N22041,N22042,N22043,N22044,N22045,N22046,N22047,N22048,
N22049,N22050,N22051,N22052,N22053,N22054,N22055,N22056,N22057,N22058,
N22059,N22060,N22061,N22062,N22063,N22064,N22065,N22066,N22067,N22068,
N22069,N22070,N22071,N22072,N22073,N22074,N22075,N22076,N22077,N22078,
N22079,N22080,N22081,N22082,N22083,N22084,N22085,N22086,N22087,N22088,
N22089,N22090,N22091,N22092,N22093,N22094,N22095,N22096,N22097,N22098,
N22099,N22100,N22101,N22102,N22103,N22104,N22105,N22106,N22107,N22108,
N22109,N22110,N22111,N22112,N22113,N22114,N22115,N22116,N22117,N22118,
N22119,N22120,N22121,N22122,N22123,N22124,N22125,N22126,N22127,N22128,
N22129,N22130,N22131,N22132,N22133,N22134,N22135,N22136,N22137,N22138,
N22139,N22140,N22141,N22142,N22143,N22144,N22145,N22146,N22147,N22148,
N22149,N22150,N22151,N22152,N22153,N22154,N22155,N22156,N22157,N22158,
N22159,N22160,N22161,N22162,N22163,N22164,N22165,N22166,N22167,N22168,
N22169,N22170,N22171,N22172,N22173,N22174,N22175,N22176,N22177,N22178,
N22179,N22180,N22181,N22182,N22183,N22184,N22185,N22186,N22187,N22188,
N22189,N22190,N22191,N22192,N22193,N22194,N22195,N22196,N22197,N22198,
N22199,N22200,N22201,N22202,N22203,N22204,N22205,N22206,N22207,N22208,
N22209,N22210,N22211,N22212,N22213,N22214,N22215,N22216,N22217,N22218,
N22219,N22220,N22221,N22222,N22223,N22224,N22225,N22226,N22227,N22228,
N22229,N22230,N22231,N22232,N22233,N22234,N22235,N22236,N22237,N22238,
N22239,N22240,N22241,N22242,N22243,N22244,N22245,N22246,N22247,N22248,
N22249,N22250,N22251,N22252,N22253,N22254,N22255,N22256,N22257,N22258,
N22259,N22260,N22261,N22262,N22263,N22264,N22265,N22266,N22267,N22268,
N22269,N22270,N22271,N22272,N22273,N22274,N22275,N22276,N22277,N22278,
N22279,N22280,N22281,N22282,N22283,N22284,N22285,N22286,N22287,N22288,
N22289,N22290,N22291,N22292,N22293,N22294,N22295,N22296,N22297,N22298,
N22299,N22300,N22301,N22302,N22303,N22304,N22305,N22306,N22307,N22308,
N22309,N22310,N22311,N22312,N22313,N22314,N22315,N22316,N22317,N22318,
N22319,N22320,N22321,N22322,N22323,N22324,N22325,N22326,N22327,N22328,
N22329,N22330,N22331,N22332,N22333,N22334,N22335,N22336,N22337,N22338,
N22339,N22340,N22341,N22342,N22343,N22344,N22345,N22346,N22347,N22348,
N22349,N22350,N22351,N22352,N22353,N22354,N22355,N22356,N22357,N22358,
N22359,N22360,N22361,N22362,N22363,N22364,N22365,N22366,N22367,N22368,
N22369,N22370,N22371,N22372,N22373,N22374,N22375,N22376,N22377,N22378,
N22379,N22380,N22381,N22382,N22383,N22384,N22385,N22386,N22387,N22388,
N22389,N22390,N22391,N22392,N22393,N22394,N22395,N22396,N22397,N22398,
N22399,N22400,N22401,N22402,N22403,N22404,N22405,N22406,N22407,N22408,
N22409,N22410,N22411,N22412,N22413,N22414,N22415,N22416,N22417,N22418,
N22419,N22420,N22421,N22422,N22423,N22424,N22425,N22426,N22427,N22428,
N22429,N22430,N22431,N22432,N22433,N22434,N22435,N22436,N22437,N22438,
N22439,N22440,N22441,N22442,N22443,N22444,N22445,N22446,N22447,N22448,
N22449,N22450,N22451,N22452,N22453,N22454,N22455,N22456,N22457,N22458,
N22459,N22460,N22461,N22462,N22463,N22464,N22465,N22466,N22467,N22468,
N22469,N22470,N22471,N22472,N22473,N22474,N22475,N22476,N22477,N22478,
N22479,N22480,N22481,N22482,N22483,N22484,N22485,N22486,N22487,N22488,
N22489,N22490,N22491,N22492,N22493,N22494,N22495,N22496,N22497,N22498,
N22499,N22500,N22501,N22502,N22503,N22504,N22505,N22506,N22507,N22508,
N22509,N22510,N22511,N22512,N22513,N22514,N22515,N22516,N22517,N22518,
N22519,N22520,N22521,N22522,N22523,N22524,N22525,N22526,N22527,N22528,
N22529,N22530,N22531,N22532,N22533,N22534,N22535,N22536,N22537,N22538,
N22539,N22540,N22541,N22542,N22543,N22544,N22545,N22546,N22547,N22548,
N22549,N22550,N22551,N22552,N22553,N22554,N22555,N22556,N22557,N22558,
N22559,N22560,N22561,N22562,N22563,N22564,N22565,N22566,N22567,N22568,
N22569,N22570,N22571,N22572,N22573,N22574,N22575,N22576,N22577,N22578,
N22579,N22580,N22581,N22582,N22583,N22584,N22585,N22586,N22587,N22588,
N22589,N22590,N22591,N22592,N22593,N22594,N22595,N22596,N22597,N22598,
N22599,N22600,N22601,N22602,N22603,N22604,N22605,N22606,N22607,N22608,
N22609,N22610,N22611,N22612,N22613,N22614,N22615,N22616,N22617,N22618,
N22619,N22620,N22621,N22622,N22623,N22624,N22625,N22626,N22627,N22628,
N22629,N22630,N22631,N22632,N22633,N22634,N22635,N22636,N22637,N22638,
N22639,N22640,N22641,N22642,N22643,N22644,N22645,N22646,N22647,N22648,
N22649,N22650,N22651,N22652,N22653,N22654,N22655,N22656,N22657,N22658,
N22659,N22660,N22661,N22662,N22663,N22664,N22665,N22666,N22667,N22668,
N22669,N22670,N22671,N22672,N22673,N22674,N22675,N22676,N22677,N22678,
N22679,N22680,N22681,N22682,N22683,N22684,N22685,N22686,N22687,N22688,
N22689,N22690,N22691,N22692,N22693,N22694,N22695,N22696,N22697,N22698,
N22699,N22700,N22701,N22702,N22703,N22704,N22705,N22706,N22707,N22708,
N22709,N22710,N22711,N22712,N22713,N22714,N22715,N22716,N22717,N22718,
N22719,N22720,N22721,N22722,N22723,N22724,N22725,N22726,N22727,N22728,
N22729,N22730,N22731,N22732,N22733,N22734,N22735,N22736,N22737,N22738,
N22739,N22740,N22741,N22742,N22743,N22744,N22745,N22746,N22747,N22748,
N22749,N22750,N22751,N22752,N22753,N22754,N22755,N22756,N22757,N22758,
N22759,N22760,N22761,N22762,N22763,N22764,N22765,N22766,N22767,N22768,
N22769,N22770,N22771,N22772,N22773,N22774,N22775,N22776,N22777,N22778,
N22779,N22780,N22781,N22782,N22783,N22784,N22785,N22786,N22787,N22788,
N22789,N22790,N22791,N22792,N22793,N22794,N22795,N22796,N22797,N22798,
N22799,N22800,N22801,N22802,N22803,N22804,N22805,N22806,N22807,N22808,
N22809,N22810,N22811,N22812,N22813,N22814,N22815,N22816,N22817,N22818,
N22819,N22820,N22821,N22822,N22823,N22824,N22825,N22826,N22827,N22828,
N22829,N22830,N22831,N22832,N22833,N22834,N22835,N22836,N22837,N22838,
N22839,N22840,N22841,N22842,N22843,N22844,N22845,N22846,N22847,N22848,
N22849,N22850,N22851,N22852,N22853,N22854,N22855,N22856,N22857,N22858,
N22859,N22860,N22861,N22862,N22863,N22864,N22865,N22866,N22867,N22868,
N22869,N22870,N22871,N22872,N22873,N22874,N22875,N22876,N22877,N22878,
N22879,N22880,N22881,N22882,N22883,N22884,N22885,N22886,N22887,N22888,
N22889,N22890,N22891,N22892,N22893,N22894,N22895,N22896,N22897,N22898,
N22899,N22900,N22901,N22902,N22903,N22904,N22905,N22906,N22907,N22908,
N22909,N22910,N22911,N22912,N22913,N22914,N22915,N22916,N22917,N22918,
N22919,N22920,N22921,N22922,N22923,N22924,N22925,N22926,N22927,N22928,
N22929,N22930,N22931,N22932,N22933,N22934,N22935,N22936,N22937,N22938,
N22939,N22940,N22941,N22942,N22943,N22944,N22945,N22946,N22947,N22948,
N22949,N22950,N22951,N22952,N22953,N22954,N22955,N22956,N22957,N22958,
N22959,N22960,N22961,N22962,N22963,N22964,N22965,N22966,N22967,N22968,
N22969,N22970,N22971,N22972,N22973,N22974,N22975,N22976,N22977,N22978,
N22979,N22980,N22981,N22982,N22983,N22984,N22985,N22986,N22987,N22988,
N22989,N22990,N22991,N22992,N22993,N22994,N22995,N22996,N22997,N22998,
N22999,N23000,N23001,N23002,N23003,N23004,N23005,N23006,N23007,N23008,
N23009,N23010,N23011,N23012,N23013,N23014,N23015,N23016,N23017,N23018,
N23019,N23020,N23021,N23022,N23023,N23024,N23025,N23026,N23027,N23028,
N23029,N23030,N23031,N23032,N23033,N23034,N23035,N23036,N23037,N23038,
N23039,N23040,N23041,N23042,N23043,N23044,N23045,N23046,N23047,N23048,
N23049,N23050,N23051,N23052,N23053,N23054,N23055,N23056,N23057,N23058,
N23059,N23060,N23061,N23062,N23063,N23064,N23065,N23066,N23067,N23068,
N23069,N23070,N23071,N23072,N23073,N23074,N23075,N23076,N23077,N23078,
N23079,N23080,N23081,N23082,N23083,N23084,N23085,N23086,N23087,N23088,
N23089,N23090,N23091,N23092,N23093,N23094,N23095,N23096,N23097,N23098,
N23099,N23100,N23101,N23102,N23103,N23104,N23105,N23106,N23107,N23108,
N23109,N23110,N23111,N23112,N23113,N23114,N23115,N23116,N23117,N23118,
N23119,N23120,N23121,N23122,N23123,N23124,N23125,N23126,N23127,N23128,
N23129,N23130,N23131,N23132,N23133,N23134,N23135,N23136,N23137,N23138,
N23139,N23140,N23141,N23142,N23143,N23144,N23145,N23146,N23147,N23148,
N23149,N23150,N23151,N23152,N23153,N23154,N23155,N23156,N23157,N23158,
N23159,N23160,N23161,N23162,N23163,N23164,N23165,N23166,N23167,N23168,
N23169,N23170,N23171,N23172,N23173,N23174,N23175,N23176,N23177,N23178,
N23179,N23180,N23181,N23182,N23183,N23184,N23185,N23186,N23187,N23188,
N23189,N23190,N23191,N23192,N23193,N23194,N23195,N23196,N23197,N23198,
N23199,N23200,N23201,N23202,N23203,N23204,N23205,N23206,N23207,N23208,
N23209,N23210,N23211,N23212,N23213,N23214,N23215,N23216,N23217,N23218,
N23219,N23220,N23221,N23222,N23223,N23224,N23225,N23226,N23227,N23228,
N23229,N23230,N23231,N23232,N23233,N23234,N23235,N23236,N23237,N23238,
N23239,N23240,N23241,N23242,N23243,N23244,N23245,N23246,N23247,N23248,
N23249,N23250,N23251,N23252,N23253,N23254,N23255,N23256,N23257,N23258,
N23259,N23260,N23261,N23262,N23263,N23264,N23265,N23266,N23267,N23268,
N23269,N23270,N23271,N23272,N23273,N23274,N23275,N23276,N23277,N23278,
N23279,N23280,N23281,N23282,N23283,N23284,N23285,N23286,N23287,N23288,
N23289,N23290,N23291,N23292,N23293,N23294,N23295,N23296,N23297,N23298,
N23299,N23300,N23301,N23302,N23303,N23304,N23305,N23306,N23307,N23308,
N23309,N23310,N23311,N23312,N23313,N23314,N23315,N23316,N23317,N23318,
N23319,N23320,N23321,N23322,N23323,N23324,N23325,N23326,N23327,N23328,
N23329,N23330,N23331,N23332,N23333,N23334,N23335,N23336,N23337,N23338,
N23339,N23340,N23341,N23342,N23343,N23344,N23345,N23346,N23347,N23348,
N23349,N23350,N23351,N23352,N23353,N23354,N23355,N23356,N23357,N23358,
N23359,N23360,N23361,N23362,N23363,N23364,N23365,N23366,N23367,N23368,
N23369,N23370,N23371,N23372,N23373,N23374,N23375,N23376,N23377,N23378,
N23379,N23380,N23381,N23382,N23383,N23384,N23385,N23386,N23387,N23388,
N23389,N23390,N23391,N23392,N23393,N23394,N23395,N23396,N23397,N23398,
N23399,N23400,N23401,N23402,N23403,N23404,N23405,N23406,N23407,N23408,
N23409,N23410,N23411,N23412,N23413,N23414,N23415,N23416,N23417,N23418,
N23419,N23420,N23421,N23422,N23423,N23424,N23425,N23426,N23427,N23428,
N23429,N23430,N23431,N23432,N23433,N23434,N23435,N23436,N23437,N23438,
N23439,N23440,N23441,N23442,N23443,N23444,N23445,N23446,N23447,N23448,
N23449,N23450,N23451,N23452,N23453,N23454,N23455,N23456,N23457,N23458,
N23459,N23460,N23461,N23462,N23463,N23464,N23465,N23466,N23467,N23468,
N23469,N23470,N23471,N23472,N23473,N23474,N23475,N23476,N23477,N23478,
N23479,N23480,N23481,N23482,N23483,N23484,N23485,N23486,N23487,N23488,
N23489,N23490,N23491,N23492,N23493,N23494,N23495,N23496,N23497,N23498,
N23499,N23500,N23501,N23502,N23503,N23504,N23505,N23506,N23507,N23508,
N23509,N23510,N23511,N23512,N23513,N23514,N23515,N23516,N23517,N23518,
N23519,N23520,N23521,N23522,N23523,N23524,N23525,N23526,N23527,N23528,
N23529,N23530,N23531,N23532,N23533,N23534,N23535,N23536,N23537,N23538,
N23539,N23540,N23541,N23542,N23543,N23544,N23545,N23546,N23547,N23548,
N23549,N23550,N23551,N23552,N23553,N23554,N23555,N23556,N23557,N23558,
N23559,N23560,N23561,N23562,N23563,N23564,N23565,N23566,N23567,N23568,
N23569,N23570,N23571,N23572,N23573,N23574,N23575,N23576,N23577,N23578,
N23579,N23580,N23581,N23582,N23583,N23584,N23585,N23586,N23587,N23588,
N23589,N23590,N23591,N23592,N23593,N23594,N23595,N23596,N23597,N23598,
N23599,N23600,N23601,N23602,N23603,N23604,N23605,N23606,N23607,N23608,
N23609,N23610,N23611,N23612,N23613,N23614,N23615,N23616,N23617,N23618,
N23619,N23620,N23621,N23622,N23623,N23624,N23625,N23626,N23627,N23628,
N23629,N23630,N23631,N23632,N23633,N23634,N23635,N23636,N23637,N23638,
N23639,N23640,N23641,N23642,N23643,N23644,N23645,N23646,N23647,N23648,
N23649,N23650,N23651,N23652,N23653,N23654,N23655,N23656,N23657,N23658,
N23659,N23660,N23661,N23662,N23663,N23664,N23665,N23666,N23667,N23668,
N23669,N23670,N23671,N23672,N23673,N23674,N23675,N23676,N23677,N23678,
N23679,N23680,N23681,N23682,N23683,N23684,N23685,N23686,N23687,N23688,
N23689,N23690,N23691,N23692,N23693,N23694,N23695,N23696,N23697,N23698,
N23699,N23700,N23701,N23702,N23703,N23704,N23705,N23706,N23707,N23708,
N23709,N23710,N23711,N23712,N23713,N23714,N23715,N23716,N23717,N23718,
N23719,N23720,N23721,N23722,N23723,N23724,N23725,N23726,N23727,N23728,
N23729,N23730,N23731,N23732,N23733,N23734,N23735,N23736,N23737,N23738,
N23739,N23740,N23741,N23742,N23743,N23744,N23745,N23746,N23747,N23748,
N23749,N23750,N23751,N23752,N23753,N23754,N23755,N23756,N23757,N23758,
N23759,N23760,N23761,N23762,N23763,N23764,N23765,N23766,N23767,N23768,
N23769,N23770,N23771,N23772,N23773,N23774,N23775,N23776,N23777,N23778,
N23779,N23780,N23781,N23782,N23783,N23784,N23785,N23786,N23787,N23788,
N23789,N23790,N23791,N23792,N23793,N23794,N23795,N23796,N23797,N23798,
N23799,N23800,N23801,N23802,N23803,N23804,N23805,N23806,N23807,N23808,
N23809,N23810,N23811,N23812,N23813,N23814,N23815,N23816,N23817,N23818,
N23819,N23820,N23821,N23822,N23823,N23824,N23825,N23826,N23827,N23828,
N23829,N23830,N23831,N23832,N23833,N23834,N23835,N23836,N23837,N23838,
N23839,N23840,N23841,N23842,N23843,N23844,N23845,N23846,N23847,N23848,
N23849,N23850,N23851,N23852,N23853,N23854,N23855,N23856,N23857,N23858,
N23859,N23860,N23861,N23862,N23863,N23864,N23865,N23866,N23867,N23868,
N23869,N23870,N23871,N23872,N23873,N23874,N23875,N23876,N23877,N23878,
N23879,N23880,N23881,N23882,N23883,N23884,N23885,N23886,N23887,N23888,
N23889,N23890,N23891,N23892,N23893,N23894,N23895,N23896,N23897,N23898,
N23899,N23900,N23901,N23902,N23903,N23904,N23905,N23906,N23907,N23908,
N23909,N23910,N23911,N23912,N23913,N23914,N23915,N23916,N23917,N23918,
N23919,N23920,N23921,N23922,N23923,N23924,N23925,N23926,N23927,N23928,
N23929,N23930,N23931,N23932,N23933,N23934,N23935,N23936,N23937,N23938,
N23939,N23940,N23941,N23942,N23943,N23944,N23945,N23946,N23947,N23948,
N23949,N23950,N23951,N23952,N23953,N23954,N23955,N23956,N23957,N23958,
N23959,N23960,N23961,N23962,N23963,N23964,N23965,N23966,N23967,N23968,
N23969,N23970,N23971,N23972,N23973,N23974,N23975,N23976,N23977,N23978,
N23979,N23980,N23981,N23982,N23983,N23984,N23985,N23986,N23987,N23988,
N23989,N23990,N23991,N23992,N23993,N23994,N23995,N23996,N23997,N23998,
N23999,N24000,N24001,N24002,N24003,N24004,N24005,N24006,N24007,N24008,
N24009,N24010,N24011,N24012,N24013,N24014,N24015,N24016,N24017,N24018,
N24019,N24020,N24021,N24022,N24023,N24024,N24025,N24026,N24027,N24028,
N24029,N24030,N24031,N24032,N24033,N24034,N24035,N24036,N24037,N24038,
N24039,N24040,N24041,N24042,N24043,N24044,N24045,N24046,N24047,N24048,
N24049,N24050,N24051,N24052,N24053,N24054,N24055,N24056,N24057,N24058,
N24059,N24060,N24061,N24062,N24063,N24064,N24065,N24066,N24067,N24068,
N24069,N24070,N24071,N24072,N24073,N24074,N24075,N24076,N24077,N24078,
N24079,N24080,N24081,N24082,N24083,N24084,N24085,N24086,N24087,N24088,
N24089,N24090,N24091,N24092,N24093,N24094,N24095,N24096,N24097,N24098,
N24099,N24100,N24101,N24102,N24103,N24104,N24105,N24106,N24107,N24108,
N24109,N24110,N24111,N24112,N24113,N24114,N24115,N24116,N24117,N24118,
N24119,N24120,N24121,N24122,N24123,N24124,N24125,N24126,N24127,N24128,
N24129,N24130,N24131,N24132,N24133,N24134,N24135,N24136,N24137,N24138,
N24139,N24140,N24141,N24142,N24143,N24144,N24145,N24146,N24147,N24148,
N24149,N24150,N24151,N24152,N24153,N24154,N24155,N24156,N24157,N24158,
N24159,N24160,N24161,N24162,N24163,N24164,N24165,N24166,N24167,N24168,
N24169,N24170,N24171,N24172,N24173,N24174,N24175,N24176,N24177,N24178,
N24179,N24180,N24181,N24182,N24183,N24184,N24185,N24186,N24187,N24188,
N24189,N24190,N24191,N24192,N24193,N24194,N24195,N24196,N24197,N24198,
N24199,N24200,N24201,N24202,N24203,N24204,N24205,N24206,N24207,N24208,
N24209,N24210,N24211,N24212,N24213,N24214,N24215,N24216,N24217,N24218,
N24219,N24220,N24221,N24222,N24223,N24224,N24225,N24226,N24227,N24228,
N24229,N24230,N24231,N24232,N24233,N24234,N24235,N24236,N24237,N24238,
N24239,N24240,N24241,N24242,N24243,N24244,N24245,N24246,N24247,N24248,
N24249,N24250,N24251,N24252,N24253,N24254,N24255,N24256,N24257,N24258,
N24259,N24260,N24261,N24262,N24263,N24264,N24265,N24266,N24267,N24268,
N24269,N24270,N24271,N24272,N24273,N24274,N24275,N24276,N24277,N24278,
N24279,N24280,N24281,N24282,N24283,N24284,N24285,N24286,N24287,N24288,
N24289,N24290,N24291,N24292,N24293,N24294,N24295,N24296,N24297,N24298,
N24299,N24300,N24301,N24302,N24303,N24304,N24305,N24306,N24307,N24308,
N24309,N24310,N24311,N24312,N24313,N24314,N24315,N24316,N24317,N24318,
N24319,N24320,N24321,N24322,N24323,N24324,N24325,N24326,N24327,N24328,
N24329,N24330,N24331,N24332,N24333,N24334,N24335,N24336,N24337,N24338,
N24339,N24340,N24341,N24342,N24343,N24344,N24345,N24346,N24347,N24348,
N24349,N24350,N24351,N24352,N24353,N24354,N24355,N24356,N24357,N24358,
N24359,N24360,N24361,N24362,N24363,N24364,N24365,N24366,N24367,N24368,
N24369,N24370,N24371,N24372,N24373,N24374,N24375,N24376,N24377,N24378,
N24379,N24380,N24381,N24382,N24383,N24384,N24385,N24386,N24387,N24388,
N24389,N24390,N24391,N24392,N24393,N24394,N24395,N24396,N24397,N24398,
N24399,N24400,N24401,N24402,N24403,N24404,N24405,N24406,N24407,N24408,
N24409,N24410,N24411,N24412,N24413,N24414,N24415,N24416,N24417,N24418,
N24419,N24420,N24421,N24422,N24423,N24424,N24425,N24426,N24427,N24428,
N24429,N24430,N24431,N24432,N24433,N24434,N24435,N24436,N24437,N24438,
N24439,N24440,N24441,N24442,N24443,N24444,N24445,N24446,N24447,N24448,
N24449,N24450,N24451,N24452,N24453,N24454,N24455,N24456,N24457,N24458,
N24459,N24460,N24461,N24462,N24463,N24464,N24465,N24466,N24467,N24468,
N24469,N24470,N24471,N24472,N24473,N24474,N24475,N24476,N24477,N24478,
N24479,N24480,N24481,N24482,N24483,N24484,N24485,N24486,N24487,N24488,
N24489,N24490,N24491,N24492,N24493,N24494,N24495,N24496,N24497,N24498,
N24499,N24500,N24501,N24502,N24503,N24504,N24505,N24506,N24507,N24508,
N24509,N24510,N24511,N24512,N24513,N24514,N24515,N24516,N24517,N24518,
N24519,N24520,N24521,N24522,N24523,N24524,N24525,N24526,N24527,N24528,
N24529,N24530,N24531,N24532,N24533,N24534,N24535,N24536,N24537,N24538,
N24539,N24540,N24541,N24542,N24543,N24544,N24545,N24546,N24547,N24548,
N24549,N24550,N24551,N24552,N24553,N24554,N24555,N24556,N24557,N24558,
N24559,N24560,N24561,N24562,N24563,N24564,N24565,N24566,N24567,N24568,
N24569,N24570,N24571,N24572,N24573,N24574,N24575,N24576,N24577,N24578,
N24579,N24580,N24581,N24582,N24583,N24584,N24585,N24586,N24587,N24588,
N24589,N24590,N24591,N24592,N24593,N24594,N24595,N24596,N24597,N24598,
N24599,N24600,N24601,N24602,N24603,N24604,N24605,N24606,N24607,N24608,
N24609,N24610,N24611,N24612,N24613,N24614,N24615,N24616,N24617,N24618,
N24619,N24620,N24621,N24622,N24623,N24624,N24625,N24626,N24627,N24628,
N24629,N24630,N24631,N24632,N24633,N24634,N24635,N24636,N24637,N24638,
N24639,N24640,N24641,N24642,N24643,N24644,N24645,N24646,N24647,N24648,
N24649,N24650,N24651,N24652,N24653,N24654,N24655,N24656,N24657,N24658,
N24659,N24660,N24661,N24662,N24663,N24664,N24665,N24666,N24667,N24668,
N24669,N24670,N24671,N24672,N24673,N24674,N24675,N24676,N24677,N24678,
N24679,N24680,N24681,N24682,N24683,N24684,N24685,N24686,N24687,N24688,
N24689,N24690,N24691,N24692,N24693,N24694,N24695,N24696,N24697,N24698,
N24699,N24700,N24701,N24702,N24703,N24704,N24705,N24706,N24707,N24708,
N24709,N24710,N24711,N24712,N24713,N24714,N24715,N24716,N24717,N24718,
N24719,N24720,N24721,N24722,N24723,N24724,N24725,N24726,N24727,N24728,
N24729,N24730,N24731,N24732,N24733,N24734,N24735,N24736,N24737,N24738,
N24739,N24740,N24741,N24742,N24743,N24744,N24745,N24746,N24747,N24748,
N24749,N24750,N24751,N24752,N24753,N24754,N24755,N24756,N24757,N24758,
N24759,N24760,N24761,N24762,N24763,N24764,N24765,N24766,N24767,N24768,
N24769,N24770,N24771,N24772,N24773,N24774,N24775,N24776,N24777,N24778,
N24779,N24780,N24781,N24782,N24783,N24784,N24785,N24786,N24787,N24788,
N24789,N24790,N24791,N24792,N24793,N24794,N24795,N24796,N24797,N24798,
N24799,N24800,N24801,N24802,N24803,N24804,N24805,N24806,N24807,N24808,
N24809,N24810,N24811,N24812,N24813,N24814,N24815,N24816,N24817,N24818,
N24819,N24820,N24821,N24822,N24823,N24824,N24825,N24826,N24827,N24828,
N24829,N24830,N24831,N24832,N24833,N24834,N24835,N24836,N24837,N24838,
N24839,N24840,N24841,N24842,N24843,N24844,N24845,N24846,N24847,N24848,
N24849,N24850,N24851,N24852,N24853,N24854,N24855,N24856,N24857,N24858,
N24859,N24860,N24861,N24862,N24863,N24864,N24865,N24866,N24867,N24868,
N24869,N24870,N24871,N24872,N24873,N24874,N24875,N24876,N24877,N24878,
N24879,N24880,N24881,N24882,N24883,N24884,N24885,N24886,N24887,N24888,
N24889,N24890,N24891,N24892,N24893,N24894,N24895,N24896,N24897,N24898,
N24899,N24900,N24901,N24902,N24903,N24904,N24905,N24906,N24907,N24908,
N24909,N24910,N24911,N24912,N24913,N24914,N24915,N24916,N24917,N24918,
N24919,N24920,N24921,N24922,N24923,N24924,N24925,N24926,N24927,N24928,
N24929,N24930,N24931,N24932,N24933,N24934,N24935,N24936,N24937,N24938,
N24939,N24940,N24941,N24942,N24943,N24944,N24945,N24946,N24947,N24948,
N24949,N24950,N24951,N24952,N24953,N24954,N24955,N24956,N24957,N24958,
N24959,N24960,N24961,N24962,N24963,N24964,N24965,N24966,N24967,N24968,
N24969,N24970,N24971,N24972,N24973,N24974,N24975,N24976,N24977,N24978,
N24979,N24980,N24981,N24982,N24983,N24984,N24985,N24986,N24987,N24988,
N24989,N24990,N24991,N24992,N24993,N24994,N24995,N24996,N24997,N24998,
N24999,N25000,N25001,N25002,N25003,N25004,N25005,N25006,N25007,N25008,
N25009,N25010,N25011,N25012,N25013,N25014,N25015,N25016,N25017,N25018,
N25019,N25020,N25021,N25022,N25023,N25024,N25025,N25026,N25027,N25028,
N25029,N25030,N25031,N25032,N25033,N25034,N25035,N25036,N25037,N25038,
N25039,N25040,N25041,N25042,N25043,N25044,N25045,N25046,N25047,N25048,
N25049,N25050,N25051,N25052,N25053,N25054,N25055,N25056,N25057,N25058,
N25059,N25060,N25061,N25062,N25063,N25064,N25065,N25066,N25067,N25068,
N25069,N25070,N25071,N25072,N25073,N25074,N25075,N25076,N25077,N25078,
N25079,N25080,N25081,N25082,N25083,N25084,N25085,N25086,N25087,N25088,
N25089,N25090,N25091,N25092,N25093,N25094,N25095,N25096,N25097,N25098,
N25099,N25100,N25101,N25102,N25103,N25104,N25105,N25106,N25107,N25108,
N25109,N25110,N25111,N25112,N25113,N25114,N25115,N25116,N25117,N25118,
N25119,N25120,N25121,N25122,N25123,N25124,N25125,N25126,N25127,N25128,
N25129,N25130,N25131,N25132,N25133,N25134,N25135,N25136,N25137,N25138,
N25139,N25140,N25141,N25142,N25143,N25144,N25145,N25146,N25147,N25148,
N25149,N25150,N25151,N25152,N25153,N25154,N25155,N25156,N25157,N25158,
N25159,N25160,N25161,N25162,N25163,N25164,N25165,N25166,N25167,N25168,
N25169,N25170,N25171,N25172,N25173,N25174,N25175,N25176,N25177,N25178,
N25179,N25180,N25181,N25182,N25183,N25184,N25185,N25186,N25187,N25188,
N25189,N25190,N25191,N25192,N25193,N25194,N25195,N25196,N25197,N25198,
N25199,N25200,N25201,N25202,N25203,N25204,N25205,N25206,N25207,N25208,
N25209,N25210,N25211,N25212,N25213,N25214,N25215,N25216,N25217,N25218,
N25219,N25220,N25221,N25222,N25223,N25224,N25225,N25226,N25227,N25228,
N25229,N25230,N25231,N25232,N25233,N25234,N25235,N25236,N25237,N25238,
N25239,N25240,N25241,N25242,N25243,N25244,N25245,N25246,N25247,N25248,
N25249,N25250,N25251,N25252,N25253,N25254,N25255,N25256,N25257,N25258,
N25259,N25260,N25261,N25262,N25263,N25264,N25265,N25266,N25267,N25268,
N25269,N25270,N25271,N25272,N25273,N25274,N25275,N25276,N25277,N25278,
N25279,N25280,N25281,N25282,N25283,N25284,N25285,N25286,N25287,N25288,
N25289,N25290,N25291,N25292,N25293,N25294,N25295,N25296,N25297,N25298,
N25299,N25300,N25301,N25302,N25303,N25304,N25305,N25306,N25307,N25308,
N25309,N25310,N25311,N25312,N25313,N25314,N25315,N25316,N25317,N25318,
N25319,N25320,N25321,N25322,N25323,N25324,N25325,N25326,N25327,N25328,
N25329,N25330,N25331,N25332,N25333,N25334,N25335,N25336,N25337,N25338,
N25339,N25340,N25341,N25342,N25343,N25344,N25345,N25346,N25347,N25348,
N25349,N25350,N25351,N25352,N25353,N25354,N25355,N25356,N25357,N25358,
N25359,N25360,N25361,N25362,N25363,N25364,N25365,N25366,N25367,N25368,
N25369,N25370,N25371,N25372,N25373,N25374,N25375,N25376,N25377,N25378,
N25379,N25380,N25381,N25382,N25383,N25384,N25385,N25386,N25387,N25388,
N25389,N25390,N25391,N25392,N25393,N25394,N25395,N25396,N25397,N25398,
N25399,N25400,N25401,N25402,N25403,N25404,N25405,N25406,N25407,N25408,
N25409,N25410,N25411,N25412,N25413,N25414,N25415,N25416,N25417,N25418,
N25419,N25420,N25421,N25422,N25423,N25424,N25425,N25426,N25427,N25428,
N25429,N25430,N25431,N25432,N25433,N25434,N25435,N25436,N25437,N25438,
N25439,N25440,N25441,N25442,N25443,N25444,N25445,N25446,N25447,N25448,
N25449,N25450,N25451,N25452,N25453,N25454,N25455,N25456,N25457,N25458,
N25459,N25460,N25461,N25462,N25463,N25464,N25465,N25466,N25467,N25468,
N25469,N25470,N25471,N25472,N25473,N25474,N25475,N25476,N25477,N25478,
N25479,N25480,N25481,N25482,N25483,N25484,N25485,N25486,N25487,N25488,
N25489,N25490,N25491,N25492,N25493,N25494,N25495,N25496,N25497,N25498,
N25499,N25500,N25501,N25502,N25503,N25504,N25505,N25506,N25507,N25508,
N25509,N25510,N25511,N25512,N25513,N25514,N25515,N25516,N25517,N25518,
N25519,N25520,N25521,N25522,N25523,N25524,N25525,N25526,N25527,N25528,
N25529,N25530,N25531,N25532,N25533,N25534,N25535,N25536,N25537,N25538,
N25539,N25540,N25541,N25542,N25543,N25544,N25545,N25546,N25547,N25548,
N25549,N25550,N25551,N25552,N25553,N25554,N25555,N25556,N25557,N25558,
N25559,N25560,N25561,N25562,N25563,N25564,N25565,N25566,N25567,N25568,
N25569,N25570,N25571,N25572,N25573,N25574,N25575,N25576,N25577,N25578,
N25579,N25580,N25581,N25582,N25583,N25584,N25585,N25586,N25587,N25588,
N25589,N25590,N25591,N25592,N25593,N25594,N25595,N25596,N25597,N25598,
N25599,N25600,N25601,N25602,N25603,N25604,N25605,N25606,N25607,N25608,
N25609,N25610,N25611,N25612,N25613,N25614,N25615,N25616,N25617,N25618,
N25619,N25620,N25621,N25622,N25623,N25624,N25625,N25626,N25627,N25628,
N25629,N25630,N25631,N25632,N25633,N25634,N25635,N25636,N25637,N25638,
N25639,N25640,N25641,N25642,N25643,N25644,N25645,N25646,N25647,N25648,
N25649,N25650,N25651,N25652,N25653,N25654,N25655,N25656,N25657,N25658,
N25659,N25660,N25661,N25662,N25663,N25664,N25665,N25666,N25667,N25668,
N25669,N25670,N25671,N25672,N25673,N25674,N25675,N25676,N25677,N25678,
N25679,N25680,N25681,N25682,N25683,N25684,N25685,N25686,N25687,N25688,
N25689,N25690,N25691,N25692,N25693,N25694,N25695,N25696,N25697,N25698,
N25699,N25700,N25701,N25702,N25703,N25704,N25705,N25706,N25707,N25708,
N25709,N25710,N25711,N25712,N25713,N25714,N25715,N25716,N25717,N25718,
N25719,N25720,N25721,N25722,N25723,N25724,N25725,N25726,N25727,N25728,
N25729,N25730,N25731,N25732,N25733,N25734,N25735,N25736,N25737,N25738,
N25739,N25740,N25741,N25742,N25743,N25744,N25745,N25746,N25747,N25748,
N25749,N25750,N25751,N25752,N25753,N25754,N25755,N25756,N25757,N25758,
N25759,N25760,N25761,N25762,N25763,N25764,N25765,N25766,N25767,N25768,
N25769,N25770,N25771,N25772,N25773,N25774,N25775,N25776,N25777,N25778,
N25779,N25780,N25781,N25782,N25783,N25784,N25785,N25786,N25787,N25788,
N25789,N25790,N25791,N25792,N25793,N25794,N25795,N25796,N25797,N25798,
N25799,N25800,N25801,N25802,N25803,N25804,N25805,N25806,N25807,N25808,
N25809,N25810,N25811,N25812,N25813,N25814,N25815,N25816,N25817,N25818,
N25819,N25820,N25821,N25822,N25823,N25824,N25825,N25826,N25827,N25828,
N25829,N25830,N25831,N25832,N25833,N25834,N25835,N25836,N25837,N25838,
N25839,N25840,N25841,N25842,N25843,N25844,N25845,N25846,N25847,N25848,
N25849,N25850,N25851,N25852,N25853,N25854,N25855,N25856,N25857,N25858,
N25859,N25860,N25861,N25862,N25863,N25864,N25865,N25866,N25867,N25868,
N25869,N25870,N25871,N25872,N25873,N25874,N25875,N25876,N25877,N25878,
N25879,N25880,N25881,N25882,N25883,N25884,N25885,N25886,N25887,N25888,
N25889,N25890,N25891,N25892,N25893,N25894,N25895,N25896,N25897,N25898,
N25899,N25900,N25901,N25902,N25903,N25904,N25905,N25906,N25907,N25908,
N25909,N25910,N25911,N25912,N25913,N25914,N25915,N25916,N25917,N25918,
N25919,N25920,N25921,N25922,N25923,N25924,N25925,N25926,N25927,N25928,
N25929,N25930,N25931,N25932,N25933,N25934,N25935,N25936,N25937,N25938,
N25939,N25940,N25941,N25942,N25943,N25944,N25945,N25946,N25947,N25948,
N25949,N25950,N25951,N25952,N25953,N25954,N25955,N25956,N25957,N25958,
N25959,N25960,N25961,N25962,N25963,N25964,N25965,N25966,N25967,N25968,
N25969,N25970,N25971,N25972,N25973,N25974,N25975,N25976,N25977,N25978,
N25979,N25980,N25981,N25982,N25983,N25984,N25985,N25986,N25987,N25988,
N25989,N25990,N25991,N25992,N25993,N25994,N25995,N25996,N25997,N25998,
N25999,N26000,N26001,N26002,N26003,N26004,N26005,N26006,N26007,N26008,
N26009,N26010,N26011,N26012,N26013,N26014,N26015,N26016,N26017,N26018,
N26019,N26020,N26021,N26022,N26023,N26024,N26025,N26026,N26027,N26028,
N26029,N26030,N26031,N26032,N26033,N26034,N26035,N26036,N26037,N26038,
N26039,N26040,N26041,N26042,N26043,N26044,N26045,N26046,N26047,N26048,
N26049,N26050,N26051,N26052,N26053,N26054,N26055,N26056,N26057,N26058,
N26059,N26060,N26061,N26062,N26063,N26064,N26065,N26066,N26067,N26068,
N26069,N26070,N26071,N26072,N26073,N26074,N26075,N26076,N26077,N26078,
N26079,N26080,N26081,N26082,N26083,N26084,N26085,N26086,N26087,N26088,
N26089,N26090,N26091,N26092,N26093,N26094,N26095,N26096,N26097,N26098,
N26099,N26100,N26101,N26102,N26103,N26104,N26105,N26106,N26107,N26108,
N26109,N26110,N26111,N26112,N26113,N26114,N26115,N26116,N26117,N26118,
N26119,N26120,N26121,N26122,N26123,N26124,N26125,N26126,N26127,N26128,
N26129,N26130,N26131,N26132,N26133,N26134,N26135,N26136,N26137,N26138,
N26139,N26140,N26141,N26142,N26143,N26144,N26145,N26146,N26147,N26148,
N26149,N26150,N26151,N26152,N26153,N26154,N26155,N26156,N26157,N26158,
N26159,N26160,N26161,N26162,N26163,N26164,N26165,N26166,N26167,N26168,
N26169,N26170,N26171,N26172,N26173,N26174,N26175,N26176,N26177,N26178,
N26179,N26180,N26181,N26182,N26183,N26184,N26185,N26186,N26187,N26188,
N26189,N26190,N26191,N26192,N26193,N26194,N26195,N26196,N26197,N26198,
N26199,N26200,N26201,N26202,N26203,N26204,N26205,N26206,N26207,N26208,
N26209,N26210,N26211,N26212,N26213,N26214,N26215,N26216,N26217,N26218,
N26219,N26220,N26221,N26222,N26223,N26224,N26225,N26226,N26227,N26228,
N26229,N26230,N26231,N26232,N26233,N26234,N26235,N26236,N26237,N26238,
N26239,N26240,N26241,N26242,N26243,N26244,N26245,N26246,N26247,N26248,
N26249,N26250,N26251,N26252,N26253,N26254,N26255,N26256,N26257,N26258,
N26259,N26260,N26261,N26262,N26263,N26264,N26265,N26266,N26267,N26268,
N26269,N26270,N26271,N26272,N26273,N26274,N26275,N26276,N26277,N26278,
N26279,N26280,N26281,N26282,N26283,N26284,N26285,N26286,N26287,N26288,
N26289,N26290,N26291,N26292,N26293,N26294,N26295,N26296,N26297,N26298,
N26299,N26300,N26301,N26302,N26303,N26304,N26305,N26306,N26307,N26308,
N26309,N26310,N26311,N26312,N26313,N26314,N26315,N26316,N26317,N26318,
N26319,N26320,N26321,N26322,N26323,N26324,N26325,N26326,N26327,N26328,
N26329,N26330,N26331,N26332,N26333,N26334,N26335,N26336,N26337,N26338,
N26339,N26340,N26341,N26342,N26343,N26344,N26345,N26346,N26347,N26348,
N26349,N26350,N26351,N26352,N26353,N26354,N26355,N26356,N26357,N26358,
N26359,N26360,N26361,N26362,N26363,N26364,N26365,N26366,N26367,N26368,
N26369,N26370,N26371,N26372,N26373,N26374,N26375,N26376,N26377,N26378,
N26379,N26380,N26381,N26382,N26383,N26384,N26385,N26386,N26387,N26388,
N26389,N26390,N26391,N26392,N26393,N26394,N26395,N26396,N26397,N26398,
N26399,N26400,N26401,N26402,N26403,N26404,N26405,N26406,N26407,N26408,
N26409,N26410,N26411,N26412,N26413,N26414,N26415,N26416,N26417,N26418,
N26419,N26420,N26421,N26422,N26423,N26424,N26425,N26426,N26427,N26428,
N26429,N26430,N26431,N26432,N26433,N26434,N26435,N26436,N26437,N26438,
N26439,N26440,N26441,N26442,N26443,N26444,N26445,N26446,N26447,N26448,
N26449,N26450,N26451,N26452,N26453,N26454,N26455,N26456,N26457,N26458,
N26459,N26460,N26461,N26462,N26463,N26464,N26465,N26466,N26467,N26468,
N26469,N26470,N26471,N26472,N26473,N26474,N26475,N26476,N26477,N26478,
N26479,N26480,N26481,N26482,N26483,N26484,N26485,N26486,N26487,N26488,
N26489,N26490,N26491,N26492,N26493,N26494,N26495,N26496,N26497,N26498,
N26499,N26500,N26501,N26502,N26503,N26504,N26505,N26506,N26507,N26508,
N26509,N26510,N26511,N26512,N26513,N26514,N26515,N26516,N26517,N26518,
N26519,N26520,N26521,N26522,N26523,N26524,N26525,N26526,N26527,N26528,
N26529,N26530,N26531,N26532,N26533,N26534,N26535,N26536,N26537,N26538,
N26539,N26540,N26541,N26542,N26543,N26544,N26545,N26546,N26547,N26548,
N26549,N26550,N26551,N26552,N26553,N26554,N26555,N26556,N26557,N26558,
N26559,N26560,N26561,N26562,N26563,N26564,N26565,N26566,N26567,N26568,
N26569,N26570,N26571,N26572,N26573,N26574,N26575,N26576,N26577,N26578,
N26579,N26580,N26581,N26582,N26583,N26584,N26585,N26586,N26587,N26588,
N26589,N26590,N26591,N26592,N26593,N26594,N26595,N26596,N26597,N26598,
N26599,N26600,N26601,N26602,N26603,N26604,N26605,N26606,N26607,N26608,
N26609,N26610,N26611,N26612,N26613,N26614,N26615,N26616,N26617,N26618,
N26619,N26620,N26621,N26622,N26623,N26624,N26625,N26626,N26627,N26628,
N26629,N26630,N26631,N26632,N26633,N26634,N26635,N26636,N26637,N26638,
N26639,N26640,N26641,N26642,N26643,N26644,N26645,N26646,N26647,N26648,
N26649,N26650,N26651,N26652,N26653,N26654,N26655,N26656,N26657,N26658,
N26659,N26660,N26661,N26662,N26663,N26664,N26665,N26666,N26667,N26668,
N26669,N26670,N26671,N26672,N26673,N26674,N26675,N26676,N26677,N26678,
N26679,N26680,N26681,N26682,N26683,N26684,N26685,N26686,N26687,N26688,
N26689,N26690,N26691,N26692,N26693,N26694,N26695,N26696,N26697,N26698,
N26699,N26700,N26701,N26702,N26703,N26704,N26705,N26706,N26707,N26708,
N26709,N26710,N26711,N26712,N26713,N26714,N26715,N26716,N26717,N26718,
N26719,N26720,N26721,N26722,N26723,N26724,N26725,N26726,N26727,N26728,
N26729,N26730,N26731,N26732,N26733,N26734,N26735,N26736,N26737,N26738,
N26739,N26740,N26741,N26742,N26743,N26744,N26745,N26746,N26747,N26748,
N26749,N26750,N26751,N26752,N26753,N26754,N26755,N26756,N26757,N26758,
N26759,N26760,N26761,N26762,N26763,N26764,N26765,N26766,N26767,N26768,
N26769,N26770,N26771,N26772,N26773,N26774,N26775,N26776,N26777,N26778,
N26779,N26780,N26781,N26782,N26783,N26784,N26785,N26786,N26787,N26788,
N26789,N26790,N26791,N26792,N26793,N26794,N26795,N26796,N26797,N26798,
N26799,N26800,N26801,N26802,N26803,N26804,N26805,N26806,N26807,N26808,
N26809,N26810,N26811,N26812,N26813,N26814,N26815,N26816,N26817,N26818,
N26819,N26820,N26821,N26822,N26823,N26824,N26825,N26826,N26827,N26828,
N26829,N26830,N26831,N26832,N26833,N26834,N26835,N26836,N26837,N26838,
N26839,N26840,N26841,N26842,N26843,N26844,N26845,N26846,N26847,N26848,
N26849,N26850,N26851,N26852,N26853,N26854,N26855,N26856,N26857,N26858,
N26859,N26860,N26861,N26862,N26863,N26864,N26865,N26866,N26867,N26868,
N26869,N26870,N26871,N26872,N26873,N26874,N26875,N26876,N26877,N26878,
N26879,N26880,N26881,N26882,N26883,N26884,N26885,N26886,N26887,N26888,
N26889,N26890,N26891,N26892,N26893,N26894,N26895,N26896,N26897,N26898,
N26899,N26900,N26901,N26902,N26903,N26904,N26905,N26906,N26907,N26908,
N26909,N26910,N26911,N26912,N26913,N26914,N26915,N26916,N26917,N26918,
N26919,N26920,N26921,N26922,N26923,N26924,N26925,N26926,N26927,N26928,
N26929,N26930,N26931,N26932,N26933,N26934,N26935,N26936,N26937,N26938,
N26939,N26940,N26941,N26942,N26943,N26944,N26945,N26946,N26947,N26948,
N26949,N26950,N26951,N26952,N26953,N26954,N26955,N26956,N26957,N26958,
N26959,N26960,N26961,N26962,N26963,N26964,N26965,N26966,N26967,N26968,
N26969,N26970,N26971,N26972,N26973,N26974,N26975,N26976,N26977,N26978,
N26979,N26980,N26981,N26982,N26983,N26984,N26985,N26986,N26987,N26988,
N26989,N26990,N26991,N26992,N26993,N26994,N26995,N26996,N26997,N26998,
N26999,N27000,N27001,N27002,N27003,N27004,N27005,N27006,N27007,N27008,
N27009,N27010,N27011,N27012,N27013,N27014,N27015,N27016,N27017,N27018,
N27019,N27020,N27021,N27022,N27023,N27024,N27025,N27026,N27027,N27028,
N27029,N27030,N27031,N27032,N27033,N27034,N27035,N27036,N27037,N27038,
N27039,N27040,N27041,N27042,N27043,N27044,N27045,N27046,N27047,N27048,
N27049,N27050,N27051,N27052,N27053,N27054,N27055,N27056,N27057,N27058,
N27059,N27060,N27061,N27062,N27063,N27064,N27065,N27066,N27067,N27068,
N27069,N27070,N27071,N27072,N27073,N27074,N27075,N27076,N27077,N27078,
N27079,N27080,N27081,N27082,N27083,N27084,N27085,N27086,N27087,N27088,
N27089,N27090,N27091,N27092,N27093,N27094,N27095,N27096,N27097,N27098,
N27099,N27100,N27101,N27102,N27103,N27104,N27105,N27106,N27107,N27108,
N27109,N27110,N27111,N27112,N27113,N27114,N27115,N27116,N27117,N27118,
N27119,N27120,N27121,N27122,N27123,N27124,N27125,N27126,N27127,N27128,
N27129,N27130,N27131,N27132,N27133,N27134,N27135,N27136,N27137,N27138,
N27139,N27140,N27141,N27142,N27143,N27144,N27145,N27146,N27147,N27148,
N27149,N27150,N27151,N27152,N27153,N27154,N27155,N27156,N27157,N27158,
N27159,N27160,N27161,N27162,N27163,N27164,N27165,N27166,N27167,N27168,
N27169,N27170,N27171,N27172,N27173,N27174,N27175,N27176,N27177,N27178,
N27179,N27180,N27181,N27182,N27183,N27184,N27185,N27186,N27187,N27188,
N27189,N27190,N27191,N27192,N27193,N27194,N27195,N27196,N27197,N27198,
N27199,N27200,N27201,N27202,N27203,N27204,N27205,N27206,N27207,N27208,
N27209,N27210,N27211,N27212,N27213,N27214,N27215,N27216,N27217,N27218,
N27219,N27220,N27221,N27222,N27223,N27224,N27225,N27226,N27227,N27228,
N27229,N27230,N27231,N27232,N27233,N27234,N27235,N27236,N27237,N27238,
N27239,N27240,N27241,N27242,N27243,N27244,N27245,N27246,N27247,N27248,
N27249,N27250,N27251,N27252,N27253,N27254,N27255,N27256,N27257,N27258,
N27259,N27260,N27261,N27262,N27263,N27264,N27265,N27266,N27267,N27268,
N27269,N27270,N27271,N27272,N27273,N27274,N27275,N27276,N27277,N27278,
N27279,N27280,N27281,N27282,N27283,N27284,N27285,N27286,N27287,N27288,
N27289,N27290,N27291,N27292,N27293,N27294,N27295,N27296,N27297,N27298,
N27299,N27300,N27301,N27302,N27303,N27304,N27305,N27306,N27307,N27308,
N27309,N27310,N27311,N27312,N27313,N27314,N27315,N27316,N27317,N27318,
N27319,N27320,N27321,N27322,N27323,N27324,N27325,N27326,N27327,N27328,
N27329,N27330,N27331,N27332,N27333,N27334,N27335,N27336,N27337,N27338,
N27339,N27340,N27341,N27342,N27343,N27344,N27345,N27346,N27347,N27348,
N27349,N27350,N27351,N27352,N27353,N27354,N27355,N27356,N27357,N27358,
N27359,N27360,N27361,N27362,N27363,N27364,N27365,N27366,N27367,N27368,
N27369,N27370,N27371,N27372,N27373,N27374,N27375,N27376,N27377,N27378,
N27379,N27380,N27381,N27382,N27383,N27384,N27385,N27386,N27387,N27388,
N27389,N27390,N27391,N27392,N27393,N27394,N27395,N27396,N27397,N27398,
N27399,N27400,N27401,N27402,N27403,N27404,N27405,N27406,N27407,N27408,
N27409,N27410,N27411,N27412,N27413,N27414,N27415,N27416,N27417,N27418,
N27419,N27420,N27421,N27422,N27423,N27424,N27425,N27426,N27427,N27428,
N27429,N27430,N27431,N27432,N27433,N27434,N27435,N27436,N27437,N27438,
N27439,N27440,N27441,N27442,N27443,N27444,N27445,N27446,N27447,N27448,
N27449,N27450,N27451,N27452,N27453,N27454,N27455,N27456,N27457,N27458,
N27459,N27460,N27461,N27462,N27463,N27464,N27465,N27466,N27467,N27468,
N27469,N27470,N27471,N27472,N27473,N27474,N27475,N27476,N27477,N27478,
N27479,N27480,N27481,N27482,N27483,N27484,N27485,N27486,N27487,N27488,
N27489,N27490,N27491,N27492,N27493,N27494,N27495,N27496,N27497,N27498,
N27499,N27500,N27501,N27502,N27503,N27504,N27505,N27506,N27507,N27508,
N27509,N27510,N27511,N27512,N27513,N27514,N27515,N27516,N27517,N27518,
N27519,N27520,N27521,N27522,N27523,N27524,N27525,N27526,N27527,N27528,
N27529,N27530,N27531,N27532,N27533,N27534,N27535,N27536,N27537,N27538,
N27539,N27540,N27541,N27542,N27543,N27544,N27545,N27546,N27547,N27548,
N27549,N27550,N27551,N27552,N27553,N27554,N27555,N27556,N27557,N27558,
N27559,N27560,N27561,N27562,N27563,N27564,N27565,N27566,N27567,N27568,
N27569,N27570,N27571,N27572,N27573,N27574,N27575,N27576,N27577,N27578,
N27579,N27580,N27581,N27582,N27583,N27584,N27585,N27586,N27587,N27588,
N27589,N27590,N27591,N27592,N27593,N27594,N27595,N27596,N27597,N27598,
N27599,N27600,N27601,N27602,N27603,N27604,N27605,N27606,N27607,N27608,
N27609,N27610,N27611,N27612,N27613,N27614,N27615,N27616,N27617,N27618,
N27619,N27620,N27621,N27622,N27623,N27624,N27625,N27626,N27627,N27628,
N27629,N27630,N27631,N27632,N27633,N27634,N27635,N27636,N27637,N27638,
N27639,N27640,N27641,N27642,N27643,N27644,N27645,N27646,N27647,N27648,
N27649,N27650,N27651,N27652,N27653,N27654,N27655,N27656,N27657,N27658,
N27659,N27660,N27661,N27662,N27663,N27664,N27665,N27666,N27667,N27668,
N27669,N27670,N27671,N27672,N27673,N27674,N27675,N27676,N27677,N27678,
N27679,N27680,N27681,N27682,N27683,N27684,N27685,N27686,N27687,N27688,
N27689,N27690,N27691,N27692,N27693,N27694,N27695,N27696,N27697,N27698,
N27699,N27700,N27701,N27702,N27703,N27704,N27705,N27706,N27707,N27708,
N27709,N27710,N27711,N27712,N27713,N27714,N27715,N27716,N27717,N27718,
N27719,N27720,N27721,N27722,N27723,N27724,N27725,N27726,N27727,N27728,
N27729,N27730,N27731,N27732,N27733,N27734,N27735,N27736,N27737,N27738,
N27739,N27740,N27741,N27742,N27743,N27744,N27745,N27746,N27747,N27748,
N27749,N27750,N27751,N27752,N27753,N27754,N27755,N27756,N27757,N27758,
N27759,N27760,N27761,N27762,N27763,N27764,N27765,N27766,N27767,N27768,
N27769,N27770,N27771,N27772,N27773,N27774,N27775,N27776,N27777,N27778,
N27779,N27780,N27781,N27782,N27783,N27784,N27785,N27786,N27787,N27788,
N27789,N27790,N27791,N27792,N27793,N27794,N27795,N27796,N27797,N27798,
N27799,N27800,N27801,N27802,N27803,N27804,N27805,N27806,N27807,N27808,
N27809,N27810,N27811,N27812,N27813,N27814,N27815,N27816,N27817,N27818,
N27819,N27820,N27821,N27822,N27823,N27824,N27825,N27826,N27827,N27828,
N27829,N27830,N27831,N27832,N27833,N27834,N27835,N27836,N27837,N27838,
N27839,N27840,N27841,N27842,N27843,N27844,N27845,N27846,N27847,N27848,
N27849,N27850,N27851,N27852,N27853,N27854,N27855,N27856,N27857,N27858,
N27859,N27860,N27861,N27862,N27863,N27864,N27865,N27866,N27867,N27868,
N27869,N27870,N27871,N27872,N27873,N27874,N27875,N27876,N27877,N27878,
N27879,N27880,N27881,N27882,N27883,N27884,N27885,N27886,N27887,N27888,
N27889,N27890,N27891,N27892,N27893,N27894,N27895,N27896,N27897,N27898,
N27899,N27900,N27901,N27902,N27903,N27904,N27905,N27906,N27907,N27908,
N27909,N27910,N27911,N27912,N27913,N27914,N27915,N27916,N27917,N27918,
N27919,N27920,N27921,N27922,N27923,N27924,N27925,N27926,N27927,N27928,
N27929,N27930,N27931,N27932,N27933,N27934,N27935,N27936,N27937,N27938,
N27939,N27940,N27941,N27942,N27943,N27944,N27945,N27946,N27947,N27948,
N27949,N27950,N27951,N27952,N27953,N27954,N27955,N27956,N27957,N27958,
N27959,N27960,N27961,N27962,N27963,N27964,N27965,N27966,N27967,N27968,
N27969,N27970,N27971,N27972,N27973,N27974,N27975,N27976,N27977,N27978,
N27979,N27980,N27981,N27982,N27983,N27984,N27985,N27986,N27987,N27988,
N27989,N27990,N27991,N27992,N27993,N27994,N27995,N27996,N27997,N27998,
N27999,N28000,N28001,N28002,N28003,N28004,N28005,N28006,N28007,N28008,
N28009,N28010,N28011,N28012,N28013,N28014,N28015,N28016,N28017,N28018,
N28019,N28020,N28021,N28022,N28023,N28024,N28025,N28026,N28027,N28028,
N28029,N28030,N28031,N28032,N28033,N28034,N28035,N28036,N28037,N28038,
N28039,N28040,N28041,N28042,N28043,N28044,N28045,N28046,N28047,N28048,
N28049,N28050,N28051,N28052,N28053,N28054,N28055,N28056,N28057,N28058,
N28059,N28060,N28061,N28062,N28063,N28064,N28065,N28066,N28067,N28068,
N28069,N28070,N28071,N28072,N28073,N28074,N28075,N28076,N28077,N28078,
N28079,N28080,N28081,N28082,N28083,N28084,N28085,N28086,N28087,N28088,
N28089,N28090,N28091,N28092,N28093,N28094,N28095,N28096,N28097,N28098,
N28099,N28100,N28101,N28102,N28103,N28104,N28105,N28106,N28107,N28108,
N28109,N28110,N28111,N28112,N28113,N28114,N28115,N28116,N28117,N28118,
N28119,N28120,N28121,N28122,N28123,N28124,N28125,N28126,N28127,N28128,
N28129,N28130,N28131,N28132,N28133,N28134,N28135,N28136,N28137,N28138,
N28139,N28140,N28141,N28142,N28143,N28144,N28145,N28146,N28147,N28148,
N28149,N28150,N28151,N28152,N28153,N28154,N28155,N28156,N28157,N28158,
N28159,N28160,N28161,N28162,N28163,N28164,N28165,N28166,N28167,N28168,
N28169,N28170,N28171,N28172,N28173,N28174,N28175,N28176,N28177,N28178,
N28179,N28180,N28181,N28182,N28183,N28184,N28185,N28186,N28187,N28188,
N28189,N28190,N28191,N28192,N28193,N28194,N28195,N28196,N28197,N28198,
N28199,N28200,N28201,N28202,N28203,N28204,N28205,N28206,N28207,N28208,
N28209,N28210,N28211,N28212,N28213,N28214,N28215,N28216,N28217,N28218,
N28219,N28220,N28221,N28222,N28223,N28224,N28225,N28226,N28227,N28228,
N28229,N28230,N28231,N28232,N28233,N28234,N28235,N28236,N28237,N28238,
N28239,N28240,N28241,N28242,N28243,N28244,N28245,N28246,N28247,N28248,
N28249,N28250,N28251,N28252,N28253,N28254,N28255,N28256,N28257,N28258,
N28259,N28260,N28261,N28262,N28263,N28264,N28265,N28266,N28267,N28268,
N28269,N28270,N28271,N28272,N28273,N28274,N28275,N28276,N28277,N28278,
N28279,N28280,N28281,N28282,N28283,N28284,N28285,N28286,N28287,N28288,
N28289,N28290,N28291,N28292,N28293,N28294,N28295,N28296,N28297,N28298,
N28299,N28300,N28301,N28302,N28303,N28304,N28305,N28306,N28307,N28308,
N28309,N28310,N28311,N28312,N28313,N28314,N28315,N28316,N28317,N28318,
N28319,N28320,N28321,N28322,N28323,N28324,N28325,N28326,N28327,N28328,
N28329,N28330,N28331,N28332,N28333,N28334,N28335,N28336,N28337,N28338,
N28339,N28340,N28341,N28342,N28343,N28344,N28345,N28346,N28347,N28348,
N28349,N28350,N28351,N28352,N28353,N28354,N28355,N28356,N28357,N28358,
N28359,N28360,N28361,N28362,N28363,N28364,N28365,N28366,N28367,N28368,
N28369,N28370,N28371,N28372,N28373,N28374,N28375,N28376,N28377,N28378,
N28379,N28380,N28381,N28382,N28383,N28384,N28385,N28386,N28387,N28388,
N28389,N28390,N28391,N28392,N28393,N28394,N28395,N28396,N28397,N28398,
N28399,N28400,N28401,N28402,N28403,N28404,N28405,N28406,N28407,N28408,
N28409,N28410,N28411,N28412,N28413,N28414,N28415,N28416,N28417,N28418,
N28419,N28420,N28421,N28422,N28423,N28424,N28425,N28426,N28427,N28428,
N28429,N28430,N28431,N28432,N28433,N28434,N28435,N28436,N28437,N28438,
N28439,N28440,N28441,N28442,N28443,N28444,N28445,N28446,N28447,N28448,
N28449,N28450,N28451,N28452,N28453,N28454,N28455,N28456,N28457,N28458,
N28459,N28460,N28461,N28462,N28463,N28464,N28465,N28466,N28467,N28468,
N28469,N28470,N28471,N28472,N28473,N28474,N28475,N28476,N28477,N28478,
N28479,N28480,N28481,N28482,N28483,N28484,N28485,N28486,N28487,N28488,
N28489,N28490,N28491,N28492,N28493,N28494,N28495,N28496,N28497,N28498,
N28499,N28500,N28501,N28502,N28503,N28504,N28505,N28506,N28507,N28508,
N28509,N28510,N28511,N28512,N28513,N28514,N28515,N28516,N28517,N28518,
N28519,N28520,N28521,N28522,N28523,N28524,N28525,N28526,N28527,N28528,
N28529,N28530,N28531,N28532,N28533,N28534,N28535,N28536,N28537,N28538,
N28539,N28540,N28541,N28542,N28543,N28544,N28545,N28546,N28547,N28548,
N28549,N28550,N28551,N28552,N28553,N28554,N28555,N28556,N28557,N28558,
N28559,N28560,N28561,N28562,N28563,N28564,N28565,N28566,N28567,N28568,
N28569,N28570,N28571,N28572,N28573,N28574,N28575,N28576,N28577,N28578,
N28579,N28580,N28581,N28582,N28583,N28584,N28585,N28586,N28587,N28588,
N28589,N28590,N28591,N28592,N28593,N28594,N28595,N28596,N28597,N28598,
N28599,N28600,N28601,N28602,N28603,N28604,N28605,N28606,N28607,N28608,
N28609,N28610,N28611,N28612,N28613,N28614,N28615,N28616,N28617,N28618,
N28619,N28620,N28621,N28622,N28623,N28624,N28625,N28626,N28627,N28628,
N28629,N28630,N28631,N28632,N28633,N28634,N28635,N28636,N28637,N28638,
N28639,N28640,N28641,N28642,N28643,N28644,N28645,N28646,N28647,N28648,
N28649,N28650,N28651,N28652,N28653,N28654,N28655,N28656,N28657,N28658,
N28659,N28660,N28661,N28662,N28663,N28664,N28665,N28666,N28667,N28668,
N28669,N28670,N28671,N28672,N28673,N28674,N28675,N28676,N28677,N28678,
N28679,N28680,N28681,N28682,N28683,N28684,N28685,N28686,N28687,N28688,
N28689,N28690,N28691,N28692,N28693,N28694,N28695,N28696,N28697,N28698,
N28699,N28700,N28701,N28702,N28703,N28704,N28705,N28706,N28707,N28708,
N28709,N28710,N28711,N28712,N28713,N28714,N28715,N28716,N28717,N28718,
N28719,N28720,N28721,N28722,N28723,N28724,N28725,N28726,N28727,N28728,
N28729,N28730,N28731,N28732,N28733,N28734,N28735,N28736,N28737,N28738,
N28739,N28740,N28741,N28742,N28743,N28744,N28745,N28746,N28747,N28748,
N28749,N28750,N28751,N28752,N28753,N28754,N28755,N28756,N28757,N28758,
N28759,N28760,N28761,N28762,N28763,N28764,N28765,N28766,N28767,N28768,
N28769,N28770,N28771,N28772,N28773,N28774,N28775,N28776,N28777,N28778,
N28779,N28780,N28781,N28782,N28783,N28784,N28785,N28786,N28787,N28788,
N28789,N28790,N28791,N28792,N28793,N28794,N28795,N28796,N28797,N28798,
N28799,N28800,N28801,N28802,N28803,N28804,N28805,N28806,N28807,N28808,
N28809,N28810,N28811,N28812,N28813,N28814,N28815,N28816,N28817,N28818,
N28819,N28820,N28821,N28822,N28823,N28824,N28825,N28826,N28827,N28828,
N28829,N28830,N28831,N28832,N28833,N28834,N28835,N28836,N28837,N28838,
N28839,N28840,N28841,N28842,N28843,N28844,N28845,N28846,N28847,N28848,
N28849,N28850,N28851,N28852,N28853,N28854,N28855,N28856,N28857,N28858,
N28859,N28860,N28861,N28862,N28863,N28864,N28865,N28866,N28867,N28868,
N28869,N28870,N28871,N28872,N28873,N28874,N28875,N28876,N28877,N28878,
N28879,N28880,N28881,N28882,N28883,N28884,N28885,N28886,N28887,N28888,
N28889,N28890,N28891,N28892,N28893,N28894,N28895,N28896,N28897,N28898,
N28899,N28900,N28901,N28902,N28903,N28904,N28905,N28906,N28907,N28908,
N28909,N28910,N28911,N28912,N28913,N28914,N28915,N28916,N28917,N28918,
N28919,N28920,N28921,N28922,N28923,N28924,N28925,N28926,N28927,N28928,
N28929,N28930,N28931,N28932,N28933,N28934,N28935,N28936,N28937,N28938,
N28939,N28940,N28941,N28942,N28943,N28944,N28945,N28946,N28947,N28948,
N28949,N28950,N28951,N28952,N28953,N28954,N28955,N28956,N28957,N28958,
N28959,N28960,N28961,N28962,N28963,N28964,N28965,N28966,N28967,N28968,
N28969,N28970,N28971,N28972,N28973,N28974,N28975,N28976,N28977,N28978,
N28979,N28980,N28981,N28982,N28983,N28984,N28985,N28986,N28987,N28988,
N28989,N28990,N28991,N28992,N28993,N28994,N28995,N28996,N28997,N28998,
N28999,N29000,N29001,N29002,N29003,N29004,N29005,N29006,N29007,N29008,
N29009,N29010,N29011,N29012,N29013,N29014,N29015,N29016,N29017,N29018,
N29019,N29020,N29021,N29022,N29023,N29024,N29025,N29026,N29027,N29028,
N29029,N29030,N29031,N29032,N29033,N29034,N29035,N29036,N29037,N29038,
N29039,N29040,N29041,N29042,N29043,N29044,N29045,N29046,N29047,N29048,
N29049,N29050,N29051,N29052,N29053,N29054,N29055,N29056,N29057,N29058,
N29059,N29060,N29061,N29062,N29063,N29064,N29065,N29066,N29067,N29068,
N29069,N29070,N29071,N29072,N29073,N29074,N29075,N29076,N29077,N29078,
N29079,N29080,N29081,N29082,N29083,N29084,N29085,N29086,N29087,N29088,
N29089,N29090,N29091,N29092,N29093,N29094,N29095,N29096,N29097,N29098,
N29099,N29100,N29101,N29102,N29103,N29104,N29105,N29106,N29107,N29108,
N29109,N29110,N29111,N29112,N29113,N29114,N29115,N29116,N29117,N29118,
N29119,N29120,N29121,N29122,N29123,N29124,N29125,N29126,N29127,N29128,
N29129,N29130,N29131,N29132,N29133,N29134,N29135,N29136,N29137,N29138,
N29139,N29140,N29141,N29142,N29143,N29144,N29145,N29146,N29147,N29148,
N29149,N29150,N29151,N29152,N29153,N29154,N29155,N29156,N29157,N29158,
N29159,N29160,N29161,N29162,N29163,N29164,N29165,N29166,N29167,N29168,
N29169,N29170,N29171,N29172,N29173,N29174,N29175,N29176,N29177,N29178,
N29179,N29180,N29181,N29182,N29183,N29184,N29185,N29186,N29187,N29188,
N29189,N29190,N29191,N29192,N29193,N29194,N29195,N29196,N29197,N29198,
N29199,N29200,N29201,N29202,N29203,N29204,N29205,N29206,N29207,N29208,
N29209,N29210,N29211,N29212,N29213,N29214,N29215,N29216,N29217,N29218,
N29219,N29220,N29221,N29222,N29223,N29224,N29225,N29226,N29227,N29228,
N29229,N29230,N29231,N29232,N29233,N29234,N29235,N29236,N29237,N29238,
N29239,N29240,N29241,N29242,N29243,N29244,N29245,N29246,N29247,N29248,
N29249,N29250,N29251,N29252,N29253,N29254,N29255,N29256,N29257,N29258,
N29259,N29260,N29261,N29262,N29263,N29264,N29265,N29266,N29267,N29268,
N29269,N29270,N29271,N29272,N29273,N29274,N29275,N29276,N29277,N29278,
N29279,N29280,N29281,N29282,N29283,N29284,N29285,N29286,N29287,N29288,
N29289,N29290,N29291,N29292,N29293,N29294,N29295,N29296,N29297,N29298,
N29299,N29300,N29301,N29302,N29303,N29304,N29305,N29306,N29307,N29308,
N29309,N29310,N29311,N29312,N29313,N29314,N29315,N29316,N29317,N29318,
N29319,N29320,N29321,N29322,N29323,N29324,N29325,N29326,N29327,N29328,
N29329,N29330,N29331,N29332,N29333,N29334,N29335,N29336,N29337,N29338,
N29339,N29340,N29341,N29342,N29343,N29344,N29345,N29346,N29347,N29348,
N29349,N29350,N29351,N29352,N29353,N29354,N29355,N29356,N29357,N29358,
N29359,N29360,N29361,N29362,N29363,N29364,N29365,N29366,N29367,N29368,
N29369,N29370,N29371,N29372,N29373,N29374,N29375,N29376,N29377,N29378,
N29379,N29380,N29381,N29382,N29383,N29384,N29385,N29386,N29387,N29388,
N29389,N29390,N29391,N29392,N29393,N29394,N29395,N29396,N29397,N29398,
N29399,N29400,N29401,N29402,N29403,N29404,N29405,N29406,N29407,N29408,
N29409,N29410,N29411,N29412,N29413,N29414,N29415,N29416,N29417,N29418,
N29419,N29420,N29421,N29422,N29423,N29424,N29425,N29426,N29427,N29428,
N29429,N29430,N29431,N29432,N29433,N29434,N29435,N29436,N29437,N29438,
N29439,N29440,N29441,N29442,N29443,N29444,N29445,N29446,N29447,N29448,
N29449,N29450,N29451,N29452,N29453,N29454,N29455,N29456,N29457,N29458,
N29459,N29460,N29461,N29462,N29463,N29464,N29465,N29466,N29467,N29468,
N29469,N29470,N29471,N29472,N29473,N29474,N29475,N29476,N29477,N29478,
N29479,N29480,N29481,N29482,N29483,N29484,N29485,N29486,N29487,N29488,
N29489,N29490,N29491,N29492,N29493,N29494,N29495,N29496,N29497,N29498,
N29499,N29500,N29501,N29502,N29503,N29504,N29505,N29506,N29507,N29508,
N29509,N29510,N29511,N29512,N29513,N29514,N29515,N29516,N29517,N29518,
N29519,N29520,N29521,N29522,N29523,N29524,N29525,N29526,N29527,N29528,
N29529,N29530,N29531,N29532,N29533,N29534,N29535,N29536,N29537,N29538,
N29539,N29540,N29541,N29542,N29543,N29544,N29545,N29546,N29547,N29548,
N29549,N29550,N29551,N29552,N29553,N29554,N29555,N29556,N29557,N29558,
N29559,N29560,N29561,N29562,N29563,N29564,N29565,N29566,N29567,N29568,
N29569,N29570,N29571,N29572,N29573,N29574,N29575,N29576,N29577,N29578,
N29579,N29580,N29581,N29582,N29583,N29584,N29585,N29586,N29587,N29588,
N29589,N29590,N29591,N29592,N29593,N29594,N29595,N29596,N29597,N29598,
N29599,N29600,N29601,N29602,N29603,N29604,N29605,N29606,N29607,N29608,
N29609,N29610,N29611,N29612,N29613,N29614,N29615,N29616,N29617,N29618,
N29619,N29620,N29621,N29622,N29623,N29624,N29625,N29626,N29627,N29628,
N29629,N29630,N29631,N29632,N29633,N29634,N29635,N29636,N29637,N29638,
N29639,N29640,N29641,N29642,N29643,N29644,N29645,N29646,N29647,N29648,
N29649,N29650,N29651,N29652,N29653,N29654,N29655,N29656,N29657,N29658,
N29659,N29660,N29661,N29662,N29663,N29664,N29665,N29666,N29667,N29668,
N29669,N29670,N29671,N29672,N29673,N29674,N29675,N29676,N29677,N29678,
N29679,N29680,N29681,N29682,N29683,N29684,N29685,N29686,N29687,N29688,
N29689,N29690,N29691,N29692,N29693,N29694,N29695,N29696,N29697,N29698,
N29699,N29700,N29701,N29702,N29703,N29704,N29705,N29706,N29707,N29708,
N29709,N29710,N29711,N29712,N29713,N29714,N29715,N29716,N29717,N29718,
N29719,N29720,N29721,N29722,N29723,N29724,N29725,N29726,N29727,N29728,
N29729,N29730,N29731,N29732,N29733,N29734,N29735,N29736,N29737,N29738,
N29739,N29740,N29741,N29742,N29743,N29744,N29745,N29746,N29747,N29748,
N29749,N29750,N29751,N29752,N29753,N29754,N29755,N29756,N29757,N29758,
N29759,N29760,N29761,N29762,N29763,N29764,N29765,N29766,N29767,N29768,
N29769,N29770,N29771,N29772,N29773,N29774,N29775,N29776,N29777,N29778,
N29779,N29780,N29781,N29782,N29783,N29784,N29785,N29786,N29787,N29788,
N29789,N29790,N29791,N29792,N29793,N29794,N29795,N29796,N29797,N29798,
N29799,N29800,N29801,N29802,N29803,N29804,N29805,N29806,N29807,N29808,
N29809,N29810,N29811,N29812,N29813,N29814,N29815,N29816,N29817,N29818,
N29819,N29820,N29821,N29822,N29823,N29824,N29825,N29826,N29827,N29828,
N29829,N29830,N29831,N29832,N29833,N29834,N29835,N29836,N29837,N29838,
N29839,N29840,N29841,N29842,N29843,N29844,N29845,N29846,N29847,N29848,
N29849,N29850,N29851,N29852,N29853,N29854,N29855,N29856,N29857,N29858,
N29859,N29860,N29861,N29862,N29863,N29864,N29865,N29866,N29867,N29868,
N29869,N29870,N29871,N29872,N29873,N29874,N29875,N29876,N29877,N29878,
N29879,N29880,N29881,N29882,N29883,N29884,N29885,N29886,N29887,N29888,
N29889,N29890,N29891,N29892,N29893,N29894,N29895,N29896,N29897,N29898,
N29899,N29900,N29901,N29902,N29903,N29904,N29905,N29906,N29907,N29908,
N29909,N29910,N29911,N29912,N29913,N29914,N29915,N29916,N29917,N29918,
N29919,N29920,N29921,N29922,N29923,N29924,N29925,N29926,N29927,N29928,
N29929,N29930,N29931,N29932,N29933,N29934,N29935,N29936,N29937,N29938,
N29939,N29940,N29941,N29942,N29943,N29944,N29945,N29946,N29947,N29948,
N29949,N29950,N29951,N29952,N29953,N29954,N29955,N29956,N29957,N29958,
N29959,N29960,N29961,N29962,N29963,N29964,N29965,N29966,N29967,N29968,
N29969,N29970,N29971,N29972,N29973,N29974,N29975,N29976,N29977,N29978,
N29979,N29980,N29981,N29982,N29983,N29984,N29985,N29986,N29987,N29988,
N29989,N29990,N29991,N29992,N29993,N29994,N29995,N29996,N29997,N29998,
N29999,N30000,N30001,N30002,N30003,N30004,N30005,N30006,N30007,N30008,
N30009,N30010,N30011,N30012,N30013,N30014,N30015,N30016,N30017,N30018,
N30019,N30020,N30021,N30022,N30023,N30024,N30025,N30026,N30027,N30028,
N30029,N30030,N30031,N30032,N30033,N30034,N30035,N30036,N30037,N30038,
N30039,N30040,N30041,N30042,N30043,N30044,N30045,N30046,N30047,N30048,
N30049,N30050,N30051,N30052,N30053,N30054,N30055,N30056,N30057,N30058,
N30059,N30060,N30061,N30062,N30063,N30064,N30065,N30066,N30067,N30068,
N30069,N30070,N30071,N30072,N30073,N30074,N30075,N30076,N30077,N30078,
N30079,N30080,N30081,N30082,N30083,N30084,N30085,N30086,N30087,N30088,
N30089,N30090,N30091,N30092,N30093,N30094,N30095,N30096,N30097,N30098,
N30099,N30100,N30101,N30102,N30103,N30104,N30105,N30106,N30107,N30108,
N30109,N30110,N30111,N30112,N30113,N30114,N30115,N30116,N30117,N30118,
N30119,N30120,N30121,N30122,N30123,N30124,N30125,N30126,N30127,N30128,
N30129,N30130,N30131,N30132,N30133,N30134,N30135,N30136,N30137,N30138,
N30139,N30140,N30141,N30142,N30143,N30144,N30145,N30146,N30147,N30148,
N30149,N30150,N30151,N30152,N30153,N30154,N30155,N30156,N30157,N30158,
N30159,N30160,N30161,N30162,N30163,N30164,N30165,N30166,N30167,N30168,
N30169,N30170,N30171,N30172,N30173,N30174,N30175,N30176,N30177,N30178,
N30179,N30180,N30181,N30182,N30183,N30184,N30185,N30186,N30187,N30188,
N30189,N30190,N30191,N30192,N30193,N30194,N30195,N30196,N30197,N30198,
N30199,N30200,N30201,N30202,N30203,N30204,N30205,N30206,N30207,N30208,
N30209,N30210,N30211,N30212,N30213,N30214,N30215,N30216,N30217,N30218,
N30219,N30220,N30221,N30222,N30223,N30224,N30225,N30226,N30227,N30228,
N30229,N30230,N30231,N30232,N30233,N30234,N30235,N30236,N30237,N30238,
N30239,N30240,N30241,N30242,N30243,N30244,N30245,N30246,N30247,N30248,
N30249,N30250,N30251,N30252,N30253,N30254,N30255,N30256,N30257,N30258,
N30259,N30260,N30261,N30262,N30263,N30264,N30265,N30266,N30267,N30268,
N30269,N30270,N30271,N30272,N30273,N30274,N30275,N30276,N30277,N30278,
N30279,N30280,N30281,N30282,N30283,N30284,N30285,N30286,N30287,N30288,
N30289,N30290,N30291,N30292,N30293,N30294,N30295,N30296,N30297,N30298,
N30299,N30300,N30301,N30302,N30303,N30304,N30305,N30306,N30307,N30308,
N30309,N30310,N30311,N30312,N30313,N30314,N30315,N30316,N30317,N30318,
N30319,N30320,N30321,N30322,N30323,N30324,N30325,N30326,N30327,N30328,
N30329,N30330,N30331,N30332,N30333,N30334,N30335,N30336,N30337,N30338,
N30339,N30340,N30341,N30342,N30343,N30344,N30345,N30346,N30347,N30348,
N30349,N30350,N30351,N30352,N30353,N30354,N30355,N30356,N30357,N30358,
N30359,N30360,N30361,N30362,N30363,N30364,N30365,N30366,N30367,N30368,
N30369,N30370,N30371,N30372,N30373,N30374,N30375,N30376,N30377,N30378,
N30379,N30380,N30381,N30382,N30383,N30384,N30385,N30386,N30387,N30388,
N30389,N30390,N30391,N30392,N30393,N30394,N30395,N30396,N30397,N30398,
N30399,N30400,N30401,N30402,N30403,N30404,N30405,N30406,N30407,N30408,
N30409,N30410,N30411,N30412,N30413,N30414,N30415,N30416,N30417,N30418,
N30419,N30420,N30421,N30422,N30423,N30424,N30425,N30426,N30427,N30428,
N30429,N30430,N30431,N30432,N30433,N30434,N30435,N30436,N30437,N30438,
N30439,N30440,N30441,N30442,N30443,N30444,N30445,N30446,N30447,N30448,
N30449,N30450,N30451,N30452,N30453,N30454,N30455,N30456,N30457,N30458,
N30459,N30460,N30461,N30462,N30463,N30464,N30465,N30466,N30467,N30468,
N30469,N30470,N30471,N30472,N30473,N30474,N30475,N30476,N30477,N30478,
N30479,N30480,N30481,N30482,N30483,N30484,N30485,N30486,N30487,N30488,
N30489,N30490,N30491,N30492,N30493,N30494,N30495,N30496,N30497,N30498,
N30499,N30500,N30501,N30502,N30503,N30504,N30505,N30506,N30507,N30508,
N30509,N30510,N30511,N30512,N30513,N30514,N30515,N30516,N30517,N30518,
N30519,N30520,N30521,N30522,N30523,N30524,N30525,N30526,N30527,N30528,
N30529,N30530,N30531,N30532,N30533,N30534,N30535,N30536,N30537,N30538,
N30539,N30540,N30541,N30542,N30543,N30544,N30545,N30546,N30547,N30548,
N30549,N30550,N30551,N30552,N30553,N30554,N30555,N30556,N30557,N30558,
N30559,N30560,N30561,N30562,N30563,N30564,N30565,N30566,N30567,N30568,
N30569,N30570,N30571,N30572,N30573,N30574,N30575,N30576,N30577,N30578,
N30579,N30580,N30581,N30582,N30583,N30584,N30585,N30586,N30587,N30588,
N30589,N30590,N30591,N30592,N30593,N30594,N30595,N30596,N30597,N30598,
N30599,N30600,N30601,N30602,N30603,N30604,N30605,N30606,N30607,N30608,
N30609,N30610,N30611,N30612,N30613,N30614,N30615,N30616,N30617,N30618,
N30619,N30620,N30621,N30622,N30623,N30624,N30625,N30626,N30627,N30628,
N30629,N30630,N30631,N30632,N30633,N30634,N30635,N30636,N30637,N30638,
N30639,N30640,N30641,N30642,N30643,N30644,N30645,N30646,N30647,N30648,
N30649,N30650,N30651,N30652,N30653,N30654,N30655,N30656,N30657,N30658,
N30659,N30660,N30661,N30662,N30663,N30664,N30665,N30666,N30667,N30668,
N30669,N30670,N30671,N30672,N30673,N30674,N30675,N30676,N30677,N30678,
N30679,N30680,N30681,N30682,N30683,N30684,N30685,N30686,N30687,N30688,
N30689,N30690,N30691,N30692,N30693,N30694,N30695,N30696,N30697,N30698,
N30699,N30700,N30701,N30702,N30703,N30704,N30705,N30706,N30707,N30708,
N30709,N30710,N30711,N30712,N30713,N30714,N30715,N30716,N30717,N30718,
N30719,N30720,N30721,N30722,N30723,N30724,N30725,N30726,N30727,N30728,
N30729,N30730,N30731,N30732,N30733,N30734,N30735,N30736,N30737,N30738,
N30739,N30740,N30741,N30742,N30743,N30744,N30745,N30746,N30747,N30748,
N30749,N30750,N30751,N30752,N30753,N30754,N30755,N30756,N30757,N30758,
N30759,N30760,N30761,N30762,N30763,N30764,N30765,N30766,N30767,N30768,
N30769,N30770,N30771,N30772,N30773,N30774,N30775,N30776,N30777,N30778,
N30779,N30780,N30781,N30782,N30783,N30784,N30785,N30786,N30787,N30788,
N30789,N30790,N30791,N30792,N30793,N30794,N30795,N30796,N30797,N30798,
N30799,N30800,N30801,N30802,N30803,N30804,N30805,N30806,N30807,N30808,
N30809,N30810,N30811,N30812,N30813,N30814,N30815,N30816,N30817,N30818,
N30819,N30820,N30821,N30822,N30823,N30824,N30825,N30826,N30827,N30828,
N30829,N30830,N30831,N30832,N30833,N30834,N30835,N30836,N30837,N30838,
N30839,N30840,N30841,N30842,N30843,N30844,N30845,N30846,N30847,N30848,
N30849,N30850,N30851,N30852,N30853,N30854,N30855,N30856,N30857,N30858,
N30859,N30860,N30861,N30862,N30863,N30864,N30865,N30866,N30867,N30868,
N30869,N30870,N30871,N30872,N30873,N30874,N30875,N30876,N30877,N30878,
N30879,N30880,N30881,N30882,N30883,N30884,N30885,N30886,N30887,N30888,
N30889,N30890,N30891,N30892,N30893,N30894,N30895,N30896,N30897,N30898,
N30899,N30900,N30901,N30902,N30903,N30904,N30905,N30906,N30907,N30908,
N30909,N30910,N30911,N30912,N30913,N30914,N30915,N30916,N30917,N30918,
N30919,N30920,N30921,N30922,N30923,N30924,N30925,N30926,N30927,N30928,
N30929,N30930,N30931,N30932,N30933,N30934,N30935,N30936,N30937,N30938,
N30939,N30940,N30941,N30942,N30943,N30944,N30945,N30946,N30947,N30948,
N30949,N30950,N30951,N30952,N30953,N30954,N30955,N30956,N30957,N30958,
N30959,N30960,N30961,N30962,N30963,N30964,N30965,N30966,N30967,N30968,
N30969,N30970,N30971,N30972,N30973,N30974,N30975,N30976,N30977,N30978,
N30979,N30980,N30981,N30982,N30983,N30984,N30985,N30986,N30987,N30988,
N30989,N30990,N30991,N30992,N30993,N30994,N30995,N30996,N30997,N30998,
N30999,N31000,N31001,N31002,N31003,N31004,N31005,N31006,N31007,N31008,
N31009,N31010,N31011,N31012,N31013,N31014,N31015,N31016,N31017,N31018,
N31019,N31020,N31021,N31022,N31023,N31024,N31025,N31026,N31027,N31028,
N31029,N31030,N31031,N31032,N31033,N31034,N31035,N31036,N31037,N31038,
N31039,N31040,N31041,N31042,N31043,N31044,N31045,N31046,N31047,N31048,
N31049,N31050,N31051,N31052,N31053,N31054,N31055,N31056,N31057,N31058,
N31059,N31060,N31061,N31062,N31063,N31064,N31065,N31066,N31067,N31068,
N31069,N31070,N31071,N31072,N31073,N31074,N31075,N31076,N31077,N31078,
N31079,N31080,N31081,N31082,N31083,N31084,N31085,N31086,N31087,N31088,
N31089,N31090,N31091,N31092,N31093,N31094,N31095,N31096,N31097,N31098,
N31099,N31100,N31101,N31102,N31103,N31104,N31105,N31106,N31107,N31108,
N31109,N31110,N31111,N31112,N31113,N31114,N31115,N31116,N31117,N31118,
N31119,N31120,N31121,N31122,N31123,N31124,N31125,N31126,N31127,N31128,
N31129,N31130,N31131,N31132,N31133,N31134,N31135,N31136,N31137,N31138,
N31139,N31140,N31141,N31142,N31143,N31144,N31145,N31146,N31147,N31148,
N31149,N31150,N31151,N31152,N31153,N31154,N31155,N31156,N31157,N31158,
N31159,N31160,N31161,N31162,N31163,N31164,N31165,N31166,N31167,N31168,
N31169,N31170,N31171,N31172,N31173,N31174,N31175,N31176,N31177,N31178,
N31179,N31180,N31181,N31182,N31183,N31184,N31185,N31186,N31187,N31188,
N31189,N31190,N31191,N31192,N31193,N31194,N31195,N31196,N31197,N31198,
N31199,N31200,N31201,N31202,N31203,N31204,N31205,N31206,N31207,N31208,
N31209,N31210,N31211,N31212,N31213,N31214,N31215,N31216,N31217,N31218,
N31219,N31220,N31221,N31222,N31223,N31224,N31225,N31226,N31227,N31228,
N31229,N31230,N31231,N31232,N31233,N31234,N31235,N31236,N31237,N31238,
N31239,N31240,N31241,N31242,N31243,N31244,N31245,N31246,N31247,N31248,
N31249,N31250,N31251,N31252,N31253,N31254,N31255,N31256,N31257,N31258,
N31259,N31260,N31261,N31262,N31263,N31264,N31265,N31266,N31267,N31268,
N31269,N31270,N31271,N31272,N31273,N31274,N31275,N31276,N31277,N31278,
N31279,N31280,N31281,N31282,N31283,N31284,N31285,N31286,N31287,N31288,
N31289,N31290,N31291,N31292,N31293,N31294,N31295,N31296,N31297,N31298,
N31299,N31300,N31301,N31302,N31303,N31304,N31305,N31306,N31307,N31308,
N31309,N31310,N31311,N31312,N31313,N31314,N31315,N31316,N31317,N31318,
N31319,N31320,N31321,N31322,N31323,N31324,N31325,N31326,N31327,N31328,
N31329,N31330,N31331,N31332,N31333,N31334,N31335,N31336,N31337,N31338,
N31339,N31340,N31341,N31342,N31343,N31344,N31345,N31346,N31347,N31348,
N31349,N31350,N31351,N31352,N31353,N31354,N31355,N31356,N31357,N31358,
N31359,N31360,N31361,N31362,N31363,N31364,N31365,N31366,N31367,N31368,
N31369,N31370,N31371,N31372,N31373,N31374,N31375,N31376,N31377,N31378,
N31379,N31380,N31381,N31382,N31383,N31384,N31385,N31386,N31387,N31388,
N31389,N31390,N31391,N31392,N31393,N31394,N31395,N31396,N31397,N31398,
N31399,N31400,N31401,N31402,N31403,N31404,N31405,N31406,N31407,N31408,
N31409,N31410,N31411,N31412,N31413,N31414,N31415,N31416,N31417,N31418,
N31419,N31420,N31421,N31422,N31423,N31424,N31425,N31426,N31427,N31428,
N31429,N31430,N31431,N31432,N31433,N31434,N31435,N31436,N31437,N31438,
N31439,N31440,N31441,N31442,N31443,N31444,N31445,N31446,N31447,N31448,
N31449,N31450,N31451,N31452,N31453,N31454,N31455,N31456,N31457,N31458,
N31459,N31460,N31461,N31462,N31463,N31464,N31465,N31466,N31467,N31468,
N31469,N31470,N31471,N31472,N31473,N31474,N31475,N31476,N31477,N31478,
N31479,N31480,N31481,N31482,N31483,N31484,N31485,N31486,N31487,N31488,
N31489,N31490,N31491,N31492,N31493,N31494,N31495,N31496,N31497,N31498,
N31499,N31500,N31501,N31502,N31503,N31504,N31505,N31506,N31507,N31508,
N31509,N31510,N31511,N31512,N31513,N31514,N31515,N31516,N31517,N31518,
N31519,N31520,N31521,N31522,N31523,N31524,N31525,N31526,N31527,N31528,
N31529,N31530,N31531,N31532,N31533,N31534,N31535,N31536,N31537,N31538,
N31539,N31540,N31541,N31542,N31543,N31544,N31545,N31546,N31547,N31548,
N31549,N31550,N31551,N31552,N31553,N31554,N31555,N31556,N31557,N31558,
N31559,N31560,N31561,N31562,N31563,N31564,N31565,N31566,N31567,N31568,
N31569,N31570,N31571,N31572,N31573,N31574,N31575,N31576,N31577,N31578,
N31579,N31580,N31581,N31582,N31583,N31584,N31585,N31586,N31587,N31588,
N31589,N31590,N31591,N31592,N31593,N31594,N31595,N31596,N31597,N31598,
N31599,N31600,N31601,N31602,N31603,N31604,N31605,N31606,N31607,N31608,
N31609,N31610,N31611,N31612,N31613,N31614,N31615,N31616,N31617,N31618,
N31619,N31620,N31621,N31622,N31623,N31624,N31625,N31626,N31627,N31628,
N31629,N31630,N31631,N31632,N31633,N31634,N31635,N31636,N31637,N31638,
N31639,N31640,N31641,N31642,N31643,N31644,N31645,N31646,N31647,N31648,
N31649,N31650,N31651,N31652,N31653,N31654,N31655,N31656,N31657,N31658,
N31659,N31660,N31661,N31662,N31663,N31664,N31665,N31666,N31667,N31668,
N31669,N31670,N31671,N31672,N31673,N31674,N31675,N31676,N31677,N31678,
N31679,N31680,N31681,N31682,N31683,N31684,N31685,N31686,N31687,N31688,
N31689,N31690,N31691,N31692,N31693,N31694,N31695,N31696,N31697,N31698,
N31699,N31700,N31701,N31702,N31703,N31704,N31705,N31706,N31707,N31708,
N31709,N31710,N31711,N31712,N31713,N31714,N31715,N31716,N31717,N31718,
N31719,N31720,N31721,N31722,N31723,N31724,N31725,N31726,N31727,N31728,
N31729,N31730,N31731,N31732,N31733,N31734,N31735,N31736,N31737,N31738,
N31739,N31740,N31741,N31742,N31743,N31744,N31745,N31746,N31747,N31748,
N31749,N31750,N31751,N31752,N31753,N31754,N31755,N31756,N31757,N31758,
N31759,N31760,N31761,N31762,N31763,N31764,N31765,N31766,N31767,N31768,
N31769,N31770,N31771,N31772,N31773,N31774,N31775,N31776,N31777,N31778,
N31779,N31780,N31781,N31782,N31783,N31784,N31785,N31786,N31787,N31788,
N31789,N31790,N31791,N31792,N31793,N31794,N31795,N31796,N31797,N31798,
N31799,N31800,N31801,N31802,N31803,N31804,N31805,N31806,N31807,N31808,
N31809,N31810,N31811,N31812,N31813,N31814,N31815,N31816,N31817,N31818,
N31819,N31820,N31821,N31822,N31823,N31824,N31825,N31826,N31827,N31828,
N31829,N31830,N31831,N31832,N31833,N31834,N31835,N31836,N31837,N31838,
N31839,N31840,N31841,N31842,N31843,N31844,N31845,N31846,N31847,N31848,
N31849,N31850,N31851,N31852,N31853,N31854,N31855,N31856,N31857,N31858,
N31859,N31860,N31861,N31862,N31863,N31864,N31865,N31866,N31867,N31868,
N31869,N31870,N31871,N31872,N31873,N31874,N31875,N31876,N31877,N31878,
N31879,N31880,N31881,N31882,N31883,N31884,N31885,N31886,N31887,N31888,
N31889,N31890,N31891,N31892,N31893,N31894,N31895,N31896,N31897,N31898,
N31899,N31900,N31901,N31902,N31903,N31904,N31905,N31906,N31907,N31908,
N31909,N31910,N31911,N31912,N31913,N31914,N31915,N31916,N31917,N31918,
N31919,N31920,N31921,N31922,N31923,N31924,N31925,N31926,N31927,N31928,
N31929,N31930,N31931,N31932,N31933,N31934,N31935,N31936,N31937,N31938,
N31939,N31940,N31941,N31942,N31943,N31944,N31945,N31946,N31947,N31948,
N31949,N31950,N31951,N31952,N31953,N31954,N31955,N31956,N31957,N31958,
N31959,N31960,N31961,N31962,N31963,N31964,N31965,N31966,N31967,N31968,
N31969,N31970,N31971,N31972,N31973,N31974,N31975,N31976,N31977,N31978,
N31979,N31980,N31981,N31982,N31983,N31984,N31985,N31986,N31987,N31988,
N31989,N31990,N31991,N31992,N31993,N31994,N31995,N31996,N31997,N31998,
N31999,N32000,N32001,N32002,N32003,N32004,N32005,N32006,N32007,N32008,
N32009,N32010,N32011,N32012,N32013,N32014,N32015,N32016,N32017,N32018,
N32019,N32020,N32021,N32022,N32023,N32024,N32025,N32026,N32027,N32028,
N32029,N32030,N32031,N32032,N32033,N32034,N32035,N32036,N32037,N32038,
N32039,N32040,N32041,N32042,N32043,N32044,N32045,N32046,N32047,N32048,
N32049,N32050,N32051,N32052,N32053,N32054,N32055,N32056,N32057,N32058,
N32059,N32060,N32061,N32062,N32063,N32064,N32065,N32066,N32067,N32068,
N32069,N32070,N32071,N32072,N32073,N32074,N32075,N32076,N32077,N32078,
N32079,N32080,N32081,N32082,N32083,N32084,N32085,N32086,N32087,N32088,
N32089,N32090,N32091,N32092,N32093,N32094,N32095,N32096,N32097,N32098,
N32099,N32100,N32101,N32102,N32103,N32104,N32105,N32106,N32107,N32108,
N32109,N32110,N32111,N32112,N32113,N32114,N32115,N32116,N32117,N32118,
N32119,N32120,N32121,N32122,N32123,N32124,N32125,N32126,N32127,N32128,
N32129,N32130,N32131,N32132,N32133,N32134,N32135,N32136,N32137,N32138,
N32139,N32140,N32141,N32142,N32143,N32144,N32145,N32146,N32147,N32148,
N32149,N32150,N32151,N32152,N32153,N32154,N32155,N32156,N32157,N32158,
N32159,N32160,N32161,N32162,N32163,N32164,N32165,N32166,N32167,N32168,
N32169,N32170,N32171,N32172,N32173,N32174,N32175,N32176,N32177,N32178,
N32179,N32180,N32181,N32182,N32183,N32184,N32185,N32186,N32187,N32188,
N32189,N32190,N32191,N32192,N32193,N32194,N32195,N32196,N32197,N32198,
N32199,N32200,N32201,N32202,N32203,N32204,N32205,N32206,N32207,N32208,
N32209,N32210,N32211,N32212,N32213,N32214,N32215,N32216,N32217,N32218,
N32219,N32220,N32221,N32222,N32223,N32224,N32225,N32226,N32227,N32228,
N32229,N32230,N32231,N32232,N32233,N32234,N32235,N32236,N32237,N32238,
N32239,N32240,N32241,N32242,N32243,N32244,N32245,N32246,N32247,N32248,
N32249,N32250,N32251,N32252,N32253,N32254,N32255,N32256,N32257,N32258,
N32259,N32260,N32261,N32262,N32263,N32264,N32265,N32266,N32267,N32268,
N32269,N32270,N32271,N32272,N32273,N32274,N32275,N32276,N32277,N32278,
N32279,N32280,N32281,N32282,N32283,N32284,N32285,N32286,N32287,N32288,
N32289,N32290,N32291,N32292,N32293,N32294,N32295,N32296,N32297,N32298,
N32299,N32300,N32301,N32302,N32303,N32304,N32305,N32306,N32307,N32308,
N32309,N32310,N32311,N32312,N32313,N32314,N32315,N32316,N32317,N32318,
N32319,N32320,N32321,N32322,N32323,N32324,N32325,N32326,N32327,N32328,
N32329,N32330,N32331,N32332,N32333,N32334,N32335,N32336,N32337,N32338,
N32339,N32340,N32341,N32342,N32343,N32344,N32345,N32346,N32347,N32348,
N32349,N32350,N32351,N32352,N32353,N32354,N32355,N32356,N32357,N32358,
N32359,N32360,N32361,N32362,N32363,N32364,N32365,N32366,N32367,N32368,
N32369,N32370,N32371,N32372,N32373,N32374,N32375,N32376,N32377,N32378,
N32379,N32380,N32381,N32382,N32383,N32384,N32385,N32386,N32387,N32388,
N32389,N32390,N32391,N32392,N32393,N32394,N32395,N32396,N32397,N32398,
N32399,N32400,N32401,N32402,N32403,N32404,N32405,N32406,N32407,N32408,
N32409,N32410,N32411,N32412,N32413,N32414,N32415,N32416,N32417,N32418,
N32419,N32420,N32421,N32422,N32423,N32424,N32425,N32426,N32427,N32428,
N32429,N32430,N32431,N32432,N32433,N32434,N32435,N32436,N32437,N32438,
N32439,N32440,N32441,N32442,N32443,N32444,N32445,N32446,N32447,N32448,
N32449,N32450,N32451,N32452,N32453,N32454,N32455,N32456,N32457,N32458,
N32459,N32460,N32461,N32462,N32463,N32464,N32465,N32466,N32467,N32468,
N32469,N32470,N32471,N32472,N32473,N32474,N32475,N32476,N32477,N32478,
N32479,N32480,N32481,N32482,N32483,N32484,N32485,N32486,N32487,N32488,
N32489,N32490,N32491,N32492,N32493,N32494,N32495,N32496,N32497,N32498,
N32499,N32500,N32501,N32502,N32503,N32504,N32505,N32506,N32507,N32508,
N32509,N32510,N32511,N32512,N32513,N32514,N32515,N32516,N32517,N32518,
N32519,N32520,N32521,N32522,N32523,N32524,N32525,N32526,N32527,N32528,
N32529,N32530,N32531,N32532,N32533,N32534,N32535,N32536,N32537,N32538,
N32539,N32540,N32541,N32542,N32543,N32544,N32545,N32546,N32547,N32548,
N32549,N32550,N32551,N32552,N32553,N32554,N32555,N32556,N32557,N32558,
N32559,N32560,N32561,N32562,N32563,N32564,N32565,N32566,N32567,N32568,
N32569,N32570,N32571,N32572,N32573,N32574,N32575,N32576,N32577,N32578,
N32579,N32580,N32581,N32582,N32583,N32584,N32585,N32586,N32587,N32588,
N32589,N32590,N32591,N32592,N32593,N32594,N32595,N32596,N32597,N32598,
N32599,N32600,N32601,N32602,N32603,N32604,N32605,N32606,N32607,N32608,
N32609,N32610,N32611,N32612,N32613,N32614,N32615,N32616,N32617,N32618,
N32619,N32620,N32621,N32622,N32623,N32624,N32625,N32626,N32627,N32628,
N32629,N32630,N32631,N32632,N32633,N32634,N32635,N32636,N32637,N32638,
N32639,N32640,N32641,N32642,N32643,N32644,N32645,N32646,N32647,N32648,
N32649,N32650,N32651,N32652,N32653,N32654,N32655,N32656,N32657,N32658,
N32659,N32660,N32661,N32662,N32663,N32664,N32665,N32666,N32667,N32668,
N32669,N32670,N32671,N32672,N32673,N32674,N32675,N32676,N32677,N32678,
N32679,N32680,N32681,N32682,N32683,N32684,N32685,N32686,N32687,N32688,
N32689,N32690,N32691,N32692,N32693,N32694,N32695,N32696,N32697,N32698,
N32699,N32700,N32701,N32702,N32703,N32704,N32705,N32706,N32707,N32708,
N32709,N32710,N32711,N32712,N32713,N32714,N32715,N32716,N32717,N32718,
N32719,N32720,N32721,N32722,N32723,N32724,N32725,N32726,N32727,N32728,
N32729,N32730,N32731,N32732,N32733,N32734,N32735,N32736,N32737,N32738,
N32739,N32740,N32741,N32742,N32743,N32744,N32745,N32746,N32747,N32748,
N32749,N32750,N32751,N32752,N32753,N32754,N32755,N32756,N32757,N32758,
N32759,N32760,N32761,N32762,N32763,N32764,N32765,N32766,N32767,N32768,
N32769,N32770,N32771,N32772,N32773,N32774,N32775,N32776,N32777,N32778,
N32779,N32780,N32781,N32782,N32783,N32784,N32785,N32786,N32787,N32788,
N32789,N32790,N32791,N32792,N32793,N32794,N32795,N32796,N32797,N32798,
N32799,N32800,N32801,N32802,N32803,N32804,N32805,N32806,N32807,N32808,
N32809,N32810,N32811,N32812,N32813,N32814,N32815,N32816,N32817,N32818,
N32819,N32820,N32821,N32822,N32823,N32824,N32825,N32826,N32827,N32828,
N32829,N32830,N32831,N32832,N32833,N32834,N32835,N32836,N32837,N32838,
N32839,N32840,N32841,N32842,N32843,N32844,N32845,N32846,N32847,N32848,
N32849,N32850,N32851,N32852,N32853,N32854,N32855,N32856,N32857,N32858,
N32859,N32860,N32861,N32862,N32863,N32864,N32865,N32866,N32867,N32868,
N32869,N32870,N32871,N32872,N32873,N32874,N32875,N32876,N32877,N32878,
N32879,N32880,N32881,N32882,N32883,N32884,N32885,N32886,N32887,N32888,
N32889,N32890,N32891,N32892,N32893,N32894,N32895,N32896,N32897,N32898,
N32899,N32900,N32901,N32902,N32903,N32904,N32905,N32906,N32907,N32908,
N32909,N32910,N32911,N32912,N32913,N32914,N32915,N32916,N32917,N32918,
N32919,N32920,N32921,N32922,N32923,N32924,N32925,N32926,N32927,N32928,
N32929,N32930,N32931,N32932,N32933,N32934,N32935,N32936,N32937,N32938,
N32939,N32940,N32941,N32942,N32943,N32944,N32945,N32946,N32947,N32948,
N32949,N32950,N32951,N32952,N32953,N32954,N32955,N32956,N32957,N32958,
N32959,N32960,N32961,N32962,N32963,N32964,N32965,N32966,N32967,N32968,
N32969,N32970,N32971,N32972,N32973,N32974,N32975,N32976,N32977,N32978,
N32979,N32980,N32981,N32982,N32983,N32984,N32985,N32986,N32987,N32988,
N32989,N32990,N32991,N32992,N32993,N32994,N32995,N32996,N32997,N32998,
N32999,N33000,N33001,N33002,N33003,N33004,N33005,N33006,N33007,N33008,
N33009,N33010,N33011,N33012,N33013,N33014,N33015,N33016,N33017,N33018,
N33019,N33020,N33021,N33022,N33023,N33024,N33025,N33026,N33027,N33028,
N33029,N33030,N33031,N33032,N33033,N33034,N33035,N33036,N33037,N33038,
N33039,N33040,N33041,N33042,N33043,N33044,N33045,N33046,N33047,N33048,
N33049,N33050,N33051,N33052,N33053,N33054,N33055,N33056,N33057,N33058,
N33059,N33060,N33061,N33062,N33063,N33064,N33065,N33066,N33067,N33068,
N33069,N33070,N33071,N33072,N33073,N33074,N33075,N33076,N33077,N33078,
N33079,N33080,N33081,N33082,N33083,N33084,N33085,N33086,N33087,N33088,
N33089,N33090,N33091,N33092,N33093,N33094,N33095,N33096,N33097,N33098,
N33099,N33100,N33101,N33102,N33103,N33104,N33105,N33106,N33107,N33108,
N33109,N33110,N33111,N33112,N33113,N33114,N33115,N33116,N33117,N33118,
N33119,N33120,N33121,N33122,N33123,N33124,N33125,N33126,N33127,N33128,
N33129,N33130,N33131,N33132,N33133,N33134,N33135,N33136,N33137,N33138,
N33139,N33140,N33141,N33142,N33143,N33144,N33145,N33146,N33147,N33148,
N33149,N33150,N33151,N33152,N33153,N33154,N33155,N33156,N33157,N33158,
N33159,N33160,N33161,N33162,N33163,N33164,N33165,N33166,N33167,N33168,
N33169,N33170,N33171,N33172,N33173,N33174,N33175,N33176,N33177,N33178,
N33179,N33180,N33181,N33182,N33183,N33184,N33185,N33186,N33187,N33188,
N33189,N33190,N33191,N33192,N33193,N33194,N33195,N33196,N33197,N33198,
N33199,N33200,N33201,N33202,N33203,N33204,N33205,N33206,N33207,N33208,
N33209,N33210,N33211,N33212,N33213,N33214,N33215,N33216,N33217,N33218,
N33219,N33220,N33221,N33222,N33223,N33224,N33225,N33226,N33227,N33228,
N33229,N33230,N33231,N33232,N33233,N33234,N33235,N33236,N33237,N33238,
N33239,N33240,N33241,N33242,N33243,N33244,N33245,N33246,N33247,N33248,
N33249,N33250,N33251,N33252,N33253,N33254,N33255,N33256,N33257,N33258,
N33259,N33260,N33261,N33262,N33263,N33264,N33265,N33266,N33267,N33268,
N33269,N33270,N33271,N33272,N33273,N33274,N33275,N33276,N33277,N33278,
N33279,N33280,N33281,N33282,N33283,N33284,N33285,N33286,N33287,N33288,
N33289,N33290,N33291,N33292,N33293,N33294,N33295,N33296,N33297,N33298,
N33299,N33300,N33301,N33302,N33303,N33304,N33305,N33306,N33307,N33308,
N33309,N33310,N33311,N33312,N33313,N33314,N33315,N33316,N33317,N33318,
N33319,N33320,N33321,N33322,N33323,N33324,N33325,N33326,N33327,N33328,
N33329,N33330,N33331,N33332,N33333,N33334,N33335,N33336,N33337,N33338,
N33339,N33340,N33341,N33342,N33343,N33344,N33345,N33346,N33347,N33348,
N33349,N33350,N33351,N33352,N33353,N33354,N33355,N33356,N33357,N33358,
N33359,N33360,N33361,N33362,N33363,N33364,N33365,N33366,N33367,N33368,
N33369,N33370,N33371,N33372,N33373,N33374,N33375,N33376,N33377,N33378,
N33379,N33380,N33381,N33382,N33383,N33384,N33385,N33386,N33387,N33388,
N33389,N33390,N33391,N33392,N33393,N33394,N33395,N33396,N33397,N33398,
N33399,N33400,N33401,N33402,N33403,N33404,N33405,N33406,N33407,N33408,
N33409,N33410,N33411,N33412,N33413,N33414,N33415,N33416,N33417,N33418,
N33419,N33420,N33421,N33422,N33423,N33424,N33425,N33426,N33427,N33428,
N33429,N33430,N33431,N33432,N33433,N33434,N33435,N33436,N33437,N33438,
N33439,N33440,N33441,N33442,N33443,N33444,N33445,N33446,N33447,N33448,
N33449,N33450,N33451,N33452,N33453,N33454,N33455,N33456,N33457,N33458,
N33459,N33460,N33461,N33462,N33463,N33464,N33465,N33466,N33467,N33468,
N33469,N33470,N33471,N33472,N33473,N33474,N33475,N33476,N33477,N33478,
N33479,N33480,N33481,N33482,N33483,N33484,N33485,N33486,N33487,N33488,
N33489,N33490,N33491,N33492,N33493,N33494,N33495,N33496,N33497,N33498,
N33499,N33500,N33501,N33502,N33503,N33504,N33505,N33506,N33507,N33508,
N33509,N33510,N33511,N33512,N33513,N33514,N33515,N33516,N33517,N33518,
N33519,N33520,N33521,N33522,N33523,N33524,N33525,N33526,N33527,N33528,
N33529,N33530,N33531,N33532,N33533,N33534,N33535,N33536,N33537,N33538,
N33539,N33540,N33541,N33542,N33543,N33544,N33545,N33546,N33547,N33548,
N33549,N33550,N33551,N33552,N33553,N33554,N33555,N33556,N33557,N33558,
N33559,N33560,N33561,N33562,N33563,N33564,N33565,N33566,N33567,N33568,
N33569,N33570,N33571,N33572,N33573,N33574,N33575,N33576,N33577,N33578,
N33579,N33580,N33581,N33582,N33583,N33584,N33585,N33586,N33587,N33588,
N33589,N33590,N33591,N33592,N33593,N33594,N33595,N33596,N33597,N33598,
N33599,N33600,N33601,N33602,N33603,N33604,N33605,N33606,N33607,N33608,
N33609,N33610,N33611,N33612,N33613,N33614,N33615,N33616,N33617,N33618,
N33619,N33620,N33621,N33622,N33623,N33624,N33625,N33626,N33627,N33628,
N33629,N33630,N33631,N33632,N33633,N33634,N33635,N33636,N33637,N33638,
N33639,N33640,N33641,N33642,N33643,N33644,N33645,N33646,N33647,N33648,
N33649,N33650,N33651,N33652,N33653,N33654,N33655,N33656,N33657,N33658,
N33659,N33660,N33661,N33662,N33663,N33664,N33665,N33666,N33667,N33668,
N33669,N33670,N33671,N33672,N33673,N33674,N33675,N33676,N33677,N33678,
N33679,N33680,N33681,N33682,N33683,N33684,N33685,N33686,N33687,N33688,
N33689,N33690,N33691,N33692,N33693,N33694,N33695,N33696,N33697,N33698,
N33699,N33700,N33701,N33702,N33703,N33704,N33705,N33706,N33707,N33708,
N33709,N33710,N33711,N33712,N33713,N33714,N33715,N33716,N33717,N33718,
N33719,N33720,N33721,N33722,N33723,N33724,N33725,N33726,N33727,N33728,
N33729,N33730,N33731,N33732,N33733,N33734,N33735,N33736,N33737,N33738,
N33739,N33740,N33741,N33742,N33743,N33744,N33745,N33746,N33747,N33748,
N33749,N33750,N33751,N33752,N33753,N33754,N33755,N33756,N33757,N33758,
N33759,N33760,N33761,N33762,N33763,N33764,N33765,N33766,N33767,N33768,
N33769,N33770,N33771,N33772,N33773,N33774,N33775,N33776,N33777,N33778,
N33779,N33780,N33781,N33782,N33783,N33784,N33785,N33786,N33787,N33788,
N33789,N33790,N33791,N33792,N33793,N33794,N33795,N33796,N33797,N33798,
N33799,N33800,N33801,N33802,N33803,N33804,N33805,N33806,N33807,N33808,
N33809,N33810,N33811,N33812,N33813,N33814,N33815,N33816,N33817,N33818,
N33819,N33820,N33821,N33822,N33823,N33824,N33825,N33826,N33827,N33828,
N33829,N33830,N33831,N33832,N33833,N33834,N33835,N33836,N33837,N33838,
N33839,N33840,N33841,N33842,N33843,N33844,N33845,N33846,N33847,N33848,
N33849,N33850,N33851,N33852,N33853,N33854,N33855,N33856,N33857,N33858,
N33859,N33860,N33861,N33862,N33863,N33864,N33865,N33866,N33867,N33868,
N33869,N33870,N33871,N33872,N33873,N33874,N33875,N33876,N33877,N33878,
N33879,N33880,N33881,N33882,N33883,N33884,N33885,N33886,N33887,N33888,
N33889,N33890,N33891,N33892,N33893,N33894,N33895,N33896,N33897,N33898,
N33899,N33900,N33901,N33902,N33903,N33904,N33905,N33906,N33907,N33908,
N33909,N33910,N33911,N33912,N33913,N33914,N33915,N33916,N33917,N33918,
N33919,N33920,N33921,N33922,N33923,N33924,N33925,N33926,N33927,N33928,
N33929,N33930,N33931,N33932,N33933,N33934,N33935,N33936,N33937,N33938,
N33939,N33940,N33941,N33942,N33943,N33944,N33945,N33946,N33947,N33948,
N33949,N33950,N33951,N33952,N33953,N33954,N33955,N33956,N33957,N33958,
N33959,N33960,N33961,N33962,N33963,N33964,N33965,N33966,N33967,N33968,
N33969,N33970,N33971,N33972,N33973,N33974,N33975,N33976,N33977,N33978,
N33979,N33980,N33981,N33982,N33983,N33984,N33985,N33986,N33987,N33988,
N33989,N33990,N33991,N33992,N33993,N33994,N33995,N33996,N33997,N33998,
N33999,N34000,N34001,N34002,N34003,N34004,N34005,N34006,N34007,N34008,
N34009,N34010,N34011,N34012,N34013,N34014,N34015,N34016,N34017,N34018,
N34019,N34020,N34021,N34022,N34023,N34024,N34025,N34026,N34027,N34028,
N34029,N34030,N34031,N34032,N34033,N34034,N34035,N34036,N34037,N34038,
N34039,N34040,N34041,N34042,N34043,N34044,N34045,N34046,N34047,N34048,
N34049,N34050,N34051,N34052,N34053,N34054,N34055,N34056,N34057,N34058,
N34059,N34060,N34061,N34062,N34063,N34064,N34065,N34066,N34067,N34068,
N34069,N34070,N34071,N34072,N34073,N34074,N34075,N34076,N34077,N34078,
N34079,N34080,N34081,N34082,N34083,N34084,N34085,N34086,N34087,N34088,
N34089,N34090,N34091,N34092,N34093,N34094,N34095,N34096,N34097,N34098,
N34099,N34100,N34101,N34102,N34103,N34104,N34105,N34106,N34107,N34108,
N34109,N34110,N34111,N34112,N34113,N34114,N34115,N34116,N34117,N34118,
N34119,N34120,N34121,N34122,N34123,N34124,N34125,N34126,N34127,N34128,
N34129,N34130,N34131,N34132,N34133,N34134,N34135,N34136,N34137,N34138,
N34139,N34140,N34141,N34142,N34143,N34144,N34145,N34146,N34147,N34148,
N34149,N34150,N34151,N34152,N34153,N34154,N34155,N34156,N34157,N34158,
N34159,N34160,N34161,N34162,N34163,N34164,N34165,N34166,N34167,N34168,
N34169,N34170,N34171,N34172,N34173,N34174,N34175,N34176,N34177,N34178,
N34179,N34180,N34181,N34182,N34183,N34184,N34185,N34186,N34187,N34188,
N34189,N34190,N34191,N34192,N34193,N34194,N34195,N34196,N34197,N34198,
N34199,N34200,N34201,N34202,N34203,N34204,N34205,N34206,N34207,N34208,
N34209,N34210,N34211,N34212,N34213,N34214,N34215,N34216,N34217,N34218,
N34219,N34220,N34221,N34222,N34223,N34224,N34225,N34226,N34227,N34228,
N34229,N34230,N34231,N34232,N34233,N34234,N34235,N34236,N34237,N34238,
N34239,N34240,N34241,N34242,N34243,N34244,N34245,N34246,N34247,N34248,
N34249,N34250,N34251,N34252,N34253,N34254,N34255,N34256,N34257,N34258,
N34259,N34260,N34261,N34262,N34263,N34264,N34265,N34266,N34267,N34268,
N34269,N34270,N34271,N34272,N34273,N34274,N34275,N34276,N34277,N34278,
N34279,N34280,N34281,N34282,N34283,N34284,N34285,N34286,N34287,N34288,
N34289,N34290,N34291,N34292,N34293,N34294,N34295,N34296,N34297,N34298,
N34299,N34300,N34301,N34302,N34303,N34304,N34305,N34306,N34307,N34308,
N34309,N34310,N34311,N34312,N34313,N34314,N34315,N34316,N34317,N34318,
N34319,N34320,N34321,N34322,N34323,N34324,N34325,N34326,N34327,N34328,
N34329,N34330,N34331,N34332,N34333,N34334,N34335,N34336,N34337,N34338,
N34339,N34340,N34341,N34342,N34343,N34344,N34345,N34346,N34347,N34348,
N34349,N34350,N34351,N34352,N34353,N34354,N34355,N34356,N34357,N34358,
N34359,N34360,N34361,N34362,N34363,N34364,N34365,N34366,N34367,N34368,
N34369,N34370,N34371,N34372,N34373,N34374,N34375,N34376,N34377,N34378,
N34379,N34380,N34381,N34382,N34383,N34384,N34385,N34386,N34387,N34388,
N34389,N34390,N34391,N34392,N34393,N34394,N34395,N34396,N34397,N34398,
N34399,N34400,N34401,N34402,N34403,N34404,N34405,N34406,N34407,N34408,
N34409,N34410,N34411,N34412,N34413,N34414,N34415,N34416,N34417,N34418,
N34419,N34420,N34421,N34422,N34423,N34424,N34425,N34426,N34427,N34428,
N34429,N34430,N34431,N34432,N34433,N34434,N34435,N34436,N34437,N34438,
N34439,N34440,N34441,N34442,N34443,N34444,N34445,N34446,N34447,N34448,
N34449,N34450,N34451,N34452,N34453,N34454,N34455,N34456,N34457,N34458,
N34459,N34460,N34461,N34462,N34463,N34464,N34465,N34466,N34467,N34468,
N34469,N34470,N34471,N34472,N34473,N34474,N34475,N34476,N34477,N34478,
N34479,N34480,N34481,N34482,N34483,N34484,N34485,N34486,N34487,N34488,
N34489,N34490,N34491,N34492,N34493,N34494,N34495,N34496,N34497,N34498,
N34499,N34500,N34501,N34502,N34503,N34504,N34505,N34506,N34507,N34508,
N34509,N34510,N34511,N34512,N34513,N34514,N34515,N34516,N34517,N34518,
N34519,N34520,N34521,N34522,N34523,N34524,N34525,N34526,N34527,N34528,
N34529,N34530,N34531,N34532,N34533,N34534,N34535,N34536,N34537,N34538,
N34539,N34540,N34541,N34542,N34543,N34544,N34545,N34546,N34547,N34548,
N34549,N34550,N34551,N34552,N34553,N34554,N34555,N34556,N34557,N34558,
N34559,N34560,N34561,N34562,N34563,N34564,N34565,N34566,N34567,N34568,
N34569,N34570,N34571,N34572,N34573,N34574,N34575,N34576,N34577,N34578,
N34579,N34580,N34581,N34582,N34583,N34584,N34585,N34586,N34587,N34588,
N34589,N34590,N34591,N34592,N34593,N34594,N34595,N34596,N34597,N34598,
N34599,N34600,N34601,N34602,N34603,N34604,N34605,N34606,N34607,N34608,
N34609,N34610,N34611,N34612,N34613,N34614,N34615,N34616,N34617,N34618,
N34619,N34620,N34621,N34622,N34623,N34624,N34625,N34626,N34627,N34628,
N34629,N34630,N34631,N34632,N34633,N34634,N34635,N34636,N34637,N34638,
N34639,N34640,N34641,N34642,N34643,N34644,N34645,N34646,N34647,N34648,
N34649,N34650,N34651,N34652,N34653,N34654,N34655,N34656,N34657,N34658,
N34659,N34660,N34661,N34662,N34663,N34664,N34665,N34666,N34667,N34668,
N34669,N34670,N34671,N34672,N34673,N34674,N34675,N34676,N34677,N34678,
N34679,N34680,N34681,N34682,N34683,N34684,N34685,N34686,N34687,N34688,
N34689,N34690,N34691,N34692,N34693,N34694,N34695,N34696,N34697,N34698,
N34699,N34700,N34701,N34702,N34703,N34704,N34705,N34706,N34707,N34708,
N34709,N34710,N34711,N34712,N34713,N34714,N34715,N34716,N34717,N34718,
N34719,N34720,N34721,N34722,N34723,N34724,N34725,N34726,N34727,N34728,
N34729,N34730,N34731,N34732,N34733,N34734,N34735,N34736,N34737,N34738,
N34739,N34740,N34741,N34742,N34743,N34744,N34745,N34746,N34747,N34748,
N34749,N34750,N34751,N34752,N34753,N34754,N34755,N34756,N34757,N34758,
N34759,N34760,N34761,N34762,N34763,N34764,N34765,N34766,N34767,N34768,
N34769,N34770,N34771,N34772,N34773,N34774,N34775,N34776,N34777,N34778,
N34779,N34780,N34781,N34782,N34783,N34784,N34785,N34786,N34787,N34788,
N34789,N34790,N34791,N34792,N34793,N34794,N34795,N34796,N34797,N34798,
N34799,N34800,N34801,N34802,N34803,N34804,N34805,N34806,N34807,N34808,
N34809,N34810,N34811,N34812,N34813,N34814,N34815,N34816,N34817,N34818,
N34819,N34820,N34821,N34822,N34823,N34824,N34825,N34826,N34827,N34828,
N34829,N34830,N34831,N34832,N34833,N34834,N34835,N34836,N34837,N34838,
N34839,N34840,N34841,N34842,N34843,N34844,N34845,N34846,N34847,N34848,
N34849,N34850,N34851,N34852,N34853,N34854,N34855,N34856,N34857,N34858,
N34859,N34860,N34861,N34862,N34863,N34864,N34865,N34866,N34867,N34868,
N34869,N34870,N34871,N34872,N34873,N34874,N34875,N34876,N34877,N34878,
N34879,N34880,N34881,N34882,N34883,N34884,N34885,N34886,N34887,N34888,
N34889,N34890,N34891,N34892,N34893,N34894,N34895,N34896,N34897,N34898,
N34899,N34900,N34901,N34902,N34903,N34904,N34905,N34906,N34907,N34908,
N34909,N34910,N34911,N34912,N34913,N34914,N34915,N34916,N34917,N34918,
N34919,N34920,N34921,N34922,N34923,N34924,N34925,N34926,N34927,N34928,
N34929,N34930,N34931,N34932,N34933,N34934,N34935,N34936,N34937,N34938,
N34939,N34940,N34941,N34942,N34943,N34944,N34945,N34946,N34947,N34948,
N34949,N34950,N34951,N34952,N34953,N34954,N34955,N34956,N34957,N34958,
N34959,N34960,N34961,N34962,N34963,N34964,N34965,N34966,N34967,N34968,
N34969,N34970,N34971,N34972,N34973,N34974,N34975,N34976,N34977,N34978,
N34979,N34980,N34981,N34982,N34983,N34984,N34985,N34986,N34987,N34988,
N34989,N34990,N34991,N34992,N34993,N34994,N34995,N34996,N34997,N34998,
N34999,N35000,N35001,N35002,N35003,N35004,N35005,N35006,N35007,N35008,
N35009,N35010,N35011,N35012,N35013,N35014,N35015,N35016,N35017,N35018,
N35019,N35020,N35021,N35022,N35023,N35024,N35025,N35026,N35027,N35028,
N35029,N35030,N35031,N35032,N35033,N35034,N35035,N35036,N35037,N35038,
N35039,N35040,N35041,N35042,N35043,N35044,N35045,N35046,N35047,N35048,
N35049,N35050,N35051,N35052,N35053,N35054,N35055,N35056,N35057,N35058,
N35059,N35060,N35061,N35062,N35063,N35064,N35065,N35066,N35067,N35068,
N35069,N35070,N35071,N35072,N35073,N35074,N35075,N35076,N35077,N35078,
N35079,N35080,N35081,N35082,N35083,N35084,N35085,N35086,N35087,N35088,
N35089,N35090,N35091,N35092,N35093,N35094,N35095,N35096,N35097,N35098,
N35099,N35100,N35101,N35102,N35103,N35104,N35105,N35106,N35107,N35108,
N35109,N35110,N35111,N35112,N35113,N35114,N35115,N35116,N35117,N35118,
N35119,N35120,N35121,N35122,N35123,N35124,N35125,N35126,N35127,N35128,
N35129,N35130,N35131,N35132,N35133,N35134,N35135,N35136,N35137,N35138,
N35139,N35140,N35141,N35142,N35143,N35144,N35145,N35146,N35147,N35148,
N35149,N35150,N35151,N35152,N35153,N35154,N35155,N35156,N35157,N35158,
N35159,N35160,N35161,N35162,N35163,N35164,N35165,N35166,N35167,N35168,
N35169,N35170,N35171,N35172,N35173,N35174,N35175,N35176,N35177,N35178,
N35179,N35180,N35181,N35182,N35183,N35184,N35185,N35186,N35187,N35188,
N35189,N35190,N35191,N35192,N35193,N35194,N35195,N35196,N35197,N35198,
N35199,N35200,N35201,N35202,N35203,N35204,N35205,N35206,N35207,N35208,
N35209,N35210,N35211,N35212,N35213,N35214,N35215,N35216,N35217,N35218,
N35219,N35220,N35221,N35222,N35223,N35224,N35225,N35226,N35227,N35228,
N35229,N35230,N35231,N35232,N35233,N35234,N35235,N35236,N35237,N35238,
N35239,N35240,N35241,N35242,N35243,N35244,N35245,N35246,N35247,N35248,
N35249,N35250,N35251,N35252,N35253,N35254,N35255,N35256,N35257,N35258,
N35259,N35260,N35261,N35262,N35263,N35264,N35265,N35266,N35267,N35268,
N35269,N35270,N35271,N35272,N35273,N35274,N35275,N35276,N35277,N35278,
N35279,N35280,N35281,N35282,N35283,N35284,N35285,N35286,N35287,N35288,
N35289,N35290,N35291,N35292,N35293,N35294,N35295,N35296,N35297,N35298,
N35299,N35300,N35301,N35302,N35303,N35304,N35305,N35306,N35307,N35308,
N35309,N35310,N35311,N35312,N35313,N35314,N35315,N35316,N35317,N35318,
N35319,N35320,N35321,N35322,N35323,N35324,N35325,N35326,N35327,N35328,
N35329,N35330,N35331,N35332,N35333,N35334,N35335,N35336,N35337,N35338,
N35339,N35340,N35341,N35342,N35343,N35344,N35345,N35346,N35347,N35348,
N35349,N35350,N35351,N35352,N35353,N35354,N35355,N35356,N35357,N35358,
N35359,N35360,N35361,N35362,N35363,N35364,N35365,N35366,N35367,N35368,
N35369,N35370,N35371,N35372,N35373,N35374,N35375,N35376,N35377,N35378,
N35379,N35380,N35381,N35382,N35383,N35384,N35385,N35386,N35387,N35388,
N35389,N35390,N35391,N35392,N35393,N35394,N35395,N35396,N35397,N35398,
N35399,N35400,N35401,N35402,N35403,N35404,N35405,N35406,N35407,N35408,
N35409,N35410,N35411,N35412,N35413,N35414,N35415,N35416,N35417,N35418,
N35419,N35420,N35421,N35422,N35423,N35424,N35425,N35426,N35427,N35428,
N35429,N35430,N35431,N35432,N35433,N35434,N35435,N35436,N35437,N35438,
N35439,N35440,N35441,N35442,N35443,N35444,N35445,N35446,N35447,N35448,
N35449,N35450,N35451,N35452,N35453,N35454,N35455,N35456,N35457,N35458,
N35459,N35460,N35461,N35462,N35463,N35464,N35465,N35466,N35467,N35468,
N35469,N35470,N35471,N35472,N35473,N35474,N35475,N35476,N35477,N35478,
N35479,N35480,N35481,N35482,N35483,N35484,N35485,N35486,N35487,N35488,
N35489,N35490,N35491,N35492,N35493,N35494,N35495,N35496,N35497,N35498,
N35499,N35500,N35501,N35502,N35503,N35504,N35505,N35506,N35507,N35508,
N35509,N35510,N35511,N35512,N35513,N35514,N35515,N35516,N35517,N35518,
N35519,N35520,N35521,N35522,N35523,N35524,N35525,N35526,N35527,N35528,
N35529,N35530,N35531,N35532,N35533,N35534,N35535,N35536,N35537,N35538,
N35539,N35540,N35541,N35542,N35543,N35544,N35545,N35546,N35547,N35548,
N35549,N35550,N35551,N35552,N35553,N35554,N35555,N35556,N35557,N35558,
N35559,N35560,N35561,N35562,N35563,N35564,N35565,N35566,N35567,N35568,
N35569,N35570,N35571,N35572,N35573,N35574,N35575,N35576,N35577,N35578,
N35579,N35580,N35581,N35582,N35583,N35584,N35585,N35586,N35587,N35588,
N35589,N35590,N35591,N35592,N35593,N35594,N35595,N35596,N35597,N35598,
N35599,N35600,N35601,N35602,N35603,N35604,N35605,N35606,N35607,N35608,
N35609,N35610,N35611,N35612,N35613,N35614,N35615,N35616,N35617,N35618,
N35619,N35620,N35621,N35622,N35623,N35624,N35625,N35626,N35627,N35628,
N35629,N35630,N35631,N35632,N35633,N35634,N35635,N35636,N35637,N35638,
N35639,N35640,N35641,N35642,N35643,N35644,N35645,N35646,N35647,N35648,
N35649,N35650,N35651,N35652,N35653,N35654,N35655,N35656,N35657,N35658,
N35659,N35660,N35661,N35662,N35663,N35664,N35665,N35666,N35667,N35668,
N35669,N35670,N35671,N35672,N35673,N35674,N35675,N35676,N35677,N35678,
N35679,N35680,N35681,N35682,N35683,N35684,N35685,N35686,N35687,N35688,
N35689,N35690,N35691,N35692,N35693,N35694,N35695,N35696,N35697,N35698,
N35699,N35700,N35701,N35702,N35703,N35704,N35705,N35706,N35707,N35708,
N35709,N35710,N35711,N35712,N35713,N35714,N35715,N35716,N35717,N35718,
N35719,N35720,N35721,N35722,N35723,N35724,N35725,N35726,N35727,N35728,
N35729,N35730,N35731,N35732,N35733,N35734,N35735,N35736,N35737,N35738,
N35739,N35740,N35741,N35742,N35743,N35744,N35745,N35746,N35747,N35748,
N35749,N35750,N35751,N35752,N35753,N35754,N35755,N35756,N35757,N35758,
N35759,N35760,N35761,N35762,N35763,N35764,N35765,N35766,N35767,N35768,
N35769,N35770,N35771,N35772,N35773,N35774,N35775,N35776,N35777,N35778,
N35779,N35780,N35781,N35782,N35783,N35784,N35785,N35786,N35787,N35788,
N35789,N35790,N35791,N35792,N35793,N35794,N35795,N35796,N35797,N35798,
N35799,N35800,N35801,N35802,N35803,N35804,N35805,N35806,N35807,N35808,
N35809,N35810,N35811,N35812,N35813,N35814,N35815,N35816,N35817,N35818,
N35819,N35820,N35821,N35822,N35823,N35824,N35825,N35826,N35827,N35828,
N35829,N35830,N35831,N35832,N35833,N35834,N35835,N35836,N35837,N35838,
N35839,N35840,N35841,N35842,N35843,N35844,N35845,N35846,N35847,N35848,
N35849,N35850,N35851,N35852,N35853,N35854,N35855,N35856,N35857,N35858,
N35859,N35860,N35861,N35862,N35863,N35864,N35865,N35866,N35867,N35868,
N35869,N35870,N35871,N35872,N35873,N35874,N35875,N35876,N35877,N35878,
N35879,N35880,N35881,N35882,N35883,N35884,N35885,N35886,N35887,N35888,
N35889,N35890,N35891,N35892,N35893,N35894,N35895,N35896,N35897,N35898,
N35899,N35900,N35901,N35902,N35903,N35904,N35905,N35906,N35907,N35908,
N35909,N35910,N35911,N35912,N35913,N35914,N35915,N35916,N35917,N35918,
N35919,N35920,N35921,N35922,N35923,N35924,N35925,N35926,N35927,N35928,
N35929,N35930,N35931,N35932,N35933,N35934,N35935,N35936,N35937,N35938,
N35939,N35940,N35941,N35942,N35943,N35944,N35945,N35946,N35947,N35948,
N35949,N35950,N35951,N35952,N35953,N35954,N35955,N35956,N35957,N35958,
N35959,N35960,N35961,N35962,N35963,N35964,N35965,N35966,N35967,N35968,
N35969,N35970,N35971,N35972,N35973,N35974,N35975,N35976,N35977,N35978,
N35979,N35980,N35981,N35982,N35983,N35984,N35985,N35986,N35987,N35988,
N35989,N35990,N35991,N35992,N35993,N35994,N35995,N35996,N35997,N35998,
N35999,N36000,N36001,N36002,N36003,N36004,N36005,N36006,N36007,N36008,
N36009,N36010,N36011,N36012,N36013,N36014,N36015,N36016,N36017,N36018,
N36019,N36020,N36021,N36022,N36023,N36024,N36025,N36026,N36027,N36028,
N36029,N36030,N36031,N36032,N36033,N36034,N36035,N36036,N36037,N36038,
N36039,N36040,N36041,N36042,N36043,N36044,N36045,N36046,N36047,N36048,
N36049,N36050,N36051,N36052,N36053,N36054,N36055,N36056,N36057,N36058,
N36059,N36060,N36061,N36062,N36063,N36064,N36065,N36066,N36067,N36068,
N36069,N36070,N36071,N36072,N36073,N36074,N36075,N36076,N36077,N36078,
N36079,N36080,N36081,N36082,N36083,N36084,N36085,N36086,N36087,N36088,
N36089,N36090,N36091,N36092,N36093,N36094,N36095,N36096,N36097,N36098,
N36099,N36100,N36101,N36102,N36103,N36104,N36105,N36106,N36107,N36108,
N36109,N36110,N36111,N36112,N36113,N36114,N36115,N36116,N36117,N36118,
N36119,N36120,N36121,N36122,N36123,N36124,N36125,N36126,N36127,N36128,
N36129,N36130,N36131,N36132,N36133,N36134,N36135,N36136,N36137,N36138,
N36139,N36140,N36141,N36142,N36143,N36144,N36145,N36146,N36147,N36148,
N36149,N36150,N36151,N36152,N36153,N36154,N36155,N36156,N36157,N36158,
N36159,N36160,N36161,N36162,N36163,N36164,N36165,N36166,N36167,N36168,
N36169,N36170,N36171,N36172,N36173,N36174,N36175,N36176,N36177,N36178,
N36179,N36180,N36181,N36182,N36183,N36184,N36185,N36186,N36187,N36188,
N36189,N36190,N36191,N36192,N36193,N36194,N36195,N36196,N36197,N36198,
N36199,N36200,N36201,N36202,N36203,N36204,N36205,N36206,N36207,N36208,
N36209,N36210,N36211,N36212,N36213,N36214,N36215,N36216,N36217,N36218,
N36219,N36220,N36221,N36222,N36223,N36224,N36225,N36226,N36227,N36228,
N36229,N36230,N36231,N36232,N36233,N36234,N36235,N36236,N36237,N36238,
N36239,N36240,N36241,N36242,N36243,N36244,N36245,N36246,N36247,N36248,
N36249,N36250,N36251,N36252,N36253,N36254,N36255,N36256,N36257,N36258,
N36259,N36260,N36261,N36262,N36263,N36264,N36265,N36266,N36267,N36268,
N36269,N36270,N36271,N36272,N36273,N36274,N36275,N36276,N36277,N36278,
N36279,N36280,N36281,N36282,N36283,N36284,N36285,N36286,N36287,N36288,
N36289,N36290,N36291,N36292,N36293,N36294,N36295,N36296,N36297,N36298,
N36299,N36300,N36301,N36302,N36303,N36304,N36305,N36306,N36307,N36308,
N36309,N36310,N36311,N36312,N36313,N36314,N36315,N36316,N36317,N36318,
N36319,N36320,N36321,N36322,N36323,N36324,N36325,N36326,N36327,N36328,
N36329,N36330,N36331,N36332,N36333,N36334,N36335,N36336,N36337,N36338,
N36339,N36340,N36341,N36342,N36343,N36344,N36345,N36346,N36347,N36348,
N36349,N36350,N36351,N36352,N36353,N36354,N36355,N36356,N36357,N36358,
N36359,N36360,N36361,N36362,N36363,N36364,N36365,N36366,N36367,N36368,
N36369,N36370,N36371,N36372,N36373,N36374,N36375,N36376,N36377,N36378,
N36379,N36380,N36381,N36382,N36383,N36384,N36385,N36386,N36387,N36388,
N36389,N36390,N36391,N36392,N36393,N36394,N36395,N36396,N36397,N36398,
N36399,N36400,N36401,N36402,N36403,N36404,N36405,N36406,N36407,N36408,
N36409,N36410,N36411,N36412,N36413,N36414,N36415,N36416,N36417,N36418,
N36419,N36420,N36421,N36422,N36423,N36424,N36425,N36426,N36427,N36428,
N36429,N36430,N36431,N36432,N36433,N36434,N36435,N36436,N36437,N36438,
N36439,N36440,N36441,N36442,N36443,N36444,N36445,N36446,N36447,N36448,
N36449,N36450,N36451,N36452,N36453,N36454,N36455,N36456,N36457,N36458,
N36459,N36460,N36461,N36462,N36463,N36464,N36465,N36466,N36467,N36468,
N36469,N36470,N36471,N36472,N36473,N36474,N36475,N36476,N36477,N36478,
N36479,N36480,N36481,N36482,N36483,N36484,N36485,N36486,N36487,N36488,
N36489,N36490,N36491,N36492,N36493,N36494,N36495,N36496,N36497,N36498,
N36499,N36500,N36501,N36502,N36503,N36504,N36505,N36506,N36507,N36508,
N36509,N36510,N36511,N36512,N36513,N36514,N36515,N36516,N36517,N36518,
N36519,N36520,N36521,N36522,N36523,N36524,N36525,N36526,N36527,N36528,
N36529,N36530,N36531,N36532,N36533,N36534,N36535,N36536,N36537,N36538,
N36539,N36540,N36541,N36542,N36543,N36544,N36545,N36546,N36547,N36548,
N36549,N36550,N36551,N36552,N36553,N36554,N36555,N36556,N36557,N36558,
N36559,N36560,N36561,N36562,N36563,N36564,N36565,N36566,N36567,N36568,
N36569,N36570,N36571,N36572,N36573,N36574,N36575,N36576,N36577,N36578,
N36579,N36580,N36581,N36582,N36583,N36584,N36585,N36586,N36587,N36588,
N36589,N36590,N36591,N36592,N36593,N36594,N36595,N36596,N36597,N36598,
N36599,N36600,N36601,N36602,N36603,N36604,N36605,N36606,N36607,N36608,
N36609,N36610,N36611,N36612,N36613,N36614,N36615,N36616,N36617,N36618,
N36619,N36620,N36621,N36622,N36623,N36624,N36625,N36626,N36627,N36628,
N36629,N36630,N36631,N36632,N36633,N36634,N36635,N36636,N36637,N36638,
N36639,N36640,N36641,N36642,N36643,N36644,N36645,N36646,N36647,N36648,
N36649,N36650,N36651,N36652,N36653,N36654,N36655,N36656,N36657,N36658,
N36659,N36660,N36661,N36662,N36663,N36664,N36665,N36666,N36667,N36668,
N36669,N36670,N36671,N36672,N36673,N36674,N36675,N36676,N36677,N36678,
N36679,N36680,N36681,N36682,N36683,N36684,N36685,N36686,N36687,N36688,
N36689,N36690,N36691,N36692,N36693,N36694,N36695,N36696,N36697,N36698,
N36699,N36700,N36701,N36702,N36703,N36704,N36705,N36706,N36707,N36708,
N36709,N36710,N36711,N36712,N36713,N36714,N36715,N36716,N36717,N36718,
N36719,N36720,N36721,N36722,N36723,N36724,N36725,N36726,N36727,N36728,
N36729,N36730,N36731,N36732,N36733,N36734,N36735,N36736,N36737,N36738,
N36739,N36740,N36741,N36742,N36743,N36744,N36745,N36746,N36747,N36748,
N36749,N36750,N36751,N36752,N36753,N36754,N36755,N36756,N36757,N36758,
N36759,N36760,N36761,N36762,N36763,N36764,N36765,N36766,N36767,N36768,
N36769,N36770,N36771,N36772,N36773,N36774,N36775,N36776,N36777,N36778,
N36779,N36780,N36781,N36782,N36783,N36784,N36785,N36786,N36787,N36788,
N36789,N36790,N36791,N36792,N36793,N36794,N36795,N36796,N36797,N36798,
N36799,N36800,N36801,N36802,N36803,N36804,N36805,N36806,N36807,N36808,
N36809,N36810,N36811,N36812,N36813,N36814,N36815,N36816,N36817,N36818,
N36819,N36820,N36821,N36822,N36823,N36824,N36825,N36826,N36827,N36828,
N36829,N36830,N36831,N36832,N36833,N36834,N36835,N36836,N36837,N36838,
N36839,N36840,N36841,N36842,N36843,N36844,N36845,N36846,N36847,N36848,
N36849,N36850,N36851,N36852,N36853,N36854,N36855,N36856,N36857,N36858,
N36859,N36860,N36861,N36862,N36863,N36864,N36865,N36866,N36867,N36868,
N36869,N36870,N36871,N36872,N36873,N36874,N36875,N36876,N36877,N36878,
N36879,N36880,N36881,N36882,N36883,N36884,N36885,N36886,N36887,N36888,
N36889,N36890,N36891,N36892,N36893,N36894,N36895,N36896,N36897,N36898,
N36899,N36900,N36901,N36902,N36903,N36904,N36905,N36906,N36907,N36908,
N36909,N36910,N36911,N36912,N36913,N36914,N36915,N36916,N36917,N36918,
N36919,N36920,N36921,N36922,N36923,N36924,N36925,N36926,N36927,N36928,
N36929,N36930,N36931,N36932,N36933,N36934,N36935,N36936,N36937,N36938,
N36939,N36940,N36941,N36942,N36943,N36944,N36945,N36946,N36947,N36948,
N36949,N36950,N36951,N36952,N36953,N36954,N36955,N36956,N36957,N36958,
N36959,N36960,N36961,N36962,N36963,N36964,N36965,N36966,N36967,N36968,
N36969,N36970,N36971,N36972,N36973,N36974,N36975,N36976,N36977,N36978,
N36979,N36980,N36981,N36982,N36983,N36984,N36985,N36986,N36987,N36988,
N36989,N36990,N36991,N36992,N36993,N36994,N36995,N36996,N36997,N36998,
N36999,N37000,N37001,N37002,N37003,N37004,N37005,N37006,N37007,N37008,
N37009,N37010,N37011,N37012,N37013,N37014,N37015,N37016,N37017,N37018,
N37019,N37020,N37021,N37022,N37023,N37024,N37025,N37026,N37027,N37028,
N37029,N37030,N37031,N37032,N37033,N37034,N37035,N37036,N37037,N37038,
N37039,N37040,N37041,N37042,N37043,N37044,N37045,N37046,N37047,N37048,
N37049,N37050,N37051,N37052,N37053,N37054,N37055,N37056,N37057,N37058,
N37059,N37060,N37061,N37062,N37063,N37064,N37065,N37066,N37067,N37068,
N37069,N37070,N37071,N37072,N37073,N37074,N37075,N37076,N37077,N37078,
N37079,N37080,N37081,N37082,N37083,N37084,N37085,N37086,N37087,N37088,
N37089,N37090,N37091,N37092,N37093,N37094,N37095,N37096,N37097,N37098,
N37099,N37100,N37101,N37102,N37103,N37104,N37105,N37106,N37107,N37108,
N37109,N37110,N37111,N37112,N37113,N37114,N37115,N37116,N37117,N37118,
N37119,N37120,N37121,N37122,N37123,N37124,N37125,N37126,N37127,N37128,
N37129,N37130,N37131,N37132,N37133,N37134,N37135,N37136,N37137,N37138,
N37139,N37140,N37141,N37142,N37143,N37144,N37145,clk,rst;

reg R0,R1,R2,R3,R4,R5,R6,R7,O0,O1,O2,O3,O4,O5;

always@(posedge clk or negedge rst)
 if(!rst)
   R0 <= N0;
   else
   R0= 1'b0;

always@(posedge clk or negedge rst)
 if(!rst)
   R1 <= N5661;
   else
   R1= 1'b0;

always@(posedge clk or negedge rst)
 if(!rst)
   R2 <= N8425;
   else
   R2= 1'b0;

always@(posedge clk or negedge rst)
 if(!rst)
   R3 <= N14726;
   else
   R3= 1'b0;

always@(posedge clk or negedge rst)
 if(!rst)
   R4 <= N20402;
   else
   R4= 1'b0;

always@(posedge clk or negedge rst)
 if(!rst)
   R5 <= N23823;
   else
   R5= 1'b0;

always@(posedge clk or negedge rst)
 if(!rst)
   R6 <= N29051;
   else
   R6= 1'b0;

always@(posedge clk or negedge rst)
 if(!rst)
   R7 <= N31564;
   else
   R7= 1'b0;

always@(posedge clk or negedge rst)
  if(!rst)
   O0 <= N34824;
  else
       O0=1'b0;
always@(posedge clk or negedge rst)
  if(!rst)
   O1 <= N35375;
  else
       O1=1'b0;
always@(posedge clk or negedge rst)
  if(!rst)
   O2 <= N35759;
  else
       O2=1'b0;
always@(posedge clk or negedge rst)
  if(!rst)
   O3 <= N35922;
  else
       O3=1'b0;
always@(posedge clk or negedge rst)
  if(!rst)
   O4 <= N36387;
  else
       O4=1'b0;
always@(posedge clk or negedge rst)
  if(!rst)
   O5 <= N36646;
  else
       O5=1'b0;

and and0(N411,N412,N413);
and and9(N428,N429,N430);
and and18(N445,N446,N447);
and and27(N462,N463,N464);
and and36(N479,N480,N481);
and and45(N496,N497,N498);
and and54(N513,N514,N515);
and and63(N530,N531,N532);
and and72(N547,N548,N549);
and and81(N564,N565,N566);
and and90(N581,N582,N583);
and and99(N598,N599,N600);
and and108(N615,N616,N617);
and and117(N631,N632,N633);
and and126(N647,N648,N649);
and and135(N663,N664,N665);
and and144(N679,N680,N681);
and and153(N695,N696,N697);
and and162(N711,N712,N713);
and and171(N727,N728,N729);
and and180(N743,N744,N745);
and and189(N759,N760,N761);
and and198(N775,N776,N777);
and and207(N791,N792,N793);
and and216(N807,N808,N809);
and and225(N822,N823,N824);
and and234(N837,N838,N839);
and and243(N852,N853,N854);
and and252(N867,N868,N869);
and and261(N882,N883,N884);
and and270(N897,N898,N899);
and and279(N912,N913,N914);
and and288(N927,N928,N929);
and and297(N942,N943,N944);
and and306(N957,N958,N959);
and and315(N972,N973,N974);
and and324(N987,N988,N989);
and and333(N1002,N1003,N1004);
and and342(N1017,N1018,N1019);
and and351(N1032,N1033,N1034);
and and360(N1047,N1048,N1049);
and and369(N1062,N1063,N1064);
and and378(N1077,N1078,N1079);
and and387(N1092,N1093,N1094);
and and396(N1107,N1108,N1109);
and and405(N1122,N1123,N1124);
and and414(N1137,N1138,N1139);
and and423(N1152,N1153,N1154);
and and432(N1167,N1168,N1169);
and and441(N1182,N1183,N1184);
and and450(N1197,N1198,N1199);
and and459(N1212,N1213,N1214);
and and468(N1227,N1228,N1229);
and and477(N1242,N1243,N1244);
and and486(N1257,N1258,N1259);
and and495(N1272,N1273,N1274);
and and504(N1287,N1288,N1289);
and and513(N1302,N1303,N1304);
and and522(N1317,N1318,N1319);
and and531(N1332,N1333,N1334);
and and540(N1347,N1348,N1349);
and and549(N1361,N1362,N1363);
and and558(N1375,N1376,N1377);
and and567(N1389,N1390,N1391);
and and576(N1403,N1404,N1405);
and and585(N1417,N1418,N1419);
and and594(N1431,N1432,N1433);
and and603(N1445,N1446,N1447);
and and612(N1459,N1460,N1461);
and and621(N1473,N1474,N1475);
and and630(N1487,N1488,N1489);
and and639(N1501,N1502,N1503);
and and648(N1515,N1516,N1517);
and and657(N1529,N1530,N1531);
and and666(N1543,N1544,N1545);
and and675(N1557,N1558,N1559);
and and684(N1571,N1572,N1573);
and and693(N1585,N1586,N1587);
and and702(N1599,N1600,N1601);
and and711(N1613,N1614,N1615);
and and720(N1627,N1628,N1629);
and and729(N1641,N1642,N1643);
and and738(N1655,N1656,N1657);
and and747(N1669,N1670,N1671);
and and756(N1683,N1684,N1685);
and and765(N1697,N1698,N1699);
and and774(N1711,N1712,N1713);
and and783(N1725,N1726,N1727);
and and792(N1738,N1739,N1740);
and and801(N1751,N1752,N1753);
and and810(N1764,N1765,N1766);
and and819(N1777,N1778,N1779);
and and828(N1790,N1791,N1792);
and and837(N1803,N1804,N1805);
and and846(N1816,N1817,N1818);
and and855(N1829,N1830,N1831);
and and864(N1842,N1843,N1844);
and and873(N1855,N1856,N1857);
and and882(N1868,N1869,N1870);
and and891(N1881,N1882,N1883);
and and900(N1894,N1895,N1896);
and and909(N1907,N1908,N1909);
and and918(N1920,N1921,N1922);
and and927(N1933,N1934,N1935);
and and936(N1946,N1947,N1948);
and and945(N1959,N1960,N1961);
and and954(N1972,N1973,N1974);
and and963(N1985,N1986,N1987);
and and972(N1998,N1999,N2000);
and and981(N2011,N2012,N2013);
and and990(N2024,N2025,N2026);
and and999(N2037,N2038,N2039);
and and1008(N2050,N2051,N2052);
and and1017(N2063,N2064,N2065);
and and1026(N2076,N2077,N2078);
and and1035(N2089,N2090,N2091);
and and1044(N2102,N2103,N2104);
and and1053(N2115,N2116,N2117);
and and1062(N2128,N2129,N2130);
and and1071(N2141,N2142,N2143);
and and1080(N2154,N2155,N2156);
and and1089(N2167,N2168,N2169);
and and1098(N2180,N2181,N2182);
and and1107(N2193,N2194,N2195);
and and1116(N2206,N2207,N2208);
and and1125(N2219,N2220,N2221);
and and1134(N2232,N2233,N2234);
and and1143(N2245,N2246,N2247);
and and1152(N2258,N2259,N2260);
and and1161(N2271,N2272,N2273);
and and1170(N2284,N2285,N2286);
and and1179(N2297,N2298,N2299);
and and1188(N2310,N2311,N2312);
and and1197(N2323,N2324,N2325);
and and1206(N2336,N2337,N2338);
and and1215(N2348,N2349,N2350);
and and1224(N2360,N2361,N2362);
and and1233(N2372,N2373,N2374);
and and1242(N2384,N2385,N2386);
and and1251(N2396,N2397,N2398);
and and1260(N2408,N2409,N2410);
and and1269(N2420,N2421,N2422);
and and1278(N2432,N2433,N2434);
and and1287(N2444,N2445,N2446);
and and1296(N2456,N2457,N2458);
and and1305(N2468,N2469,N2470);
and and1314(N2480,N2481,N2482);
and and1323(N2492,N2493,N2494);
and and1332(N2504,N2505,N2506);
and and1341(N2516,N2517,N2518);
and and1350(N2528,N2529,N2530);
and and1359(N2540,N2541,N2542);
and and1368(N2552,N2553,N2554);
and and1377(N2564,N2565,N2566);
and and1386(N2575,N2576,N2577);
and and1395(N2586,N2587,N2588);
and and1404(N2597,N2598,N2599);
and and1413(N2608,N2609,N2610);
and and1422(N2619,N2620,N2621);
and and1431(N2630,N2631,N2632);
and and1440(N2641,N2642,N2643);
and and1449(N2652,N2653,N2654);
and and1458(N2663,N2664,N2665);
and and1467(N2674,N2675,N2676);
and and1476(N2685,N2686,N2687);
and and1485(N2696,N2697,N2698);
and and1494(N2707,N2708,N2709);
and and1503(N2718,N2719,N2720);
and and1512(N2729,N2730,N2731);
and and1521(N2740,N2741,N2742);
and and1530(N2751,N2752,N2753);
and and1539(N2762,N2763,N2764);
and and1548(N2773,N2774,N2775);
and and1557(N2784,N2785,N2786);
and and1566(N2793,N2794,N2795);
and and1575(N2802,N2803,N2804);
and and1583(N2818,N2819,N2820);
and and1591(N2834,N2835,N2836);
and and1599(N2850,N2851,N2852);
and and1607(N2866,N2867,N2868);
and and1615(N2881,N2882,N2883);
and and1623(N2896,N2897,N2898);
and and1631(N2911,N2912,N2913);
and and1639(N2926,N2927,N2928);
and and1647(N2941,N2942,N2943);
and and1655(N2956,N2957,N2958);
and and1663(N2971,N2972,N2973);
and and1671(N2985,N2986,N2987);
and and1679(N2999,N3000,N3001);
and and1687(N3013,N3014,N3015);
and and1695(N3027,N3028,N3029);
and and1703(N3041,N3042,N3043);
and and1711(N3055,N3056,N3057);
and and1719(N3069,N3070,N3071);
and and1727(N3083,N3084,N3085);
and and1735(N3097,N3098,N3099);
and and1743(N3111,N3112,N3113);
and and1751(N3125,N3126,N3127);
and and1759(N3139,N3140,N3141);
and and1767(N3153,N3154,N3155);
and and1775(N3167,N3168,N3169);
and and1783(N3181,N3182,N3183);
and and1791(N3195,N3196,N3197);
and and1799(N3209,N3210,N3211);
and and1807(N3223,N3224,N3225);
and and1815(N3237,N3238,N3239);
and and1823(N3251,N3252,N3253);
and and1831(N3265,N3266,N3267);
and and1839(N3279,N3280,N3281);
and and1847(N3293,N3294,N3295);
and and1855(N3307,N3308,N3309);
and and1863(N3321,N3322,N3323);
and and1871(N3335,N3336,N3337);
and and1879(N3349,N3350,N3351);
and and1887(N3363,N3364,N3365);
and and1895(N3377,N3378,N3379);
and and1903(N3391,N3392,N3393);
and and1911(N3405,N3406,N3407);
and and1919(N3419,N3420,N3421);
and and1927(N3433,N3434,N3435);
and and1935(N3447,N3448,N3449);
and and1943(N3461,N3462,N3463);
and and1951(N3475,N3476,N3477);
and and1959(N3488,N3489,N3490);
and and1967(N3501,N3502,N3503);
and and1975(N3514,N3515,N3516);
and and1983(N3527,N3528,N3529);
and and1991(N3540,N3541,N3542);
and and1999(N3553,N3554,N3555);
and and2007(N3566,N3567,N3568);
and and2015(N3579,N3580,N3581);
and and2023(N3592,N3593,N3594);
and and2031(N3605,N3606,N3607);
and and2039(N3618,N3619,N3620);
and and2047(N3631,N3632,N3633);
and and2055(N3644,N3645,N3646);
and and2063(N3657,N3658,N3659);
and and2071(N3670,N3671,N3672);
and and2079(N3683,N3684,N3685);
and and2087(N3696,N3697,N3698);
and and2095(N3709,N3710,N3711);
and and2103(N3722,N3723,N3724);
and and2111(N3735,N3736,N3737);
and and2119(N3748,N3749,N3750);
and and2127(N3761,N3762,N3763);
and and2135(N3774,N3775,N3776);
and and2143(N3787,N3788,N3789);
and and2151(N3800,N3801,N3802);
and and2159(N3813,N3814,N3815);
and and2167(N3826,N3827,N3828);
and and2175(N3839,N3840,N3841);
and and2183(N3852,N3853,N3854);
and and2191(N3865,N3866,N3867);
and and2199(N3878,N3879,N3880);
and and2207(N3891,N3892,N3893);
and and2215(N3904,N3905,N3906);
and and2223(N3917,N3918,N3919);
and and2231(N3930,N3931,N3932);
and and2239(N3943,N3944,N3945);
and and2247(N3956,N3957,N3958);
and and2255(N3969,N3970,N3971);
and and2263(N3981,N3982,N3983);
and and2271(N3993,N3994,N3995);
and and2279(N4005,N4006,N4007);
and and2287(N4017,N4018,N4019);
and and2295(N4029,N4030,N4031);
and and2303(N4041,N4042,N4043);
and and2311(N4053,N4054,N4055);
and and2319(N4065,N4066,N4067);
and and2327(N4077,N4078,N4079);
and and2335(N4089,N4090,N4091);
and and2343(N4101,N4102,N4103);
and and2351(N4113,N4114,N4115);
and and2359(N4125,N4126,N4127);
and and2367(N4137,N4138,N4139);
and and2375(N4149,N4150,N4151);
and and2383(N4161,N4162,N4163);
and and2391(N4173,N4174,N4175);
and and2399(N4185,N4186,N4187);
and and2407(N4197,N4198,N4199);
and and2415(N4209,N4210,N4211);
and and2423(N4221,N4222,N4223);
and and2431(N4233,N4234,N4235);
and and2439(N4245,N4246,N4247);
and and2447(N4257,N4258,N4259);
and and2455(N4269,N4270,N4271);
and and2463(N4281,N4282,N4283);
and and2471(N4293,N4294,N4295);
and and2479(N4305,N4306,N4307);
and and2487(N4317,N4318,N4319);
and and2495(N4329,N4330,N4331);
and and2503(N4341,N4342,N4343);
and and2511(N4353,N4354,N4355);
and and2519(N4365,N4366,N4367);
and and2527(N4377,N4378,N4379);
and and2535(N4389,N4390,N4391);
and and2543(N4401,N4402,N4403);
and and2551(N4413,N4414,N4415);
and and2559(N4425,N4426,N4427);
and and2567(N4437,N4438,N4439);
and and2575(N4449,N4450,N4451);
and and2583(N4461,N4462,N4463);
and and2591(N4473,N4474,N4475);
and and2599(N4485,N4486,N4487);
and and2607(N4497,N4498,N4499);
and and2615(N4509,N4510,N4511);
and and2623(N4521,N4522,N4523);
and and2631(N4533,N4534,N4535);
and and2639(N4545,N4546,N4547);
and and2647(N4557,N4558,N4559);
and and2655(N4569,N4570,N4571);
and and2663(N4581,N4582,N4583);
and and2671(N4593,N4594,N4595);
and and2679(N4604,N4605,N4606);
and and2687(N4615,N4616,N4617);
and and2695(N4626,N4627,N4628);
and and2703(N4637,N4638,N4639);
and and2711(N4648,N4649,N4650);
and and2719(N4659,N4660,N4661);
and and2727(N4670,N4671,N4672);
and and2735(N4681,N4682,N4683);
and and2743(N4692,N4693,N4694);
and and2751(N4703,N4704,N4705);
and and2759(N4714,N4715,N4716);
and and2767(N4725,N4726,N4727);
and and2775(N4736,N4737,N4738);
and and2783(N4747,N4748,N4749);
and and2791(N4758,N4759,N4760);
and and2799(N4769,N4770,N4771);
and and2807(N4780,N4781,N4782);
and and2815(N4791,N4792,N4793);
and and2823(N4802,N4803,N4804);
and and2831(N4813,N4814,N4815);
and and2839(N4824,N4825,N4826);
and and2847(N4835,N4836,N4837);
and and2855(N4846,N4847,N4848);
and and2863(N4857,N4858,N4859);
and and2871(N4868,N4869,N4870);
and and2879(N4879,N4880,N4881);
and and2887(N4890,N4891,N4892);
and and2895(N4900,N4901,N4902);
and and2903(N4910,N4911,N4912);
and and2911(N4920,N4921,N4922);
and and2919(N4930,N4931,N4932);
and and2927(N4940,N4941,N4942);
and and2935(N4950,N4951,N4952);
and and2943(N4960,N4961,N4962);
and and2951(N4970,N4971,N4972);
and and2959(N4980,N4981,N4982);
and and2967(N4990,N4991,N4992);
and and2975(N5000,N5001,N5002);
and and2983(N5010,N5011,N5012);
and and2991(N5020,N5021,N5022);
and and2999(N5030,N5031,N5032);
and and3007(N5040,N5041,N5042);
and and3015(N5050,N5051,N5052);
and and3023(N5060,N5061,N5062);
and and3031(N5070,N5071,N5072);
and and3039(N5079,N5080,N5081);
and and3047(N5088,N5089,N5090);
and and3055(N5097,N5098,N5099);
and and3063(N5106,N5107,N5108);
and and3071(N5115,N5116,N5117);
and and3079(N5124,N5125,N5126);
and and3086(N5138,N5139,N5140);
and and3093(N5152,N5153,N5154);
and and3100(N5166,N5167,N5168);
and and3107(N5179,N5180,N5181);
and and3114(N5192,N5193,N5194);
and and3121(N5205,N5206,N5207);
and and3128(N5218,N5219,N5220);
and and3135(N5231,N5232,N5233);
and and3142(N5243,N5244,N5245);
and and3149(N5255,N5256,N5257);
and and3156(N5267,N5268,N5269);
and and3163(N5279,N5280,N5281);
and and3170(N5291,N5292,N5293);
and and3177(N5303,N5304,N5305);
and and3184(N5315,N5316,N5317);
and and3191(N5327,N5328,N5329);
and and3198(N5338,N5339,N5340);
and and3205(N5349,N5350,N5351);
and and3212(N5360,N5361,N5362);
and and3219(N5371,N5372,N5373);
and and3226(N5382,N5383,N5384);
and and3233(N5393,N5394,N5395);
and and3240(N5404,N5405,N5406);
and and3247(N5415,N5416,N5417);
and and3254(N5426,N5427,N5428);
and and3261(N5437,N5438,N5439);
and and3268(N5448,N5449,N5450);
and and3275(N5459,N5460,N5461);
and and3282(N5470,N5471,N5472);
and and3289(N5481,N5482,N5483);
and and3296(N5491,N5492,N5493);
and and3303(N5501,N5502,N5503);
and and3310(N5511,N5512,N5513);
and and3317(N5521,N5522,N5523);
and and3324(N5531,N5532,N5533);
and and3331(N5541,N5542,N5543);
and and3338(N5551,N5552,N5553);
and and3345(N5561,N5562,N5563);
and and3352(N5571,N5572,N5573);
and and3359(N5581,N5582,N5583);
and and3366(N5591,N5592,N5593);
and and3373(N5601,N5602,N5603);
and and3380(N5610,N5611,N5612);
and and3387(N5619,N5620,N5621);
and and3394(N5628,N5629,N5630);
and and3401(N5637,N5638,N5639);
and and3408(N5646,N5647,N5648);
and and3415(N5654,N5655,N5656);
and and1(N412,N414,N415);
and and2(N413,N416,N417);
and and10(N429,N431,N432);
and and11(N430,N433,N434);
and and19(N446,N448,N449);
and and20(N447,N450,N451);
and and28(N463,N465,N466);
and and29(N464,N467,N468);
and and37(N480,N482,N483);
and and38(N481,N484,N485);
and and46(N497,N499,N500);
and and47(N498,N501,N502);
and and55(N514,N516,N517);
and and56(N515,N518,N519);
and and64(N531,N533,N534);
and and65(N532,N535,N536);
and and73(N548,N550,N551);
and and74(N549,N552,N553);
and and82(N565,N567,N568);
and and83(N566,N569,N570);
and and91(N582,N584,N585);
and and92(N583,N586,N587);
and and100(N599,N601,N602);
and and101(N600,N603,N604);
and and109(N616,N618,N619);
and and110(N617,N620,N621);
and and118(N632,N634,N635);
and and119(N633,N636,N637);
and and127(N648,N650,N651);
and and128(N649,N652,N653);
and and136(N664,N666,N667);
and and137(N665,N668,N669);
and and145(N680,N682,N683);
and and146(N681,N684,N685);
and and154(N696,N698,N699);
and and155(N697,N700,N701);
and and163(N712,N714,N715);
and and164(N713,N716,N717);
and and172(N728,N730,N731);
and and173(N729,N732,N733);
and and181(N744,N746,N747);
and and182(N745,N748,N749);
and and190(N760,N762,N763);
and and191(N761,N764,N765);
and and199(N776,N778,N779);
and and200(N777,N780,N781);
and and208(N792,N794,N795);
and and209(N793,N796,N797);
and and217(N808,N810,N811);
and and218(N809,N812,N813);
and and226(N823,N825,N826);
and and227(N824,N827,N828);
and and235(N838,N840,N841);
and and236(N839,N842,N843);
and and244(N853,N855,N856);
and and245(N854,N857,N858);
and and253(N868,N870,N871);
and and254(N869,N872,N873);
and and262(N883,N885,N886);
and and263(N884,N887,N888);
and and271(N898,N900,N901);
and and272(N899,N902,N903);
and and280(N913,N915,N916);
and and281(N914,N917,N918);
and and289(N928,N930,N931);
and and290(N929,N932,N933);
and and298(N943,N945,N946);
and and299(N944,N947,N948);
and and307(N958,N960,N961);
and and308(N959,N962,N963);
and and316(N973,N975,N976);
and and317(N974,N977,N978);
and and325(N988,N990,N991);
and and326(N989,N992,N993);
and and334(N1003,N1005,N1006);
and and335(N1004,N1007,N1008);
and and343(N1018,N1020,N1021);
and and344(N1019,N1022,N1023);
and and352(N1033,N1035,N1036);
and and353(N1034,N1037,N1038);
and and361(N1048,N1050,N1051);
and and362(N1049,N1052,N1053);
and and370(N1063,N1065,N1066);
and and371(N1064,N1067,N1068);
and and379(N1078,N1080,N1081);
and and380(N1079,N1082,N1083);
and and388(N1093,N1095,N1096);
and and389(N1094,N1097,N1098);
and and397(N1108,N1110,N1111);
and and398(N1109,N1112,N1113);
and and406(N1123,N1125,N1126);
and and407(N1124,N1127,N1128);
and and415(N1138,N1140,N1141);
and and416(N1139,N1142,N1143);
and and424(N1153,N1155,N1156);
and and425(N1154,N1157,N1158);
and and433(N1168,N1170,N1171);
and and434(N1169,N1172,N1173);
and and442(N1183,N1185,N1186);
and and443(N1184,N1187,N1188);
and and451(N1198,N1200,N1201);
and and452(N1199,N1202,N1203);
and and460(N1213,N1215,N1216);
and and461(N1214,N1217,N1218);
and and469(N1228,N1230,N1231);
and and470(N1229,N1232,N1233);
and and478(N1243,N1245,N1246);
and and479(N1244,N1247,N1248);
and and487(N1258,N1260,N1261);
and and488(N1259,N1262,N1263);
and and496(N1273,N1275,N1276);
and and497(N1274,N1277,N1278);
and and505(N1288,N1290,N1291);
and and506(N1289,N1292,N1293);
and and514(N1303,N1305,N1306);
and and515(N1304,N1307,N1308);
and and523(N1318,N1320,N1321);
and and524(N1319,N1322,N1323);
and and532(N1333,N1335,N1336);
and and533(N1334,N1337,N1338);
and and541(N1348,N1350,N1351);
and and542(N1349,N1352,N1353);
and and550(N1362,N1364,N1365);
and and551(N1363,N1366,N1367);
and and559(N1376,N1378,N1379);
and and560(N1377,N1380,N1381);
and and568(N1390,N1392,N1393);
and and569(N1391,N1394,N1395);
and and577(N1404,N1406,N1407);
and and578(N1405,N1408,N1409);
and and586(N1418,N1420,N1421);
and and587(N1419,N1422,N1423);
and and595(N1432,N1434,N1435);
and and596(N1433,N1436,N1437);
and and604(N1446,N1448,N1449);
and and605(N1447,N1450,N1451);
and and613(N1460,N1462,N1463);
and and614(N1461,N1464,N1465);
and and622(N1474,N1476,N1477);
and and623(N1475,N1478,N1479);
and and631(N1488,N1490,N1491);
and and632(N1489,N1492,N1493);
and and640(N1502,N1504,N1505);
and and641(N1503,N1506,N1507);
and and649(N1516,N1518,N1519);
and and650(N1517,N1520,N1521);
and and658(N1530,N1532,N1533);
and and659(N1531,N1534,N1535);
and and667(N1544,N1546,N1547);
and and668(N1545,N1548,N1549);
and and676(N1558,N1560,N1561);
and and677(N1559,N1562,N1563);
and and685(N1572,N1574,N1575);
and and686(N1573,N1576,N1577);
and and694(N1586,N1588,N1589);
and and695(N1587,N1590,N1591);
and and703(N1600,N1602,N1603);
and and704(N1601,N1604,N1605);
and and712(N1614,N1616,N1617);
and and713(N1615,N1618,N1619);
and and721(N1628,N1630,N1631);
and and722(N1629,N1632,N1633);
and and730(N1642,N1644,N1645);
and and731(N1643,N1646,N1647);
and and739(N1656,N1658,N1659);
and and740(N1657,N1660,N1661);
and and748(N1670,N1672,N1673);
and and749(N1671,N1674,N1675);
and and757(N1684,N1686,N1687);
and and758(N1685,N1688,N1689);
and and766(N1698,N1700,N1701);
and and767(N1699,N1702,N1703);
and and775(N1712,N1714,N1715);
and and776(N1713,N1716,N1717);
and and784(N1726,N1728,N1729);
and and785(N1727,N1730,N1731);
and and793(N1739,N1741,N1742);
and and794(N1740,N1743,N1744);
and and802(N1752,N1754,N1755);
and and803(N1753,N1756,N1757);
and and811(N1765,N1767,N1768);
and and812(N1766,N1769,N1770);
and and820(N1778,N1780,N1781);
and and821(N1779,N1782,N1783);
and and829(N1791,N1793,N1794);
and and830(N1792,N1795,N1796);
and and838(N1804,N1806,N1807);
and and839(N1805,N1808,N1809);
and and847(N1817,N1819,N1820);
and and848(N1818,N1821,N1822);
and and856(N1830,N1832,N1833);
and and857(N1831,N1834,N1835);
and and865(N1843,N1845,N1846);
and and866(N1844,N1847,N1848);
and and874(N1856,N1858,N1859);
and and875(N1857,N1860,N1861);
and and883(N1869,N1871,N1872);
and and884(N1870,N1873,N1874);
and and892(N1882,N1884,N1885);
and and893(N1883,N1886,N1887);
and and901(N1895,N1897,N1898);
and and902(N1896,N1899,N1900);
and and910(N1908,N1910,N1911);
and and911(N1909,N1912,N1913);
and and919(N1921,N1923,N1924);
and and920(N1922,N1925,N1926);
and and928(N1934,N1936,N1937);
and and929(N1935,N1938,N1939);
and and937(N1947,N1949,N1950);
and and938(N1948,N1951,N1952);
and and946(N1960,N1962,N1963);
and and947(N1961,N1964,N1965);
and and955(N1973,N1975,N1976);
and and956(N1974,N1977,N1978);
and and964(N1986,N1988,N1989);
and and965(N1987,N1990,N1991);
and and973(N1999,N2001,N2002);
and and974(N2000,N2003,N2004);
and and982(N2012,N2014,N2015);
and and983(N2013,N2016,N2017);
and and991(N2025,N2027,N2028);
and and992(N2026,N2029,N2030);
and and1000(N2038,N2040,N2041);
and and1001(N2039,N2042,N2043);
and and1009(N2051,N2053,N2054);
and and1010(N2052,N2055,N2056);
and and1018(N2064,N2066,N2067);
and and1019(N2065,N2068,N2069);
and and1027(N2077,N2079,N2080);
and and1028(N2078,N2081,N2082);
and and1036(N2090,N2092,N2093);
and and1037(N2091,N2094,N2095);
and and1045(N2103,N2105,N2106);
and and1046(N2104,N2107,N2108);
and and1054(N2116,N2118,N2119);
and and1055(N2117,N2120,N2121);
and and1063(N2129,N2131,N2132);
and and1064(N2130,N2133,N2134);
and and1072(N2142,N2144,N2145);
and and1073(N2143,N2146,N2147);
and and1081(N2155,N2157,N2158);
and and1082(N2156,N2159,N2160);
and and1090(N2168,N2170,N2171);
and and1091(N2169,N2172,N2173);
and and1099(N2181,N2183,N2184);
and and1100(N2182,N2185,N2186);
and and1108(N2194,N2196,N2197);
and and1109(N2195,N2198,N2199);
and and1117(N2207,N2209,N2210);
and and1118(N2208,N2211,N2212);
and and1126(N2220,N2222,N2223);
and and1127(N2221,N2224,N2225);
and and1135(N2233,N2235,N2236);
and and1136(N2234,N2237,N2238);
and and1144(N2246,N2248,N2249);
and and1145(N2247,N2250,N2251);
and and1153(N2259,N2261,N2262);
and and1154(N2260,N2263,N2264);
and and1162(N2272,N2274,N2275);
and and1163(N2273,N2276,N2277);
and and1171(N2285,N2287,N2288);
and and1172(N2286,N2289,N2290);
and and1180(N2298,N2300,N2301);
and and1181(N2299,N2302,N2303);
and and1189(N2311,N2313,N2314);
and and1190(N2312,N2315,N2316);
and and1198(N2324,N2326,N2327);
and and1199(N2325,N2328,N2329);
and and1207(N2337,N2339,N2340);
and and1208(N2338,N2341,N2342);
and and1216(N2349,N2351,N2352);
and and1217(N2350,N2353,N2354);
and and1225(N2361,N2363,N2364);
and and1226(N2362,N2365,N2366);
and and1234(N2373,N2375,N2376);
and and1235(N2374,N2377,N2378);
and and1243(N2385,N2387,N2388);
and and1244(N2386,N2389,N2390);
and and1252(N2397,N2399,N2400);
and and1253(N2398,N2401,N2402);
and and1261(N2409,N2411,N2412);
and and1262(N2410,N2413,N2414);
and and1270(N2421,N2423,N2424);
and and1271(N2422,N2425,N2426);
and and1279(N2433,N2435,N2436);
and and1280(N2434,N2437,N2438);
and and1288(N2445,N2447,N2448);
and and1289(N2446,N2449,N2450);
and and1297(N2457,N2459,N2460);
and and1298(N2458,N2461,N2462);
and and1306(N2469,N2471,N2472);
and and1307(N2470,N2473,N2474);
and and1315(N2481,N2483,N2484);
and and1316(N2482,N2485,N2486);
and and1324(N2493,N2495,N2496);
and and1325(N2494,N2497,N2498);
and and1333(N2505,N2507,N2508);
and and1334(N2506,N2509,N2510);
and and1342(N2517,N2519,N2520);
and and1343(N2518,N2521,N2522);
and and1351(N2529,N2531,N2532);
and and1352(N2530,N2533,N2534);
and and1360(N2541,N2543,N2544);
and and1361(N2542,N2545,N2546);
and and1369(N2553,N2555,N2556);
and and1370(N2554,N2557,N2558);
and and1378(N2565,N2567,N2568);
and and1379(N2566,N2569,N2570);
and and1387(N2576,N2578,N2579);
and and1388(N2577,N2580,N2581);
and and1396(N2587,N2589,N2590);
and and1397(N2588,N2591,N2592);
and and1405(N2598,N2600,N2601);
and and1406(N2599,N2602,N2603);
and and1414(N2609,N2611,N2612);
and and1415(N2610,N2613,N2614);
and and1423(N2620,N2622,N2623);
and and1424(N2621,N2624,N2625);
and and1432(N2631,N2633,N2634);
and and1433(N2632,N2635,N2636);
and and1441(N2642,N2644,N2645);
and and1442(N2643,N2646,N2647);
and and1450(N2653,N2655,N2656);
and and1451(N2654,N2657,N2658);
and and1459(N2664,N2666,N2667);
and and1460(N2665,N2668,N2669);
and and1468(N2675,N2677,N2678);
and and1469(N2676,N2679,N2680);
and and1477(N2686,N2688,N2689);
and and1478(N2687,N2690,N2691);
and and1486(N2697,N2699,N2700);
and and1487(N2698,N2701,N2702);
and and1495(N2708,N2710,N2711);
and and1496(N2709,N2712,N2713);
and and1504(N2719,N2721,N2722);
and and1505(N2720,N2723,N2724);
and and1513(N2730,N2732,N2733);
and and1514(N2731,N2734,N2735);
and and1522(N2741,N2743,N2744);
and and1523(N2742,N2745,N2746);
and and1531(N2752,N2754,N2755);
and and1532(N2753,N2756,N2757);
and and1540(N2763,N2765,N2766);
and and1541(N2764,N2767,N2768);
and and1549(N2774,N2776,N2777);
and and1550(N2775,N2778,N2779);
and and1558(N2785,N2787,N2788);
and and1559(N2786,N2789,N2790);
and and1567(N2794,N2796,N2797);
and and1568(N2795,N2798,N2799);
and and1576(N2803,N2805,N2806);
and and1577(N2804,N2807,N2808);
and and1584(N2819,N2821,N2822);
and and1585(N2820,N2823,N2824);
and and1592(N2835,N2837,N2838);
and and1593(N2836,N2839,N2840);
and and1600(N2851,N2853,N2854);
and and1601(N2852,N2855,N2856);
and and1608(N2867,N2869,N2870);
and and1609(N2868,N2871,N2872);
and and1616(N2882,N2884,N2885);
and and1617(N2883,N2886,N2887);
and and1624(N2897,N2899,N2900);
and and1625(N2898,N2901,N2902);
and and1632(N2912,N2914,N2915);
and and1633(N2913,N2916,N2917);
and and1640(N2927,N2929,N2930);
and and1641(N2928,N2931,N2932);
and and1648(N2942,N2944,N2945);
and and1649(N2943,N2946,N2947);
and and1656(N2957,N2959,N2960);
and and1657(N2958,N2961,N2962);
and and1664(N2972,N2974,N2975);
and and1665(N2973,N2976,N2977);
and and1672(N2986,N2988,N2989);
and and1673(N2987,N2990,N2991);
and and1680(N3000,N3002,N3003);
and and1681(N3001,N3004,N3005);
and and1688(N3014,N3016,N3017);
and and1689(N3015,N3018,N3019);
and and1696(N3028,N3030,N3031);
and and1697(N3029,N3032,N3033);
and and1704(N3042,N3044,N3045);
and and1705(N3043,N3046,N3047);
and and1712(N3056,N3058,N3059);
and and1713(N3057,N3060,N3061);
and and1720(N3070,N3072,N3073);
and and1721(N3071,N3074,N3075);
and and1728(N3084,N3086,N3087);
and and1729(N3085,N3088,N3089);
and and1736(N3098,N3100,N3101);
and and1737(N3099,N3102,N3103);
and and1744(N3112,N3114,N3115);
and and1745(N3113,N3116,N3117);
and and1752(N3126,N3128,N3129);
and and1753(N3127,N3130,N3131);
and and1760(N3140,N3142,N3143);
and and1761(N3141,N3144,N3145);
and and1768(N3154,N3156,N3157);
and and1769(N3155,N3158,N3159);
and and1776(N3168,N3170,N3171);
and and1777(N3169,N3172,N3173);
and and1784(N3182,N3184,N3185);
and and1785(N3183,N3186,N3187);
and and1792(N3196,N3198,N3199);
and and1793(N3197,N3200,N3201);
and and1800(N3210,N3212,N3213);
and and1801(N3211,N3214,N3215);
and and1808(N3224,N3226,N3227);
and and1809(N3225,N3228,N3229);
and and1816(N3238,N3240,N3241);
and and1817(N3239,N3242,N3243);
and and1824(N3252,N3254,N3255);
and and1825(N3253,N3256,N3257);
and and1832(N3266,N3268,N3269);
and and1833(N3267,N3270,N3271);
and and1840(N3280,N3282,N3283);
and and1841(N3281,N3284,N3285);
and and1848(N3294,N3296,N3297);
and and1849(N3295,N3298,N3299);
and and1856(N3308,N3310,N3311);
and and1857(N3309,N3312,N3313);
and and1864(N3322,N3324,N3325);
and and1865(N3323,N3326,N3327);
and and1872(N3336,N3338,N3339);
and and1873(N3337,N3340,N3341);
and and1880(N3350,N3352,N3353);
and and1881(N3351,N3354,N3355);
and and1888(N3364,N3366,N3367);
and and1889(N3365,N3368,N3369);
and and1896(N3378,N3380,N3381);
and and1897(N3379,N3382,N3383);
and and1904(N3392,N3394,N3395);
and and1905(N3393,N3396,N3397);
and and1912(N3406,N3408,N3409);
and and1913(N3407,N3410,N3411);
and and1920(N3420,N3422,N3423);
and and1921(N3421,N3424,N3425);
and and1928(N3434,N3436,N3437);
and and1929(N3435,N3438,N3439);
and and1936(N3448,N3450,N3451);
and and1937(N3449,N3452,N3453);
and and1944(N3462,N3464,N3465);
and and1945(N3463,N3466,N3467);
and and1952(N3476,N3478,N3479);
and and1953(N3477,N3480,N3481);
and and1960(N3489,N3491,N3492);
and and1961(N3490,N3493,N3494);
and and1968(N3502,N3504,N3505);
and and1969(N3503,N3506,N3507);
and and1976(N3515,N3517,N3518);
and and1977(N3516,N3519,N3520);
and and1984(N3528,N3530,N3531);
and and1985(N3529,N3532,N3533);
and and1992(N3541,N3543,N3544);
and and1993(N3542,N3545,N3546);
and and2000(N3554,N3556,N3557);
and and2001(N3555,N3558,N3559);
and and2008(N3567,N3569,N3570);
and and2009(N3568,N3571,N3572);
and and2016(N3580,N3582,N3583);
and and2017(N3581,N3584,N3585);
and and2024(N3593,N3595,N3596);
and and2025(N3594,N3597,N3598);
and and2032(N3606,N3608,N3609);
and and2033(N3607,N3610,N3611);
and and2040(N3619,N3621,N3622);
and and2041(N3620,N3623,N3624);
and and2048(N3632,N3634,N3635);
and and2049(N3633,N3636,N3637);
and and2056(N3645,N3647,N3648);
and and2057(N3646,N3649,N3650);
and and2064(N3658,N3660,N3661);
and and2065(N3659,N3662,N3663);
and and2072(N3671,N3673,N3674);
and and2073(N3672,N3675,N3676);
and and2080(N3684,N3686,N3687);
and and2081(N3685,N3688,N3689);
and and2088(N3697,N3699,N3700);
and and2089(N3698,N3701,N3702);
and and2096(N3710,N3712,N3713);
and and2097(N3711,N3714,N3715);
and and2104(N3723,N3725,N3726);
and and2105(N3724,N3727,N3728);
and and2112(N3736,N3738,N3739);
and and2113(N3737,N3740,N3741);
and and2120(N3749,N3751,N3752);
and and2121(N3750,N3753,N3754);
and and2128(N3762,N3764,N3765);
and and2129(N3763,N3766,N3767);
and and2136(N3775,N3777,N3778);
and and2137(N3776,N3779,N3780);
and and2144(N3788,N3790,N3791);
and and2145(N3789,N3792,N3793);
and and2152(N3801,N3803,N3804);
and and2153(N3802,N3805,N3806);
and and2160(N3814,N3816,N3817);
and and2161(N3815,N3818,N3819);
and and2168(N3827,N3829,N3830);
and and2169(N3828,N3831,N3832);
and and2176(N3840,N3842,N3843);
and and2177(N3841,N3844,N3845);
and and2184(N3853,N3855,N3856);
and and2185(N3854,N3857,N3858);
and and2192(N3866,N3868,N3869);
and and2193(N3867,N3870,N3871);
and and2200(N3879,N3881,N3882);
and and2201(N3880,N3883,N3884);
and and2208(N3892,N3894,N3895);
and and2209(N3893,N3896,N3897);
and and2216(N3905,N3907,N3908);
and and2217(N3906,N3909,N3910);
and and2224(N3918,N3920,N3921);
and and2225(N3919,N3922,N3923);
and and2232(N3931,N3933,N3934);
and and2233(N3932,N3935,N3936);
and and2240(N3944,N3946,N3947);
and and2241(N3945,N3948,N3949);
and and2248(N3957,N3959,N3960);
and and2249(N3958,N3961,N3962);
and and2256(N3970,N3972,N3973);
and and2257(N3971,N3974,N3975);
and and2264(N3982,N3984,N3985);
and and2265(N3983,N3986,N3987);
and and2272(N3994,N3996,N3997);
and and2273(N3995,N3998,N3999);
and and2280(N4006,N4008,N4009);
and and2281(N4007,N4010,N4011);
and and2288(N4018,N4020,N4021);
and and2289(N4019,N4022,N4023);
and and2296(N4030,N4032,N4033);
and and2297(N4031,N4034,N4035);
and and2304(N4042,N4044,N4045);
and and2305(N4043,N4046,N4047);
and and2312(N4054,N4056,N4057);
and and2313(N4055,N4058,N4059);
and and2320(N4066,N4068,N4069);
and and2321(N4067,N4070,N4071);
and and2328(N4078,N4080,N4081);
and and2329(N4079,N4082,N4083);
and and2336(N4090,N4092,N4093);
and and2337(N4091,N4094,N4095);
and and2344(N4102,N4104,N4105);
and and2345(N4103,N4106,N4107);
and and2352(N4114,N4116,N4117);
and and2353(N4115,N4118,N4119);
and and2360(N4126,N4128,N4129);
and and2361(N4127,N4130,N4131);
and and2368(N4138,N4140,N4141);
and and2369(N4139,N4142,N4143);
and and2376(N4150,N4152,N4153);
and and2377(N4151,N4154,N4155);
and and2384(N4162,N4164,N4165);
and and2385(N4163,N4166,N4167);
and and2392(N4174,N4176,N4177);
and and2393(N4175,N4178,N4179);
and and2400(N4186,N4188,N4189);
and and2401(N4187,N4190,N4191);
and and2408(N4198,N4200,N4201);
and and2409(N4199,N4202,N4203);
and and2416(N4210,N4212,N4213);
and and2417(N4211,N4214,N4215);
and and2424(N4222,N4224,N4225);
and and2425(N4223,N4226,N4227);
and and2432(N4234,N4236,N4237);
and and2433(N4235,N4238,N4239);
and and2440(N4246,N4248,N4249);
and and2441(N4247,N4250,N4251);
and and2448(N4258,N4260,N4261);
and and2449(N4259,N4262,N4263);
and and2456(N4270,N4272,N4273);
and and2457(N4271,N4274,N4275);
and and2464(N4282,N4284,N4285);
and and2465(N4283,N4286,N4287);
and and2472(N4294,N4296,N4297);
and and2473(N4295,N4298,N4299);
and and2480(N4306,N4308,N4309);
and and2481(N4307,N4310,N4311);
and and2488(N4318,N4320,N4321);
and and2489(N4319,N4322,N4323);
and and2496(N4330,N4332,N4333);
and and2497(N4331,N4334,N4335);
and and2504(N4342,N4344,N4345);
and and2505(N4343,N4346,N4347);
and and2512(N4354,N4356,N4357);
and and2513(N4355,N4358,N4359);
and and2520(N4366,N4368,N4369);
and and2521(N4367,N4370,N4371);
and and2528(N4378,N4380,N4381);
and and2529(N4379,N4382,N4383);
and and2536(N4390,N4392,N4393);
and and2537(N4391,N4394,N4395);
and and2544(N4402,N4404,N4405);
and and2545(N4403,N4406,N4407);
and and2552(N4414,N4416,N4417);
and and2553(N4415,N4418,N4419);
and and2560(N4426,N4428,N4429);
and and2561(N4427,N4430,N4431);
and and2568(N4438,N4440,N4441);
and and2569(N4439,N4442,N4443);
and and2576(N4450,N4452,N4453);
and and2577(N4451,N4454,N4455);
and and2584(N4462,N4464,N4465);
and and2585(N4463,N4466,N4467);
and and2592(N4474,N4476,N4477);
and and2593(N4475,N4478,N4479);
and and2600(N4486,N4488,N4489);
and and2601(N4487,N4490,N4491);
and and2608(N4498,N4500,N4501);
and and2609(N4499,N4502,N4503);
and and2616(N4510,N4512,N4513);
and and2617(N4511,N4514,N4515);
and and2624(N4522,N4524,N4525);
and and2625(N4523,N4526,N4527);
and and2632(N4534,N4536,N4537);
and and2633(N4535,N4538,N4539);
and and2640(N4546,N4548,N4549);
and and2641(N4547,N4550,N4551);
and and2648(N4558,N4560,N4561);
and and2649(N4559,N4562,N4563);
and and2656(N4570,N4572,N4573);
and and2657(N4571,N4574,N4575);
and and2664(N4582,N4584,N4585);
and and2665(N4583,N4586,N4587);
and and2672(N4594,N4596,N4597);
and and2673(N4595,N4598,N4599);
and and2680(N4605,N4607,N4608);
and and2681(N4606,N4609,N4610);
and and2688(N4616,N4618,N4619);
and and2689(N4617,N4620,N4621);
and and2696(N4627,N4629,N4630);
and and2697(N4628,N4631,N4632);
and and2704(N4638,N4640,N4641);
and and2705(N4639,N4642,N4643);
and and2712(N4649,N4651,N4652);
and and2713(N4650,N4653,N4654);
and and2720(N4660,N4662,N4663);
and and2721(N4661,N4664,N4665);
and and2728(N4671,N4673,N4674);
and and2729(N4672,N4675,N4676);
and and2736(N4682,N4684,N4685);
and and2737(N4683,N4686,N4687);
and and2744(N4693,N4695,N4696);
and and2745(N4694,N4697,N4698);
and and2752(N4704,N4706,N4707);
and and2753(N4705,N4708,N4709);
and and2760(N4715,N4717,N4718);
and and2761(N4716,N4719,N4720);
and and2768(N4726,N4728,N4729);
and and2769(N4727,N4730,N4731);
and and2776(N4737,N4739,N4740);
and and2777(N4738,N4741,N4742);
and and2784(N4748,N4750,N4751);
and and2785(N4749,N4752,N4753);
and and2792(N4759,N4761,N4762);
and and2793(N4760,N4763,N4764);
and and2800(N4770,N4772,N4773);
and and2801(N4771,N4774,N4775);
and and2808(N4781,N4783,N4784);
and and2809(N4782,N4785,N4786);
and and2816(N4792,N4794,N4795);
and and2817(N4793,N4796,N4797);
and and2824(N4803,N4805,N4806);
and and2825(N4804,N4807,N4808);
and and2832(N4814,N4816,N4817);
and and2833(N4815,N4818,N4819);
and and2840(N4825,N4827,N4828);
and and2841(N4826,N4829,N4830);
and and2848(N4836,N4838,N4839);
and and2849(N4837,N4840,N4841);
and and2856(N4847,N4849,N4850);
and and2857(N4848,N4851,N4852);
and and2864(N4858,N4860,N4861);
and and2865(N4859,N4862,N4863);
and and2872(N4869,N4871,N4872);
and and2873(N4870,N4873,N4874);
and and2880(N4880,N4882,N4883);
and and2881(N4881,N4884,N4885);
and and2888(N4891,N4893,N4894);
and and2889(N4892,N4895,N4896);
and and2896(N4901,N4903,N4904);
and and2897(N4902,N4905,N4906);
and and2904(N4911,N4913,N4914);
and and2905(N4912,N4915,N4916);
and and2912(N4921,N4923,N4924);
and and2913(N4922,N4925,N4926);
and and2920(N4931,N4933,N4934);
and and2921(N4932,N4935,N4936);
and and2928(N4941,N4943,N4944);
and and2929(N4942,N4945,N4946);
and and2936(N4951,N4953,N4954);
and and2937(N4952,N4955,N4956);
and and2944(N4961,N4963,N4964);
and and2945(N4962,N4965,N4966);
and and2952(N4971,N4973,N4974);
and and2953(N4972,N4975,N4976);
and and2960(N4981,N4983,N4984);
and and2961(N4982,N4985,N4986);
and and2968(N4991,N4993,N4994);
and and2969(N4992,N4995,N4996);
and and2976(N5001,N5003,N5004);
and and2977(N5002,N5005,N5006);
and and2984(N5011,N5013,N5014);
and and2985(N5012,N5015,N5016);
and and2992(N5021,N5023,N5024);
and and2993(N5022,N5025,N5026);
and and3000(N5031,N5033,N5034);
and and3001(N5032,N5035,N5036);
and and3008(N5041,N5043,N5044);
and and3009(N5042,N5045,N5046);
and and3016(N5051,N5053,N5054);
and and3017(N5052,N5055,N5056);
and and3024(N5061,N5063,N5064);
and and3025(N5062,N5065,N5066);
and and3032(N5071,N5073,N5074);
and and3033(N5072,N5075,N5076);
and and3040(N5080,N5082,N5083);
and and3041(N5081,N5084,N5085);
and and3048(N5089,N5091,N5092);
and and3049(N5090,N5093,N5094);
and and3056(N5098,N5100,N5101);
and and3057(N5099,N5102,N5103);
and and3064(N5107,N5109,N5110);
and and3065(N5108,N5111,N5112);
and and3072(N5116,N5118,N5119);
and and3073(N5117,N5120,N5121);
and and3080(N5125,N5127,N5128);
and and3081(N5126,N5129,N5130);
and and3087(N5139,N5141,N5142);
and and3088(N5140,N5143,N5144);
and and3094(N5153,N5155,N5156);
and and3095(N5154,N5157,N5158);
and and3101(N5167,N5169,N5170);
and and3102(N5168,N5171,N5172);
and and3108(N5180,N5182,N5183);
and and3109(N5181,N5184,N5185);
and and3115(N5193,N5195,N5196);
and and3116(N5194,N5197,N5198);
and and3122(N5206,N5208,N5209);
and and3123(N5207,N5210,N5211);
and and3129(N5219,N5221,N5222);
and and3130(N5220,N5223,N5224);
and and3136(N5232,N5234,N5235);
and and3137(N5233,N5236,N5237);
and and3143(N5244,N5246,N5247);
and and3144(N5245,N5248,N5249);
and and3150(N5256,N5258,N5259);
and and3151(N5257,N5260,N5261);
and and3157(N5268,N5270,N5271);
and and3158(N5269,N5272,N5273);
and and3164(N5280,N5282,N5283);
and and3165(N5281,N5284,N5285);
and and3171(N5292,N5294,N5295);
and and3172(N5293,N5296,N5297);
and and3178(N5304,N5306,N5307);
and and3179(N5305,N5308,N5309);
and and3185(N5316,N5318,N5319);
and and3186(N5317,N5320,N5321);
and and3192(N5328,N5330,N5331);
and and3193(N5329,N5332,N5333);
and and3199(N5339,N5341,N5342);
and and3200(N5340,N5343,N5344);
and and3206(N5350,N5352,N5353);
and and3207(N5351,N5354,N5355);
and and3213(N5361,N5363,N5364);
and and3214(N5362,N5365,N5366);
and and3220(N5372,N5374,N5375);
and and3221(N5373,N5376,N5377);
and and3227(N5383,N5385,N5386);
and and3228(N5384,N5387,N5388);
and and3234(N5394,N5396,N5397);
and and3235(N5395,N5398,N5399);
and and3241(N5405,N5407,N5408);
and and3242(N5406,N5409,N5410);
and and3248(N5416,N5418,N5419);
and and3249(N5417,N5420,N5421);
and and3255(N5427,N5429,N5430);
and and3256(N5428,N5431,N5432);
and and3262(N5438,N5440,N5441);
and and3263(N5439,N5442,N5443);
and and3269(N5449,N5451,N5452);
and and3270(N5450,N5453,N5454);
and and3276(N5460,N5462,N5463);
and and3277(N5461,N5464,N5465);
and and3283(N5471,N5473,N5474);
and and3284(N5472,N5475,N5476);
and and3290(N5482,N5484,N5485);
and and3291(N5483,N5486,N5487);
and and3297(N5492,N5494,N5495);
and and3298(N5493,N5496,N5497);
and and3304(N5502,N5504,N5505);
and and3305(N5503,N5506,N5507);
and and3311(N5512,N5514,N5515);
and and3312(N5513,N5516,N5517);
and and3318(N5522,N5524,N5525);
and and3319(N5523,N5526,N5527);
and and3325(N5532,N5534,N5535);
and and3326(N5533,N5536,N5537);
and and3332(N5542,N5544,N5545);
and and3333(N5543,N5546,N5547);
and and3339(N5552,N5554,N5555);
and and3340(N5553,N5556,N5557);
and and3346(N5562,N5564,N5565);
and and3347(N5563,N5566,N5567);
and and3353(N5572,N5574,N5575);
and and3354(N5573,N5576,N5577);
and and3360(N5582,N5584,N5585);
and and3361(N5583,N5586,N5587);
and and3367(N5592,N5594,N5595);
and and3368(N5593,N5596,N5597);
and and3374(N5602,N5604,N5605);
and and3375(N5603,N5606,N5607);
and and3381(N5611,N5613,N5614);
and and3382(N5612,N5615,N5616);
and and3388(N5620,N5622,N5623);
and and3389(N5621,N5624,N5625);
and and3395(N5629,N5631,N5632);
and and3396(N5630,N5633,N5634);
and and3402(N5638,N5640,N5641);
and and3403(N5639,N5642,N5643);
and and3409(N5647,N5649,N5650);
and and3410(N5648,N5651,N5652);
and and3416(N5655,N5657,N5658);
and and3417(N5656,N5659,N5660);
and and3(N414,N418,N419);
and and4(N415,N420,N421);
and and5(N416,in2,N422);
and and6(N417,R1,N423);
and and12(N431,N435,N436);
and and13(N432,N437,in2);
and and14(N433,N438,N439);
and and15(N434,N440,N441);
and and21(N448,N452,N453);
and and22(N449,in0,N454);
and and23(N450,N455,N456);
and and24(N451,N457,N458);
and and30(N465,N469,N470);
and and31(N466,in1,N471);
and and32(N467,N472,N473);
and and33(N468,N474,N475);
and and39(N482,N486,N487);
and and40(N483,in1,N488);
and and41(N484,N489,N490);
and and42(N485,N491,R3);
and and48(N499,N503,N504);
and and49(N500,N505,in2);
and and50(N501,N506,N507);
and and51(N502,N508,R3);
and and57(N516,N520,N521);
and and58(N517,N522,N523);
and and59(N518,N524,N525);
and and60(N519,N526,R2);
and and66(N533,N537,N538);
and and67(N534,N539,N540);
and and68(N535,N541,N542);
and and69(N536,N543,R2);
and and75(N550,N554,N555);
and and76(N551,N556,N557);
and and77(N552,N558,N559);
and and78(N553,N560,N561);
and and84(N567,N571,N572);
and and85(N568,N573,N574);
and and86(N569,N575,N576);
and and87(N570,N577,N578);
and and93(N584,N588,N589);
and and94(N585,N590,N591);
and and95(N586,N592,N593);
and and96(N587,N594,R3);
and and102(N601,N605,N606);
and and103(N602,N607,N608);
and and104(N603,N609,N610);
and and105(N604,N611,R2);
and and111(N618,N622,N623);
and and112(N619,N624,in1);
and and113(N620,in2,R0);
and and114(N621,N625,N626);
and and120(N634,N638,N639);
and and121(N635,in0,in1);
and and122(N636,N640,N641);
and and123(N637,N642,N643);
and and129(N650,N654,N655);
and and130(N651,N656,in1);
and and131(N652,in2,N657);
and and132(N653,N658,N659);
and and138(N666,N670,N671);
and and139(N667,N672,N673);
and and140(N668,N674,R1);
and and141(N669,R2,N675);
and and147(N682,N686,N687);
and and148(N683,N688,N689);
and and149(N684,in2,R1);
and and150(N685,R2,N690);
and and156(N698,N702,N703);
and and157(N699,N704,in1);
and and158(N700,R0,N705);
and and159(N701,N706,R3);
and and165(N714,N718,N719);
and and166(N715,N720,N721);
and and167(N716,R0,N722);
and and168(N717,N723,N724);
and and174(N730,N734,N735);
and and175(N731,N736,N737);
and and176(N732,N738,N739);
and and177(N733,N740,R3);
and and183(N746,N750,N751);
and and184(N747,N752,in1);
and and185(N748,N753,N754);
and and186(N749,N755,N756);
and and192(N762,N766,N767);
and and193(N763,N768,N769);
and and194(N764,in2,N770);
and and195(N765,R1,N771);
and and201(N778,N782,N783);
and and202(N779,in0,N784);
and and203(N780,N785,N786);
and and204(N781,N787,N788);
and and210(N794,N798,N799);
and and211(N795,N800,N801);
and and212(N796,in2,N802);
and and213(N797,N803,R2);
and and219(N810,N814,N815);
and and220(N811,N816,N817);
and and221(N812,N818,R1);
and and222(N813,R2,N819);
and and228(N825,N829,N830);
and and229(N826,in0,in1);
and and230(N827,in2,N831);
and and231(N828,N832,N833);
and and237(N840,N844,N845);
and and238(N841,in0,in1);
and and239(N842,R0,N846);
and and240(N843,N847,N848);
and and246(N855,N859,N860);
and and247(N856,N861,N862);
and and248(N857,in2,R0);
and and249(N858,N863,N864);
and and255(N870,N874,N875);
and and256(N871,in0,N876);
and and257(N872,in2,R0);
and and258(N873,N877,N878);
and and264(N885,N889,N890);
and and265(N886,N891,in1);
and and266(N887,in2,R0);
and and267(N888,N892,N893);
and and273(N900,N904,N905);
and and274(N901,N906,in1);
and and275(N902,in2,N907);
and and276(N903,R1,R2);
and and282(N915,N919,N920);
and and283(N916,N921,in2);
and and284(N917,N922,N923);
and and285(N918,N924,N925);
and and291(N930,N934,N935);
and and292(N931,N936,N937);
and and293(N932,in2,R0);
and and294(N933,N938,R3);
and and300(N945,N949,N950);
and and301(N946,in1,N951);
and and302(N947,N952,N953);
and and303(N948,R2,N954);
and and309(N960,N964,N965);
and and310(N961,in0,N966);
and and311(N962,N967,N968);
and and312(N963,R2,N969);
and and318(N975,N979,N980);
and and319(N976,in1,N981);
and and320(N977,N982,N983);
and and321(N978,N984,R3);
and and327(N990,N994,N995);
and and328(N991,N996,N997);
and and329(N992,in2,R0);
and and330(N993,N998,R2);
and and336(N1005,N1009,N1010);
and and337(N1006,N1011,in2);
and and338(N1007,N1012,N1013);
and and339(N1008,R2,R3);
and and345(N1020,N1024,N1025);
and and346(N1021,N1026,N1027);
and and347(N1022,N1028,R1);
and and348(N1023,R2,N1029);
and and354(N1035,N1039,N1040);
and and355(N1036,N1041,in1);
and and356(N1037,N1042,N1043);
and and357(N1038,R2,N1044);
and and363(N1050,N1054,N1055);
and and364(N1051,N1056,N1057);
and and365(N1052,in2,R0);
and and366(N1053,N1058,R2);
and and372(N1065,N1069,N1070);
and and373(N1066,N1071,in1);
and and374(N1067,N1072,R0);
and and375(N1068,N1073,R2);
and and381(N1080,N1084,N1085);
and and382(N1081,N1086,in1);
and and383(N1082,N1087,R0);
and and384(N1083,N1088,N1089);
and and390(N1095,N1099,N1100);
and and391(N1096,N1101,in1);
and and392(N1097,in2,N1102);
and and393(N1098,N1103,N1104);
and and399(N1110,N1114,N1115);
and and400(N1111,N1116,N1117);
and and401(N1112,N1118,R0);
and and402(N1113,N1119,R2);
and and408(N1125,N1129,N1130);
and and409(N1126,N1131,in1);
and and410(N1127,in2,N1132);
and and411(N1128,N1133,N1134);
and and417(N1140,N1144,N1145);
and and418(N1141,N1146,N1147);
and and419(N1142,in2,N1148);
and and420(N1143,R1,R2);
and and426(N1155,N1159,N1160);
and and427(N1156,N1161,N1162);
and and428(N1157,in2,N1163);
and and429(N1158,R2,R3);
and and435(N1170,N1174,N1175);
and and436(N1171,N1176,N1177);
and and437(N1172,R0,R1);
and and438(N1173,N1178,N1179);
and and444(N1185,N1189,N1190);
and and445(N1186,N1191,N1192);
and and446(N1187,N1193,N1194);
and and447(N1188,N1195,R2);
and and453(N1200,N1204,N1205);
and and454(N1201,N1206,in1);
and and455(N1202,N1207,R0);
and and456(N1203,N1208,N1209);
and and462(N1215,N1219,N1220);
and and463(N1216,N1221,N1222);
and and464(N1217,in2,R0);
and and465(N1218,N1223,N1224);
and and471(N1230,N1234,N1235);
and and472(N1231,N1236,N1237);
and and473(N1232,in2,R0);
and and474(N1233,R1,N1238);
and and480(N1245,N1249,N1250);
and and481(N1246,in0,in1);
and and482(N1247,N1251,N1252);
and and483(N1248,N1253,N1254);
and and489(N1260,N1264,N1265);
and and490(N1261,N1266,N1267);
and and491(N1262,N1268,N1269);
and and492(N1263,R1,N1270);
and and498(N1275,N1279,N1280);
and and499(N1276,in0,N1281);
and and500(N1277,in2,N1282);
and and501(N1278,N1283,N1284);
and and507(N1290,N1294,N1295);
and and508(N1291,N1296,in1);
and and509(N1292,in2,N1297);
and and510(N1293,N1298,N1299);
and and516(N1305,N1309,N1310);
and and517(N1306,N1311,N1312);
and and518(N1307,in2,N1313);
and and519(N1308,N1314,R2);
and and525(N1320,N1324,N1325);
and and526(N1321,N1326,in1);
and and527(N1322,N1327,N1328);
and and528(N1323,N1329,R2);
and and534(N1335,N1339,N1340);
and and535(N1336,N1341,N1342);
and and536(N1337,N1343,R0);
and and537(N1338,R1,N1344);
and and543(N1350,N1354,N1355);
and and544(N1351,N1356,in1);
and and545(N1352,N1357,N1358);
and and546(N1353,R2,R3);
and and552(N1364,N1368,N1369);
and and553(N1365,N1370,in1);
and and554(N1366,in2,R0);
and and555(N1367,R1,R2);
and and561(N1378,N1382,N1383);
and and562(N1379,N1384,N1385);
and and563(N1380,in2,R0);
and and564(N1381,N1386,R2);
and and570(N1392,N1396,N1397);
and and571(N1393,N1398,in2);
and and572(N1394,N1399,N1400);
and and573(N1395,N1401,R3);
and and579(N1406,N1410,N1411);
and and580(N1407,in1,N1412);
and and581(N1408,N1413,R1);
and and582(N1409,R2,N1414);
and and588(N1420,N1424,N1425);
and and589(N1421,N1426,N1427);
and and590(N1422,in2,N1428);
and and591(N1423,R1,R2);
and and597(N1434,N1438,N1439);
and and598(N1435,N1440,in1);
and and599(N1436,in2,N1441);
and and600(N1437,R1,R2);
and and606(N1448,N1452,N1453);
and and607(N1449,N1454,N1455);
and and608(N1450,in2,R1);
and and609(N1451,N1456,R3);
and and615(N1462,N1466,N1467);
and and616(N1463,in0,in2);
and and617(N1464,N1468,N1469);
and and618(N1465,N1470,R3);
and and624(N1476,N1480,N1481);
and and625(N1477,N1482,in1);
and and626(N1478,in2,N1483);
and and627(N1479,N1484,R3);
and and633(N1490,N1494,N1495);
and and634(N1491,N1496,N1497);
and and635(N1492,N1498,R0);
and and636(N1493,R1,R2);
and and642(N1504,N1508,N1509);
and and643(N1505,N1510,N1511);
and and644(N1506,R0,N1512);
and and645(N1507,R2,N1513);
and and651(N1518,N1522,N1523);
and and652(N1519,N1524,in2);
and and653(N1520,N1525,R1);
and and654(N1521,N1526,R3);
and and660(N1532,N1536,N1537);
and and661(N1533,N1538,in2);
and and662(N1534,N1539,N1540);
and and663(N1535,R2,N1541);
and and669(N1546,N1550,N1551);
and and670(N1547,N1552,N1553);
and and671(N1548,in2,N1554);
and and672(N1549,R1,R2);
and and678(N1560,N1564,N1565);
and and679(N1561,N1566,in1);
and and680(N1562,in2,R0);
and and681(N1563,N1567,R2);
and and687(N1574,N1578,N1579);
and and688(N1575,N1580,N1581);
and and689(N1576,in2,R0);
and and690(N1577,R1,R2);
and and696(N1588,N1592,N1593);
and and697(N1589,N1594,in1);
and and698(N1590,in2,R0);
and and699(N1591,N1595,N1596);
and and705(N1602,N1606,N1607);
and and706(N1603,N1608,in1);
and and707(N1604,N1609,N1610);
and and708(N1605,N1611,R3);
and and714(N1616,N1620,N1621);
and and715(N1617,N1622,in2);
and and716(N1618,N1623,N1624);
and and717(N1619,R2,N1625);
and and723(N1630,N1634,N1635);
and and724(N1631,N1636,N1637);
and and725(N1632,in2,R0);
and and726(N1633,R1,N1638);
and and732(N1644,N1648,N1649);
and and733(N1645,N1650,in1);
and and734(N1646,N1651,R0);
and and735(N1647,N1652,N1653);
and and741(N1658,N1662,N1663);
and and742(N1659,N1664,in1);
and and743(N1660,in2,R0);
and and744(N1661,N1665,N1666);
and and750(N1672,N1676,N1677);
and and751(N1673,in0,N1678);
and and752(N1674,N1679,N1680);
and and753(N1675,R2,R3);
and and759(N1686,N1690,N1691);
and and760(N1687,in0,N1692);
and and761(N1688,N1693,N1694);
and and762(N1689,N1695,R2);
and and768(N1700,N1704,N1705);
and and769(N1701,N1706,in1);
and and770(N1702,N1707,R0);
and and771(N1703,R1,N1708);
and and777(N1714,N1718,N1719);
and and778(N1715,N1720,N1721);
and and779(N1716,in2,R0);
and and780(N1717,R1,N1722);
and and786(N1728,N1732,N1733);
and and787(N1729,N1734,in2);
and and788(N1730,R0,N1735);
and and789(N1731,R2,R3);
and and795(N1741,N1745,N1746);
and and796(N1742,in0,in2);
and and797(N1743,N1747,N1748);
and and798(N1744,R2,R3);
and and804(N1754,N1758,N1759);
and and805(N1755,N1760,in2);
and and806(N1756,R0,R1);
and and807(N1757,R2,N1761);
and and813(N1767,N1771,N1772);
and and814(N1768,in1,in2);
and and815(N1769,N1773,N1774);
and and816(N1770,R2,R3);
and and822(N1780,N1784,N1785);
and and823(N1781,N1786,in2);
and and824(N1782,R0,N1787);
and and825(N1783,R2,N1788);
and and831(N1793,N1797,N1798);
and and832(N1794,N1799,in1);
and and833(N1795,N1800,R0);
and and834(N1796,N1801,R2);
and and840(N1806,N1810,N1811);
and and841(N1807,in1,in2);
and and842(N1808,R0,R1);
and and843(N1809,R2,N1812);
and and849(N1819,N1823,N1824);
and and850(N1820,in0,N1825);
and and851(N1821,in2,N1826);
and and852(N1822,R1,R2);
and and858(N1832,N1836,N1837);
and and859(N1833,in0,in1);
and and860(N1834,in2,N1838);
and and861(N1835,R2,N1839);
and and867(N1845,N1849,N1850);
and and868(N1846,in1,N1851);
and and869(N1847,R0,N1852);
and and870(N1848,R2,R3);
and and876(N1858,N1862,N1863);
and and877(N1859,in0,in2);
and and878(N1860,N1864,R1);
and and879(N1861,R2,N1865);
and and885(N1871,N1875,N1876);
and and886(N1872,N1877,N1878);
and and887(N1873,R0,N1879);
and and888(N1874,R2,R3);
and and894(N1884,N1888,N1889);
and and895(N1885,N1890,N1891);
and and896(N1886,in2,R0);
and and897(N1887,N1892,N1893);
and and903(N1897,N1901,N1902);
and and904(N1898,in0,in1);
and and905(N1899,in2,R0);
and and906(N1900,R1,N1903);
and and912(N1910,N1914,N1915);
and and913(N1911,in0,in2);
and and914(N1912,R0,N1916);
and and915(N1913,R2,N1917);
and and921(N1923,N1927,N1928);
and and922(N1924,N1929,in1);
and and923(N1925,R0,R1);
and and924(N1926,R2,R3);
and and930(N1936,N1940,N1941);
and and931(N1937,in0,in2);
and and932(N1938,N1942,R1);
and and933(N1939,R2,N1943);
and and939(N1949,N1953,N1954);
and and940(N1950,in0,N1955);
and and941(N1951,R0,R1);
and and942(N1952,R2,R3);
and and948(N1962,N1966,N1967);
and and949(N1963,in0,in1);
and and950(N1964,in2,R0);
and and951(N1965,N1968,R2);
and and957(N1975,N1979,N1980);
and and958(N1976,in0,in1);
and and959(N1977,in2,R0);
and and960(N1978,N1981,N1982);
and and966(N1988,N1992,N1993);
and and967(N1989,N1994,in1);
and and968(N1990,R0,N1995);
and and969(N1991,R2,R3);
and and975(N2001,N2005,N2006);
and and976(N2002,N2007,in2);
and and977(N2003,R0,N2008);
and and978(N2004,R2,R3);
and and984(N2014,N2018,N2019);
and and985(N2015,in0,N2020);
and and986(N2016,R0,N2021);
and and987(N2017,R2,R3);
and and993(N2027,N2031,N2032);
and and994(N2028,N2033,in1);
and and995(N2029,in2,R0);
and and996(N2030,R1,N2034);
and and1002(N2040,N2044,N2045);
and and1003(N2041,N2046,in1);
and and1004(N2042,in2,R0);
and and1005(N2043,N2047,N2048);
and and1011(N2053,N2057,N2058);
and and1012(N2054,N2059,N2060);
and and1013(N2055,in2,R0);
and and1014(N2056,N2061,N2062);
and and1020(N2066,N2070,N2071);
and and1021(N2067,N2072,in1);
and and1022(N2068,N2073,R1);
and and1023(N2069,N2074,R3);
and and1029(N2079,N2083,N2084);
and and1030(N2080,in0,in1);
and and1031(N2081,in2,R0);
and and1032(N2082,N2085,N2086);
and and1038(N2092,N2096,N2097);
and and1039(N2093,in0,N2098);
and and1040(N2094,R0,R1);
and and1041(N2095,N2099,R3);
and and1047(N2105,N2109,N2110);
and and1048(N2106,in0,N2111);
and and1049(N2107,in2,R0);
and and1050(N2108,R1,N2112);
and and1056(N2118,N2122,N2123);
and and1057(N2119,in0,in1);
and and1058(N2120,R0,R1);
and and1059(N2121,N2124,N2125);
and and1065(N2131,N2135,N2136);
and and1066(N2132,N2137,in1);
and and1067(N2133,in2,R0);
and and1068(N2134,R1,N2138);
and and1074(N2144,N2148,N2149);
and and1075(N2145,N2150,N2151);
and and1076(N2146,R0,R1);
and and1077(N2147,R2,N2152);
and and1083(N2157,N2161,N2162);
and and1084(N2158,N2163,N2164);
and and1085(N2159,in2,R1);
and and1086(N2160,R2,N2165);
and and1092(N2170,N2174,N2175);
and and1093(N2171,N2176,in1);
and and1094(N2172,in2,N2177);
and and1095(N2173,N2178,R2);
and and1101(N2183,N2187,N2188);
and and1102(N2184,N2189,N2190);
and and1103(N2185,in2,R0);
and and1104(N2186,N2191,R3);
and and1110(N2196,N2200,N2201);
and and1111(N2197,N2202,in1);
and and1112(N2198,N2203,N2204);
and and1113(N2199,N2205,R2);
and and1119(N2209,N2213,N2214);
and and1120(N2210,in0,in1);
and and1121(N2211,N2215,N2216);
and and1122(N2212,R1,R2);
and and1128(N2222,N2226,N2227);
and and1129(N2223,in0,in1);
and and1130(N2224,N2228,N2229);
and and1131(N2225,N2230,R2);
and and1137(N2235,N2239,N2240);
and and1138(N2236,in1,in2);
and and1139(N2237,R0,R1);
and and1140(N2238,N2241,N2242);
and and1146(N2248,N2252,N2253);
and and1147(N2249,N2254,in2);
and and1148(N2250,N2255,N2256);
and and1149(N2251,R2,R3);
and and1155(N2261,N2265,N2266);
and and1156(N2262,N2267,in1);
and and1157(N2263,in2,N2268);
and and1158(N2264,N2269,N2270);
and and1164(N2274,N2278,N2279);
and and1165(N2275,in0,N2280);
and and1166(N2276,in2,N2281);
and and1167(N2277,N2282,R2);
and and1173(N2287,N2291,N2292);
and and1174(N2288,in0,in1);
and and1175(N2289,N2293,N2294);
and and1176(N2290,N2295,R2);
and and1182(N2300,N2304,N2305);
and and1183(N2301,in0,N2306);
and and1184(N2302,in2,N2307);
and and1185(N2303,N2308,R2);
and and1191(N2313,N2317,N2318);
and and1192(N2314,in0,in1);
and and1193(N2315,N2319,N2320);
and and1194(N2316,N2321,R2);
and and1200(N2326,N2330,N2331);
and and1201(N2327,N2332,in1);
and and1202(N2328,in2,R0);
and and1203(N2329,R1,N2333);
and and1209(N2339,N2343,N2344);
and and1210(N2340,in1,N2345);
and and1211(N2341,R0,R1);
and and1212(N2342,R2,R3);
and and1218(N2351,N2355,N2356);
and and1219(N2352,in1,N2357);
and and1220(N2353,N2358,R1);
and and1221(N2354,R2,R3);
and and1227(N2363,N2367,N2368);
and and1228(N2364,N2369,in1);
and and1229(N2365,in2,N2370);
and and1230(N2366,R1,R2);
and and1236(N2375,N2379,N2380);
and and1237(N2376,in0,in1);
and and1238(N2377,in2,R0);
and and1239(N2378,R1,R2);
and and1245(N2387,N2391,N2392);
and and1246(N2388,N2393,in1);
and and1247(N2389,R0,N2394);
and and1248(N2390,N2395,R3);
and and1254(N2399,N2403,N2404);
and and1255(N2400,N2405,in1);
and and1256(N2401,in2,R0);
and and1257(N2402,N2406,R2);
and and1263(N2411,N2415,N2416);
and and1264(N2412,N2417,N2418);
and and1265(N2413,in2,R1);
and and1266(N2414,R2,R3);
and and1272(N2423,N2427,N2428);
and and1273(N2424,in1,in2);
and and1274(N2425,R0,N2429);
and and1275(N2426,N2430,R3);
and and1281(N2435,N2439,N2440);
and and1282(N2436,N2441,in1);
and and1283(N2437,in2,R0);
and and1284(N2438,N2442,R3);
and and1290(N2447,N2451,N2452);
and and1291(N2448,N2453,in2);
and and1292(N2449,R0,R1);
and and1293(N2450,N2454,R3);
and and1299(N2459,N2463,N2464);
and and1300(N2460,N2465,in2);
and and1301(N2461,R0,R1);
and and1302(N2462,N2466,R3);
and and1308(N2471,N2475,N2476);
and and1309(N2472,in1,in2);
and and1310(N2473,R0,R1);
and and1311(N2474,R2,R3);
and and1317(N2483,N2487,N2488);
and and1318(N2484,in0,in1);
and and1319(N2485,N2489,N2490);
and and1320(N2486,R1,R2);
and and1326(N2495,N2499,N2500);
and and1327(N2496,N2501,in1);
and and1328(N2497,in2,R0);
and and1329(N2498,R1,R2);
and and1335(N2507,N2511,N2512);
and and1336(N2508,in1,in2);
and and1337(N2509,R0,R1);
and and1338(N2510,N2513,R3);
and and1344(N2519,N2523,N2524);
and and1345(N2520,in0,in2);
and and1346(N2521,R0,N2525);
and and1347(N2522,N2526,R3);
and and1353(N2531,N2535,N2536);
and and1354(N2532,in0,in1);
and and1355(N2533,in2,N2537);
and and1356(N2534,R2,R3);
and and1362(N2543,N2547,N2548);
and and1363(N2544,N2549,in1);
and and1364(N2545,in2,R0);
and and1365(N2546,R1,N2550);
and and1371(N2555,N2559,N2560);
and and1372(N2556,in0,N2561);
and and1373(N2557,N2562,R0);
and and1374(N2558,R1,R2);
and and1380(N2567,N2571,N2572);
and and1381(N2568,in0,in1);
and and1382(N2569,in2,R0);
and and1383(N2570,R2,R3);
and and1389(N2578,N2582,N2583);
and and1390(N2579,in1,in2);
and and1391(N2580,N2584,R1);
and and1392(N2581,R2,R3);
and and1398(N2589,N2593,N2594);
and and1399(N2590,in0,in1);
and and1400(N2591,in2,R0);
and and1401(N2592,R1,R2);
and and1407(N2600,N2604,N2605);
and and1408(N2601,in0,in1);
and and1409(N2602,in2,N2606);
and and1410(N2603,R1,R2);
and and1416(N2611,N2615,N2616);
and and1417(N2612,in0,in1);
and and1418(N2613,N2617,N2618);
and and1419(N2614,R2,R3);
and and1425(N2622,N2626,N2627);
and and1426(N2623,in0,in1);
and and1427(N2624,in2,R0);
and and1428(N2625,N2628,R2);
and and1434(N2633,N2637,N2638);
and and1435(N2634,in0,in1);
and and1436(N2635,in2,R0);
and and1437(N2636,R1,N2639);
and and1443(N2644,N2648,N2649);
and and1444(N2645,in0,in1);
and and1445(N2646,in2,R0);
and and1446(N2647,R1,R2);
and and1452(N2655,N2659,N2660);
and and1453(N2656,N2661,in1);
and and1454(N2657,in2,R0);
and and1455(N2658,R1,N2662);
and and1461(N2666,N2670,N2671);
and and1462(N2667,in0,in1);
and and1463(N2668,in2,N2672);
and and1464(N2669,R1,R2);
and and1470(N2677,N2681,N2682);
and and1471(N2678,in0,in1);
and and1472(N2679,in2,R0);
and and1473(N2680,R1,R2);
and and1479(N2688,N2692,N2693);
and and1480(N2689,in0,in1);
and and1481(N2690,in2,R0);
and and1482(N2691,N2694,R2);
and and1488(N2699,N2703,N2704);
and and1489(N2700,in0,in1);
and and1490(N2701,in2,N2705);
and and1491(N2702,R1,N2706);
and and1497(N2710,N2714,N2715);
and and1498(N2711,N2716,in2);
and and1499(N2712,R0,R1);
and and1500(N2713,R2,R3);
and and1506(N2721,N2725,N2726);
and and1507(N2722,in0,in1);
and and1508(N2723,R0,R1);
and and1509(N2724,R2,N2727);
and and1515(N2732,N2736,N2737);
and and1516(N2733,in0,in2);
and and1517(N2734,R0,R1);
and and1518(N2735,R2,N2738);
and and1524(N2743,N2747,N2748);
and and1525(N2744,in0,in1);
and and1526(N2745,N2749,R0);
and and1527(N2746,R1,R2);
and and1533(N2754,N2758,N2759);
and and1534(N2755,in0,in1);
and and1535(N2756,in2,N2760);
and and1536(N2757,N2761,R2);
and and1542(N2765,N2769,N2770);
and and1543(N2766,in0,in1);
and and1544(N2767,in2,R0);
and and1545(N2768,N2771,R2);
and and1551(N2776,N2780,N2781);
and and1552(N2777,in0,in2);
and and1553(N2778,R0,R1);
and and1554(N2779,R2,R3);
and and1560(N2787,N2791,N2792);
and and1561(N2788,in0,in1);
and and1562(N2789,in2,R1);
and and1563(N2790,R2,R3);
and and1569(N2796,N2800,N2801);
and and1570(N2797,in0,in1);
and and1571(N2798,in2,R0);
and and1572(N2799,R1,R2);
and and1578(N2805,N2809,N2810);
and and1579(N2806,N2811,N2812);
and and1580(N2807,N2813,N2814);
and and1581(N2808,N2815,N2816);
and and1586(N2821,N2825,N2826);
and and1587(N2822,N2827,N2828);
and and1588(N2823,R2,N2829);
and and1589(N2824,N2830,N2831);
and and1594(N2837,N2841,N2842);
and and1595(N2838,N2843,N2844);
and and1596(N2839,N2845,N2846);
and and1597(N2840,N2847,R5);
and and1602(N2853,N2857,in0);
and and1603(N2854,N2858,N2859);
and and1604(N2855,N2860,N2861);
and and1605(N2856,N2862,N2863);
and and1610(N2869,N2873,N2874);
and and1611(N2870,N2875,R1);
and and1612(N2871,N2876,N2877);
and and1613(N2872,N2878,N2879);
and and1618(N2884,N2888,in1);
and and1619(N2885,N2889,N2890);
and and1620(N2886,N2891,N2892);
and and1621(N2887,R4,N2893);
and and1626(N2899,N2903,N2904);
and and1627(N2900,N2905,N2906);
and and1628(N2901,R0,R2);
and and1629(N2902,N2907,N2908);
and and1634(N2914,N2918,N2919);
and and1635(N2915,N2920,R0);
and and1636(N2916,N2921,N2922);
and and1637(N2917,R3,N2923);
and and1642(N2929,N2933,N2934);
and and1643(N2930,N2935,R0);
and and1644(N2931,N2936,N2937);
and and1645(N2932,N2938,N2939);
and and1650(N2944,N2948,N2949);
and and1651(N2945,N2950,N2951);
and and1652(N2946,R1,N2952);
and and1653(N2947,N2953,R5);
and and1658(N2959,N2963,N2964);
and and1659(N2960,N2965,N2966);
and and1660(N2961,N2967,N2968);
and and1661(N2962,R3,N2969);
and and1666(N2974,N2978,in0);
and and1667(N2975,in2,R0);
and and1668(N2976,N2979,N2980);
and and1669(N2977,N2981,N2982);
and and1674(N2988,N2992,N2993);
and and1675(N2989,in2,N2994);
and and1676(N2990,N2995,R2);
and and1677(N2991,N2996,N2997);
and and1682(N3002,N3006,in0);
and and1683(N3003,N3007,R0);
and and1684(N3004,N3008,N3009);
and and1685(N3005,N3010,N3011);
and and1690(N3016,N3020,N3021);
and and1691(N3017,N3022,N3023);
and and1692(N3018,R1,R2);
and and1693(N3019,R3,N3024);
and and1698(N3030,N3034,in0);
and and1699(N3031,N3035,N3036);
and and1700(N3032,R1,R2);
and and1701(N3033,N3037,N3038);
and and1706(N3044,N3048,N3049);
and and1707(N3045,in2,R0);
and and1708(N3046,N3050,R2);
and and1709(N3047,N3051,N3052);
and and1714(N3058,N3062,N3063);
and and1715(N3059,N3064,N3065);
and and1716(N3060,N3066,R3);
and and1717(N3061,R4,N3067);
and and1722(N3072,N3076,in0);
and and1723(N3073,N3077,N3078);
and and1724(N3074,N3079,R2);
and and1725(N3075,N3080,N3081);
and and1730(N3086,N3090,in1);
and and1731(N3087,N3091,N3092);
and and1732(N3088,N3093,R2);
and and1733(N3089,N3094,N3095);
and and1738(N3100,N3104,N3105);
and and1739(N3101,in2,N3106);
and and1740(N3102,N3107,R2);
and and1741(N3103,N3108,N3109);
and and1746(N3114,N3118,N3119);
and and1747(N3115,N3120,N3121);
and and1748(N3116,R1,N3122);
and and1749(N3117,N3123,R5);
and and1754(N3128,N3132,in0);
and and1755(N3129,N3133,N3134);
and and1756(N3130,N3135,R2);
and and1757(N3131,N3136,R5);
and and1762(N3142,N3146,in1);
and and1763(N3143,N3147,N3148);
and and1764(N3144,N3149,R2);
and and1765(N3145,N3150,R5);
and and1770(N3156,N3160,N3161);
and and1771(N3157,N3162,N3163);
and and1772(N3158,R1,R3);
and and1773(N3159,R4,N3164);
and and1778(N3170,N3174,N3175);
and and1779(N3171,in1,N3176);
and and1780(N3172,N3177,N3178);
and and1781(N3173,N3179,R5);
and and1786(N3184,N3188,N3189);
and and1787(N3185,N3190,R0);
and and1788(N3186,N3191,N3192);
and and1789(N3187,N3193,N3194);
and and1794(N3198,N3202,in0);
and and1795(N3199,N3203,N3204);
and and1796(N3200,N3205,N3206);
and and1797(N3201,R4,R5);
and and1802(N3212,N3216,N3217);
and and1803(N3213,N3218,R0);
and and1804(N3214,R2,N3219);
and and1805(N3215,R4,N3220);
and and1810(N3226,N3230,N3231);
and and1811(N3227,in1,N3232);
and and1812(N3228,R1,N3233);
and and1813(N3229,N3234,R5);
and and1818(N3240,N3244,N3245);
and and1819(N3241,N3246,R0);
and and1820(N3242,R1,N3247);
and and1821(N3243,N3248,R5);
and and1826(N3254,N3258,N3259);
and and1827(N3255,N3260,in2);
and and1828(N3256,N3261,R3);
and and1829(N3257,N3262,N3263);
and and1834(N3268,N3272,N3273);
and and1835(N3269,N3274,N3275);
and and1836(N3270,N3276,R2);
and and1837(N3271,N3277,R4);
and and1842(N3282,N3286,in0);
and and1843(N3283,N3287,N3288);
and and1844(N3284,R2,N3289);
and and1845(N3285,R4,N3290);
and and1850(N3296,N3300,N3301);
and and1851(N3297,N3302,R0);
and and1852(N3298,R2,N3303);
and and1853(N3299,N3304,N3305);
and and1858(N3310,N3314,N3315);
and and1859(N3311,N3316,R0);
and and1860(N3312,N3317,R3);
and and1861(N3313,N3318,N3319);
and and1866(N3324,N3328,N3329);
and and1867(N3325,N3330,R0);
and and1868(N3326,R1,R3);
and and1869(N3327,N3331,N3332);
and and1874(N3338,N3342,in0);
and and1875(N3339,N3343,N3344);
and and1876(N3340,N3345,R3);
and and1877(N3341,N3346,R5);
and and1882(N3352,N3356,N3357);
and and1883(N3353,N3358,N3359);
and and1884(N3354,N3360,R2);
and and1885(N3355,N3361,R4);
and and1890(N3366,N3370,in0);
and and1891(N3367,N3371,R0);
and and1892(N3368,N3372,N3373);
and and1893(N3369,N3374,N3375);
and and1898(N3380,N3384,in0);
and and1899(N3381,N3385,N3386);
and and1900(N3382,N3387,R1);
and and1901(N3383,R2,N3388);
and and1906(N3394,N3398,N3399);
and and1907(N3395,in2,R1);
and and1908(N3396,N3400,N3401);
and and1909(N3397,N3402,N3403);
and and1914(N3408,N3412,in0);
and and1915(N3409,N3413,R0);
and and1916(N3410,N3414,N3415);
and and1917(N3411,R3,N3416);
and and1922(N3422,N3426,in0);
and and1923(N3423,N3427,R0);
and and1924(N3424,N3428,N3429);
and and1925(N3425,R3,N3430);
and and1930(N3436,N3440,N3441);
and and1931(N3437,in1,N3442);
and and1932(N3438,N3443,R2);
and and1933(N3439,N3444,R5);
and and1938(N3450,N3454,N3455);
and and1939(N3451,N3456,R0);
and and1940(N3452,R2,N3457);
and and1941(N3453,R4,N3458);
and and1946(N3464,N3468,N3469);
and and1947(N3465,R0,N3470);
and and1948(N3466,N3471,N3472);
and and1949(N3467,N3473,N3474);
and and1954(N3478,N3482,in1);
and and1955(N3479,in2,N3483);
and and1956(N3480,R1,R3);
and and1957(N3481,N3484,N3485);
and and1962(N3491,N3495,in0);
and and1963(N3492,N3496,in2);
and and1964(N3493,R1,R3);
and and1965(N3494,N3497,N3498);
and and1970(N3504,N3508,in0);
and and1971(N3505,in1,N3509);
and and1972(N3506,N3510,R1);
and and1973(N3507,R3,N3511);
and and1978(N3517,N3521,in0);
and and1979(N3518,in1,in2);
and and1980(N3519,N3522,N3523);
and and1981(N3520,R2,N3524);
and and1986(N3530,N3534,in0);
and and1987(N3531,in1,in2);
and and1988(N3532,N3535,N3536);
and and1989(N3533,N3537,N3538);
and and1994(N3543,N3547,in0);
and and1995(N3544,N3548,R0);
and and1996(N3545,R1,R2);
and and1997(N3546,N3549,N3550);
and and2002(N3556,N3560,in0);
and and2003(N3557,in1,in2);
and and2004(N3558,N3561,N3562);
and and2005(N3559,R3,N3563);
and and2010(N3569,N3573,N3574);
and and2011(N3570,in1,N3575);
and and2012(N3571,R1,N3576);
and and2013(N3572,N3577,R5);
and and2018(N3582,N3586,N3587);
and and2019(N3583,N3588,in2);
and and2020(N3584,N3589,R1);
and and2021(N3585,N3590,R5);
and and2026(N3595,N3599,in0);
and and2027(N3596,N3600,R0);
and and2028(N3597,N3601,N3602);
and and2029(N3598,N3603,R4);
and and2034(N3608,N3612,N3613);
and and2035(N3609,in1,N3614);
and and2036(N3610,N3615,R1);
and and2037(N3611,R3,R4);
and and2042(N3621,N3625,N3626);
and and2043(N3622,N3627,in2);
and and2044(N3623,N3628,R1);
and and2045(N3624,R3,R4);
and and2050(N3634,N3638,in0);
and and2051(N3635,N3639,R0);
and and2052(N3636,N3640,R2);
and and2053(N3637,N3641,R5);
and and2058(N3647,N3651,in0);
and and2059(N3648,N3652,R0);
and and2060(N3649,N3653,N3654);
and and2061(N3650,N3655,R5);
and and2066(N3660,N3664,N3665);
and and2067(N3661,N3666,R1);
and and2068(N3662,N3667,R3);
and and2069(N3663,R4,R5);
and and2074(N3673,N3677,N3678);
and and2075(N3674,R0,R1);
and and2076(N3675,N3679,N3680);
and and2077(N3676,R4,N3681);
and and2082(N3686,N3690,N3691);
and and2083(N3687,N3692,R0);
and and2084(N3688,N3693,N3694);
and and2085(N3689,N3695,R4);
and and2090(N3699,N3703,N3704);
and and2091(N3700,in2,R0);
and and2092(N3701,N3705,N3706);
and and2093(N3702,R3,R4);
and and2098(N3712,N3716,N3717);
and and2099(N3713,in1,R0);
and and2100(N3714,N3718,N3719);
and and2101(N3715,R3,R4);
and and2106(N3725,N3729,N3730);
and and2107(N3726,N3731,N3732);
and and2108(N3727,N3733,N3734);
and and2109(N3728,R3,R4);
and and2114(N3738,N3742,in0);
and and2115(N3739,in2,N3743);
and and2116(N3740,R1,N3744);
and and2117(N3741,N3745,R5);
and and2122(N3751,N3755,in0);
and and2123(N3752,in1,N3756);
and and2124(N3753,R1,N3757);
and and2125(N3754,N3758,R5);
and and2130(N3764,N3768,N3769);
and and2131(N3765,in1,in2);
and and2132(N3766,N3770,R1);
and and2133(N3767,N3771,N3772);
and and2138(N3777,N3781,N3782);
and and2139(N3778,N3783,N3784);
and and2140(N3779,R2,N3785);
and and2141(N3780,N3786,R5);
and and2146(N3790,N3794,in0);
and and2147(N3791,in2,N3795);
and and2148(N3792,N3796,N3797);
and and2149(N3793,R3,N3798);
and and2154(N3803,N3807,in0);
and and2155(N3804,in2,N3808);
and and2156(N3805,N3809,N3810);
and and2157(N3806,R3,N3811);
and and2162(N3816,N3820,in0);
and and2163(N3817,N3821,N3822);
and and2164(N3818,N3823,R2);
and and2165(N3819,N3824,R4);
and and2170(N3829,N3833,N3834);
and and2171(N3830,in1,in2);
and and2172(N3831,N3835,R2);
and and2173(N3832,N3836,R4);
and and2178(N3842,N3846,in0);
and and2179(N3843,N3847,R0);
and and2180(N3844,N3848,R2);
and and2181(N3845,N3849,N3850);
and and2186(N3855,N3859,in1);
and and2187(N3856,R0,N3860);
and and2188(N3857,R2,N3861);
and and2189(N3858,N3862,N3863);
and and2194(N3868,N3872,N3873);
and and2195(N3869,N3874,R0);
and and2196(N3870,N3875,R2);
and and2197(N3871,N3876,R4);
and and2202(N3881,N3885,N3886);
and and2203(N3882,in1,N3887);
and and2204(N3883,N3888,R1);
and and2205(N3884,R3,N3889);
and and2210(N3894,N3898,in0);
and and2211(N3895,N3899,N3900);
and and2212(N3896,R1,N3901);
and and2213(N3897,R3,N3902);
and and2218(N3907,N3911,in0);
and and2219(N3908,N3912,R0);
and and2220(N3909,R1,R2);
and and2221(N3910,N3913,N3914);
and and2226(N3920,N3924,in0);
and and2227(N3921,in2,N3925);
and and2228(N3922,N3926,R2);
and and2229(N3923,N3927,N3928);
and and2234(N3933,N3937,N3938);
and and2235(N3934,N3939,in2);
and and2236(N3935,R0,R2);
and and2237(N3936,N3940,N3941);
and and2242(N3946,N3950,in0);
and and2243(N3947,in1,N3951);
and and2244(N3948,R0,N3952);
and and2245(N3949,R2,N3953);
and and2250(N3959,N3963,N3964);
and and2251(N3960,N3965,N3966);
and and2252(N3961,R0,R1);
and and2253(N3962,N3967,R5);
and and2258(N3972,N3976,in0);
and and2259(N3973,N3977,N3978);
and and2260(N3974,R2,R3);
and and2261(N3975,R4,R5);
and and2266(N3984,N3988,in0);
and and2267(N3985,in1,N3989);
and and2268(N3986,R1,R2);
and and2269(N3987,N3990,N3991);
and and2274(N3996,N4000,in0);
and and2275(N3997,in1,in2);
and and2276(N3998,R1,R2);
and and2277(N3999,N4001,N4002);
and and2282(N4008,N4012,in0);
and and2283(N4009,N4013,N4014);
and and2284(N4010,N4015,R3);
and and2285(N4011,N4016,R5);
and and2290(N4020,N4024,N4025);
and and2291(N4021,N4026,R0);
and and2292(N4022,R1,R3);
and and2293(N4023,R4,N4027);
and and2298(N4032,N4036,N4037);
and and2299(N4033,N4038,R0);
and and2300(N4034,N4039,R3);
and and2301(N4035,R4,N4040);
and and2306(N4044,N4048,in0);
and and2307(N4045,N4049,R1);
and and2308(N4046,R2,N4050);
and and2309(N4047,N4051,R5);
and and2314(N4056,N4060,N4061);
and and2315(N4057,N4062,R0);
and and2316(N4058,N4063,N4064);
and and2317(N4059,R3,R5);
and and2322(N4068,N4072,in0);
and and2323(N4069,in2,N4073);
and and2324(N4070,R1,R2);
and and2325(N4071,N4074,R5);
and and2330(N4080,N4084,in0);
and and2331(N4081,in1,N4085);
and and2332(N4082,R1,R2);
and and2333(N4083,N4086,R5);
and and2338(N4092,N4096,in1);
and and2339(N4093,in2,R0);
and and2340(N4094,N4097,N4098);
and and2341(N4095,N4099,R4);
and and2346(N4104,N4108,in0);
and and2347(N4105,in1,N4109);
and and2348(N4106,R0,N4110);
and and2349(N4107,N4111,R4);
and and2354(N4116,N4120,in0);
and and2355(N4117,N4121,R0);
and and2356(N4118,R2,N4122);
and and2357(N4119,R4,R5);
and and2362(N4128,N4132,N4133);
and and2363(N4129,R0,N4134);
and and2364(N4130,R2,R3);
and and2365(N4131,R4,N4135);
and and2370(N4140,N4144,in0);
and and2371(N4141,N4145,in2);
and and2372(N4142,R1,N4146);
and and2373(N4143,R3,R4);
and and2378(N4152,N4156,N4157);
and and2379(N4153,in1,in2);
and and2380(N4154,R1,N4158);
and and2381(N4155,R3,R4);
and and2386(N4164,N4168,in0);
and and2387(N4165,N4169,N4170);
and and2388(N4166,R1,R2);
and and2389(N4167,R4,N4171);
and and2394(N4176,N4180,N4181);
and and2395(N4177,N4182,N4183);
and and2396(N4178,R1,R2);
and and2397(N4179,R4,N4184);
and and2402(N4188,N4192,in0);
and and2403(N4189,in1,N4193);
and and2404(N4190,R0,N4194);
and and2405(N4191,N4195,R5);
and and2410(N4200,N4204,in1);
and and2411(N4201,in2,R0);
and and2412(N4202,N4205,N4206);
and and2413(N4203,R4,N4207);
and and2418(N4212,N4216,in1);
and and2419(N4213,N4217,R0);
and and2420(N4214,R1,N4218);
and and2421(N4215,N4219,R4);
and and2426(N4224,N4228,in0);
and and2427(N4225,N4229,R0);
and and2428(N4226,R1,R2);
and and2429(N4227,R4,N4230);
and and2434(N4236,N4240,N4241);
and and2435(N4237,in1,R0);
and and2436(N4238,R1,R2);
and and2437(N4239,R3,N4242);
and and2442(N4248,N4252,N4253);
and and2443(N4249,N4254,R0);
and and2444(N4250,R1,N4255);
and and2445(N4251,R3,N4256);
and and2450(N4260,N4264,in0);
and and2451(N4261,N4265,N4266);
and and2452(N4262,N4267,R2);
and and2453(N4263,R4,N4268);
and and2458(N4272,N4276,in1);
and and2459(N4273,in2,R1);
and and2460(N4274,N4277,R3);
and and2461(N4275,N4278,N4279);
and and2466(N4284,N4288,N4289);
and and2467(N4285,N4290,N4291);
and and2468(N4286,R1,R2);
and and2469(N4287,R4,R5);
and and2474(N4296,N4300,in0);
and and2475(N4297,N4301,N4302);
and and2476(N4298,N4303,R2);
and and2477(N4299,R3,R4);
and and2482(N4308,N4312,in0);
and and2483(N4309,in2,R0);
and and2484(N4310,R1,N4313);
and and2485(N4311,N4314,R5);
and and2490(N4320,N4324,in1);
and and2491(N4321,in2,R0);
and and2492(N4322,R1,N4325);
and and2493(N4323,N4326,R5);
and and2498(N4332,N4336,in0);
and and2499(N4333,N4337,N4338);
and and2500(N4334,R2,R3);
and and2501(N4335,R4,N4339);
and and2506(N4344,N4348,N4349);
and and2507(N4345,in2,N4350);
and and2508(N4346,R1,R2);
and and2509(N4347,R3,N4351);
and and2514(N4356,N4360,N4361);
and and2515(N4357,in2,R0);
and and2516(N4358,R1,N4362);
and and2517(N4359,N4363,R5);
and and2522(N4368,N4372,in1);
and and2523(N4369,in2,N4373);
and and2524(N4370,N4374,R2);
and and2525(N4371,N4375,R4);
and and2530(N4380,N4384,in0);
and and2531(N4381,N4385,in2);
and and2532(N4382,N4386,N4387);
and and2533(N4383,R2,R4);
and and2538(N4392,N4396,N4397);
and and2539(N4393,N4398,N4399);
and and2540(N4394,R2,R3);
and and2541(N4395,R4,R5);
and and2546(N4404,N4408,in0);
and and2547(N4405,N4409,N4410);
and and2548(N4406,N4411,R3);
and and2549(N4407,R4,R5);
and and2554(N4416,N4420,in0);
and and2555(N4417,in1,R0);
and and2556(N4418,N4421,R3);
and and2557(N4419,N4422,N4423);
and and2562(N4428,N4432,in0);
and and2563(N4429,N4433,R1);
and and2564(N4430,N4434,R3);
and and2565(N4431,R4,N4435);
and and2570(N4440,N4444,in0);
and and2571(N4441,in1,N4445);
and and2572(N4442,N4446,N4447);
and and2573(N4443,R2,R4);
and and2578(N4452,N4456,in0);
and and2579(N4453,N4457,R0);
and and2580(N4454,R1,R3);
and and2581(N4455,N4458,R5);
and and2586(N4464,N4468,in1);
and and2587(N4465,in2,N4469);
and and2588(N4466,R1,R2);
and and2589(N4467,R3,N4470);
and and2594(N4476,N4480,in0);
and and2595(N4477,N4481,R1);
and and2596(N4478,R2,N4482);
and and2597(N4479,N4483,R5);
and and2602(N4488,N4492,in0);
and and2603(N4489,in1,R0);
and and2604(N4490,R1,N4493);
and and2605(N4491,R4,N4494);
and and2610(N4500,N4504,in1);
and and2611(N4501,in2,N4505);
and and2612(N4502,R1,N4506);
and and2613(N4503,N4507,R5);
and and2618(N4512,N4516,in0);
and and2619(N4513,in1,in2);
and and2620(N4514,N4517,N4518);
and and2621(N4515,R3,R4);
and and2626(N4524,N4528,in0);
and and2627(N4525,in1,in2);
and and2628(N4526,N4529,N4530);
and and2629(N4527,N4531,R3);
and and2634(N4536,N4540,N4541);
and and2635(N4537,in1,N4542);
and and2636(N4538,R1,R3);
and and2637(N4539,N4543,R5);
and and2642(N4548,N4552,in0);
and and2643(N4549,N4553,R1);
and and2644(N4550,N4554,R3);
and and2645(N4551,R4,R5);
and and2650(N4560,N4564,N4565);
and and2651(N4561,N4566,in2);
and and2652(N4562,N4567,R1);
and and2653(N4563,R3,R4);
and and2658(N4572,N4576,in0);
and and2659(N4573,N4577,N4578);
and and2660(N4574,N4579,R2);
and and2661(N4575,R3,R4);
and and2666(N4584,N4588,in0);
and and2667(N4585,N4589,N4590);
and and2668(N4586,N4591,R3);
and and2669(N4587,R4,R5);
and and2674(N4596,N4600,in1);
and and2675(N4597,in2,R0);
and and2676(N4598,N4601,R2);
and and2677(N4599,N4602,R5);
and and2682(N4607,N4611,N4612);
and and2683(N4608,N4613,N4614);
and and2684(N4609,R2,R3);
and and2685(N4610,R4,R5);
and and2690(N4618,N4622,in1);
and and2691(N4619,R0,R1);
and and2692(N4620,N4623,R3);
and and2693(N4621,R4,N4624);
and and2698(N4629,N4633,in0);
and and2699(N4630,R0,R1);
and and2700(N4631,N4634,R3);
and and2701(N4632,N4635,R5);
and and2706(N4640,N4644,in0);
and and2707(N4641,in1,in2);
and and2708(N4642,R0,N4645);
and and2709(N4643,R2,N4646);
and and2714(N4651,N4655,in0);
and and2715(N4652,in1,in2);
and and2716(N4653,N4656,R2);
and and2717(N4654,R3,N4657);
and and2722(N4662,N4666,N4667);
and and2723(N4663,N4668,in2);
and and2724(N4664,R1,N4669);
and and2725(N4665,R3,R5);
and and2730(N4673,N4677,N4678);
and and2731(N4674,N4679,R0);
and and2732(N4675,R1,R3);
and and2733(N4676,R4,R5);
and and2738(N4684,N4688,in0);
and and2739(N4685,N4689,R1);
and and2740(N4686,R2,R3);
and and2741(N4687,R4,R5);
and and2746(N4695,N4699,in0);
and and2747(N4696,in1,N4700);
and and2748(N4697,R0,R1);
and and2749(N4698,R2,R4);
and and2754(N4706,N4710,N4711);
and and2755(N4707,R0,R1);
and and2756(N4708,R2,R3);
and and2757(N4709,N4712,R5);
and and2762(N4717,N4721,N4722);
and and2763(N4718,N4723,R0);
and and2764(N4719,R1,R2);
and and2765(N4720,R4,N4724);
and and2770(N4728,N4732,in0);
and and2771(N4729,in1,N4733);
and and2772(N4730,R0,N4734);
and and2773(N4731,N4735,R3);
and and2778(N4739,N4743,in0);
and and2779(N4740,in2,N4744);
and and2780(N4741,N4745,N4746);
and and2781(N4742,R3,R4);
and and2786(N4750,N4754,in0);
and and2787(N4751,in1,N4755);
and and2788(N4752,N4756,N4757);
and and2789(N4753,R3,R4);
and and2794(N4761,N4765,N4766);
and and2795(N4762,in2,R0);
and and2796(N4763,R1,R2);
and and2797(N4764,R4,N4767);
and and2802(N4772,N4776,in0);
and and2803(N4773,N4777,N4778);
and and2804(N4774,R0,R1);
and and2805(N4775,R2,R4);
and and2810(N4783,N4787,in0);
and and2811(N4784,in1,in2);
and and2812(N4785,R1,R3);
and and2813(N4786,N4788,N4789);
and and2818(N4794,N4798,in0);
and and2819(N4795,N4799,R0);
and and2820(N4796,R2,N4800);
and and2821(N4797,R4,R5);
and and2826(N4805,N4809,in0);
and and2827(N4806,N4810,R0);
and and2828(N4807,R1,R3);
and and2829(N4808,R4,N4811);
and and2834(N4816,N4820,in0);
and and2835(N4817,N4821,R0);
and and2836(N4818,N4822,R3);
and and2837(N4819,R4,N4823);
and and2842(N4827,N4831,in0);
and and2843(N4828,in2,R0);
and and2844(N4829,N4832,R3);
and and2845(N4830,R4,N4833);
and and2850(N4838,N4842,N4843);
and and2851(N4839,N4844,R0);
and and2852(N4840,R1,R3);
and and2853(N4841,R4,R5);
and and2858(N4849,N4853,in0);
and and2859(N4850,N4854,in2);
and and2860(N4851,N4855,R1);
and and2861(N4852,R2,R3);
and and2866(N4860,N4864,in0);
and and2867(N4861,in1,N4865);
and and2868(N4862,R0,R1);
and and2869(N4863,R3,N4866);
and and2874(N4871,N4875,in0);
and and2875(N4872,in1,N4876);
and and2876(N4873,N4877,R2);
and and2877(N4874,R4,N4878);
and and2882(N4882,N4886,in0);
and and2883(N4883,in1,N4887);
and and2884(N4884,R0,R2);
and and2885(N4885,N4888,R4);
and and2890(N4893,N4897,in0);
and and2891(N4894,N4898,N4899);
and and2892(N4895,R1,R2);
and and2893(N4896,R3,R4);
and and2898(N4903,N4907,in0);
and and2899(N4904,N4908,R0);
and and2900(N4905,R2,R3);
and and2901(N4906,N4909,R5);
and and2906(N4913,N4917,in0);
and and2907(N4914,in2,R0);
and and2908(N4915,N4918,N4919);
and and2909(N4916,R3,R5);
and and2914(N4923,N4927,N4928);
and and2915(N4924,N4929,R1);
and and2916(N4925,R2,R3);
and and2917(N4926,R4,R5);
and and2922(N4933,N4937,N4938);
and and2923(N4934,in1,R1);
and and2924(N4935,R2,N4939);
and and2925(N4936,R4,R5);
and and2930(N4943,N4947,in1);
and and2931(N4944,in2,N4948);
and and2932(N4945,R1,N4949);
and and2933(N4946,R3,R5);
and and2938(N4953,N4957,in0);
and and2939(N4954,in1,N4958);
and and2940(N4955,R0,R1);
and and2941(N4956,R2,R3);
and and2946(N4963,N4967,in0);
and and2947(N4964,in1,R0);
and and2948(N4965,N4968,R3);
and and2949(N4966,R4,R5);
and and2954(N4973,N4977,in0);
and and2955(N4974,N4978,R0);
and and2956(N4975,R1,R2);
and and2957(N4976,R3,R5);
and and2962(N4983,N4987,N4988);
and and2963(N4984,R0,R1);
and and2964(N4985,R2,R3);
and and2965(N4986,R4,R5);
and and2970(N4993,N4997,in0);
and and2971(N4994,N4998,in2);
and and2972(N4995,R1,R2);
and and2973(N4996,R4,R5);
and and2978(N5003,N5007,in0);
and and2979(N5004,in1,N5008);
and and2980(N5005,R1,R2);
and and2981(N5006,R4,R5);
and and2986(N5013,N5017,in1);
and and2987(N5014,in2,N5018);
and and2988(N5015,R1,R2);
and and2989(N5016,R4,R5);
and and2994(N5023,N5027,in0);
and and2995(N5024,in1,in2);
and and2996(N5025,N5028,R2);
and and2997(N5026,R3,R4);
and and3002(N5033,N5037,in0);
and and3003(N5034,in1,in2);
and and3004(N5035,N5038,R2);
and and3005(N5036,R3,R4);
and and3010(N5043,N5047,in0);
and and3011(N5044,in1,in2);
and and3012(N5045,R0,R1);
and and3013(N5046,R3,R5);
and and3018(N5053,N5057,in0);
and and3019(N5054,in1,N5058);
and and3020(N5055,R0,R3);
and and3021(N5056,R4,R5);
and and3026(N5063,N5067,in0);
and and3027(N5064,in2,R0);
and and3028(N5065,R1,R2);
and and3029(N5066,R4,N5068);
and and3034(N5073,N5077,in1);
and and3035(N5074,R0,R1);
and and3036(N5075,R2,R3);
and and3037(N5076,N5078,R5);
and and3042(N5082,N5086,in0);
and and3043(N5083,in1,R0);
and and3044(N5084,R2,R3);
and and3045(N5085,R4,N5087);
and and3050(N5091,N5095,in0);
and and3051(N5092,in2,N5096);
and and3052(N5093,R2,R3);
and and3053(N5094,R4,R5);
and and3058(N5100,N5104,N5105);
and and3059(N5101,in2,R0);
and and3060(N5102,R2,R3);
and and3061(N5103,R4,R5);
and and3066(N5109,N5113,N5114);
and and3067(N5110,in1,R0);
and and3068(N5111,R2,R3);
and and3069(N5112,R4,R5);
and and3074(N5118,N5122,in0);
and and3075(N5119,in2,R0);
and and3076(N5120,R1,R2);
and and3077(N5121,R3,R5);
and and3082(N5127,N5131,R0);
and and3083(N5128,N5132,N5133);
and and3084(N5129,N5134,N5135);
and and3085(N5130,N5136,N5137);
and and3089(N5141,in0,N5145);
and and3090(N5142,N5146,N5147);
and and3091(N5143,N5148,N5149);
and and3092(N5144,N5150,N5151);
and and3096(N5155,in1,N5159);
and and3097(N5156,N5160,N5161);
and and3098(N5157,N5162,N5163);
and and3099(N5158,N5164,N5165);
and and3103(N5169,N5173,R0);
and and3104(N5170,N5174,N5175);
and and3105(N5171,N5176,N5177);
and and3106(N5172,N5178,R7);
and and3110(N5182,in1,N5186);
and and3111(N5183,N5187,R2);
and and3112(N5184,N5188,N5189);
and and3113(N5185,N5190,N5191);
and and3117(N5195,N5199,N5200);
and and3118(N5196,N5201,N5202);
and and3119(N5197,R3,R4);
and and3120(N5198,N5203,N5204);
and and3124(N5208,in0,N5212);
and and3125(N5209,N5213,N5214);
and and3126(N5210,N5215,N5216);
and and3127(N5211,N5217,R7);
and and3131(N5221,in0,N5225);
and and3132(N5222,N5226,N5227);
and and3133(N5223,N5228,N5229);
and and3134(N5224,N5230,R7);
and and3138(N5234,in1,N5238);
and and3139(N5235,N5239,R2);
and and3140(N5236,N5240,N5241);
and and3141(N5237,N5242,R7);
and and3145(N5246,in0,N5250);
and and3146(N5247,N5251,R2);
and and3147(N5248,N5252,N5253);
and and3148(N5249,N5254,R7);
and and3152(N5258,in0,R0);
and and3153(N5259,N5262,R2);
and and3154(N5260,N5263,N5264);
and and3155(N5261,N5265,N5266);
and and3159(N5270,N5274,R0);
and and3160(N5271,R1,N5275);
and and3161(N5272,R4,N5276);
and and3162(N5273,N5277,N5278);
and and3166(N5282,in0,N5286);
and and3167(N5283,N5287,R2);
and and3168(N5284,R3,N5288);
and and3169(N5285,N5289,N5290);
and and3173(N5294,N5298,N5299);
and and3174(N5295,N5300,R3);
and and3175(N5296,R4,N5301);
and and3176(N5297,R6,N5302);
and and3180(N5306,in0,in1);
and and3181(N5307,N5310,N5311);
and and3182(N5308,N5312,N5313);
and and3183(N5309,N5314,R7);
and and3187(N5318,in0,N5322);
and and3188(N5319,N5323,N5324);
and and3189(N5320,R3,R4);
and and3190(N5321,N5325,N5326);
and and3194(N5330,in1,N5334);
and and3195(N5331,R0,R1);
and and3196(N5332,N5335,N5336);
and and3197(N5333,N5337,R7);
and and3201(N5341,in0,N5345);
and and3202(N5342,R0,R1);
and and3203(N5343,N5346,N5347);
and and3204(N5344,N5348,R7);
and and3208(N5352,N5356,R0);
and and3209(N5353,N5357,R3);
and and3210(N5354,R4,N5358);
and and3211(N5355,N5359,R7);
and and3215(N5363,N5367,N5368);
and and3216(N5364,N5369,R1);
and and3217(N5365,R3,N5370);
and and3218(N5366,R5,R6);
and and3222(N5374,in0,R0);
and and3223(N5375,N5378,N5379);
and and3224(N5376,R4,N5380);
and and3225(N5377,R6,N5381);
and and3229(N5385,in0,R0);
and and3230(N5386,N5389,R3);
and and3231(N5387,N5390,N5391);
and and3232(N5388,N5392,R7);
and and3236(N5396,in0,R0);
and and3237(N5397,N5400,R3);
and and3238(N5398,R4,N5401);
and and3239(N5399,N5402,N5403);
and and3243(N5407,in0,R0);
and and3244(N5408,N5411,R2);
and and3245(N5409,N5412,R4);
and and3246(N5410,N5413,N5414);
and and3250(N5418,in0,R1);
and and3251(N5419,N5422,R3);
and and3252(N5420,N5423,N5424);
and and3253(N5421,R6,N5425);
and and3257(N5429,in0,R0);
and and3258(N5430,N5433,N5434);
and and3259(N5431,R4,R5);
and and3260(N5432,N5435,N5436);
and and3264(N5440,N5444,N5445);
and and3265(N5441,R2,R3);
and and3266(N5442,R4,N5446);
and and3267(N5443,R6,N5447);
and and3271(N5451,in0,N5455);
and and3272(N5452,R0,N5456);
and and3273(N5453,R3,N5457);
and and3274(N5454,N5458,R6);
and and3278(N5462,in0,in1);
and and3279(N5463,in2,N5466);
and and3280(N5464,N5467,R2);
and and3281(N5465,N5468,N5469);
and and3285(N5473,N5477,R0);
and and3286(N5474,N5478,R3);
and and3287(N5475,R4,N5479);
and and3288(N5476,N5480,R7);
and and3292(N5484,in0,N5488);
and and3293(N5485,R2,R3);
and and3294(N5486,N5489,R5);
and and3295(N5487,N5490,R7);
and and3299(N5494,in0,R1);
and and3300(N5495,R2,N5498);
and and3301(N5496,N5499,N5500);
and and3302(N5497,R6,R7);
and and3306(N5504,in0,N5508);
and and3307(N5505,R1,R2);
and and3308(N5506,R3,N5509);
and and3309(N5507,R6,N5510);
and and3313(N5514,R0,R1);
and and3314(N5515,R2,N5518);
and and3315(N5516,R4,N5519);
and and3316(N5517,R6,N5520);
and and3320(N5524,in0,in1);
and and3321(N5525,N5528,R0);
and and3322(N5526,R1,N5529);
and and3323(N5527,R5,N5530);
and and3327(N5534,in0,N5538);
and and3328(N5535,N5539,R2);
and and3329(N5536,N5540,R5);
and and3330(N5537,R6,R7);
and and3334(N5544,in0,N5548);
and and3335(N5545,N5549,R0);
and and3336(N5546,R1,R5);
and and3337(N5547,N5550,R7);
and and3341(N5554,in0,N5558);
and and3342(N5555,R0,N5559);
and and3343(N5556,R3,R5);
and and3344(N5557,R6,N5560);
and and3348(N5564,in0,N5568);
and and3349(N5565,R0,N5569);
and and3350(N5566,R3,R5);
and and3351(N5567,N5570,R7);
and and3355(N5574,in0,in1);
and and3356(N5575,R0,R1);
and and3357(N5576,R3,N5578);
and and3358(N5577,N5579,N5580);
and and3362(N5584,in0,N5588);
and and3363(N5585,in2,N5589);
and and3364(N5586,R2,R4);
and and3365(N5587,N5590,R7);
and and3369(N5594,in0,in1);
and and3370(N5595,N5598,R0);
and and3371(N5596,N5599,R2);
and and3372(N5597,N5600,R7);
and and3376(N5604,in0,N5608);
and and3377(N5605,R1,N5609);
and and3378(N5606,R3,R5);
and and3379(N5607,R6,R7);
and and3383(N5613,in0,in2);
and and3384(N5614,R0,R3);
and and3385(N5615,N5617,R5);
and and3386(N5616,N5618,R7);
and and3390(N5622,in0,N5626);
and and3391(N5623,R1,R2);
and and3392(N5624,R3,N5627);
and and3393(N5625,R5,R7);
and and3397(N5631,in0,in2);
and and3398(N5632,N5635,R2);
and and3399(N5633,N5636,R5);
and and3400(N5634,R6,R7);
and and3404(N5640,in0,in1);
and and3405(N5641,N5644,R0);
and and3406(N5642,N5645,R3);
and and3407(N5643,R5,R7);
and and3411(N5649,in0,R0);
and and3412(N5650,R1,R2);
and and3413(N5651,N5653,R4);
and and3414(N5652,R6,R7);
and and3418(N5657,in0,R0);
and and3419(N5658,R1,R3);
and and3420(N5659,R4,R5);
and and3421(N5660,R6,R7);
and and7(N418,N424,N425);
and and8(N419,N426,N427);
and and16(N435,R4,N442);
and and17(N436,N443,N444);
and and25(N452,R4,N459);
and and26(N453,N460,N461);
and and34(N469,N476,R5);
and and35(N470,N477,N478);
and and43(N486,N492,N493);
and and44(N487,N494,N495);
and and52(N503,N509,N510);
and and53(N504,N511,N512);
and and61(N520,N527,N528);
and and62(N521,R6,N529);
and and70(N537,N544,N545);
and and71(N538,R5,N546);
and and79(N554,N562,R5);
and and80(N555,N563,R7);
and and88(N571,R4,R5);
and and89(N572,N579,N580);
and and97(N588,N595,N596);
and and98(N589,N597,R7);
and and106(N605,R4,N612);
and and107(N606,N613,N614);
and and115(N622,N627,N628);
and and116(N623,N629,N630);
and and124(N638,N644,N645);
and and125(N639,R6,N646);
and and133(N654,N660,N661);
and and134(N655,R6,N662);
and and142(N670,N676,N677);
and and143(N671,N678,R7);
and and151(N686,N691,N692);
and and152(N687,N693,N694);
and and160(N702,N707,N708);
and and161(N703,N709,N710);
and and169(N718,R4,N725);
and and170(N719,N726,R7);
and and178(N734,N741,R5);
and and179(N735,N742,R7);
and and187(N750,R4,R5);
and and188(N751,N757,N758);
and and196(N766,N772,R5);
and and197(N767,N773,N774);
and and205(N782,R3,N789);
and and206(N783,N790,R7);
and and214(N798,N804,R4);
and and215(N799,N805,N806);
and and223(N814,R4,R5);
and and224(N815,N820,N821);
and and232(N829,R4,N834);
and and233(N830,N835,N836);
and and241(N844,N849,N850);
and and242(N845,N851,R7);
and and250(N859,N865,R5);
and and251(N860,N866,R7);
and and259(N874,R4,N879);
and and260(N875,N880,N881);
and and268(N889,N894,N895);
and and269(N890,R5,N896);
and and277(N904,N908,N909);
and and278(N905,N910,N911);
and and286(N919,R4,R5);
and and287(N920,N926,R7);
and and295(N934,N939,R5);
and and296(N935,N940,N941);
and and304(N949,N955,R5);
and and305(N950,R6,N956);
and and313(N964,N970,R5);
and and314(N965,R6,N971);
and and322(N979,N985,R5);
and and323(N980,R6,N986);
and and331(N994,N999,N1000);
and and332(N995,N1001,R7);
and and340(N1009,N1014,R5);
and and341(N1010,N1015,N1016);
and and349(N1024,R4,N1030);
and and350(N1025,N1031,R7);
and and358(N1039,N1045,N1046);
and and359(N1040,R6,R7);
and and367(N1054,N1059,R5);
and and368(N1055,N1060,N1061);
and and376(N1069,N1074,N1075);
and and377(N1070,R5,N1076);
and and385(N1084,R4,N1090);
and and386(N1085,R6,N1091);
and and394(N1099,R3,R4);
and and395(N1100,N1105,N1106);
and and403(N1114,R3,N1120);
and and404(N1115,R6,N1121);
and and412(N1129,R4,R5);
and and413(N1130,N1135,N1136);
and and421(N1144,N1149,R4);
and and422(N1145,N1150,N1151);
and and430(N1159,R4,N1164);
and and431(N1160,N1165,N1166);
and and439(N1174,R4,R5);
and and440(N1175,N1180,N1181);
and and448(N1189,R3,R4);
and and449(N1190,N1196,R7);
and and457(N1204,R4,R5);
and and458(N1205,N1210,N1211);
and and466(N1219,N1225,R4);
and and467(N1220,R5,N1226);
and and475(N1234,N1239,R5);
and and476(N1235,N1240,N1241);
and and484(N1249,R3,N1255);
and and485(N1250,N1256,R6);
and and493(N1264,R3,R4);
and and494(N1265,N1271,R7);
and and502(N1279,R3,N1285);
and and503(N1280,R5,N1286);
and and511(N1294,R3,N1300);
and and512(N1295,R5,N1301);
and and520(N1309,R4,N1315);
and and521(N1310,N1316,R7);
and and529(N1324,R4,N1330);
and and530(N1325,N1331,R7);
and and538(N1339,R3,N1345);
and and539(N1340,R5,N1346);
and and547(N1354,R4,R5);
and and548(N1355,N1359,N1360);
and and556(N1368,N1371,N1372);
and and557(N1369,N1373,N1374);
and and565(N1382,R3,N1387);
and and566(N1383,N1388,R7);
and and574(N1396,N1402,R5);
and and575(N1397,R6,R7);
and and583(N1410,N1415,R5);
and and584(N1411,N1416,R7);
and and592(N1424,N1429,R5);
and and593(N1425,R6,N1430);
and and601(N1438,N1442,N1443);
and and602(N1439,R5,N1444);
and and610(N1452,N1457,R5);
and and611(N1453,R6,N1458);
and and619(N1466,N1471,N1472);
and and620(N1467,R6,R7);
and and628(N1480,N1485,N1486);
and and629(N1481,R6,R7);
and and637(N1494,R3,R4);
and and638(N1495,N1499,N1500);
and and646(N1508,R4,R5);
and and647(N1509,N1514,R7);
and and655(N1522,R4,R5);
and and656(N1523,N1527,N1528);
and and664(N1536,R4,R5);
and and665(N1537,R6,N1542);
and and673(N1550,R3,N1555);
and and674(N1551,R5,N1556);
and and682(N1564,N1568,R4);
and and683(N1565,N1569,N1570);
and and691(N1578,R3,N1582);
and and692(N1579,N1583,N1584);
and and700(N1592,N1597,N1598);
and and701(N1593,R6,R7);
and and709(N1606,R4,R5);
and and710(N1607,R6,N1612);
and and718(N1620,N1626,R5);
and and719(N1621,R6,R7);
and and727(N1634,R3,N1639);
and and728(N1635,N1640,R7);
and and736(N1648,R3,N1654);
and and737(N1649,R5,R7);
and and745(N1662,R3,N1667);
and and746(N1663,R6,N1668);
and and754(N1676,N1681,N1682);
and and755(N1677,R6,R7);
and and763(N1690,R3,N1696);
and and764(N1691,R5,R6);
and and772(N1704,R3,N1709);
and and773(N1705,R5,N1710);
and and781(N1718,R3,N1723);
and and782(N1719,R5,N1724);
and and790(N1732,R4,R5);
and and791(N1733,N1736,N1737);
and and799(N1745,R4,R5);
and and800(N1746,N1749,N1750);
and and808(N1758,R4,R5);
and and809(N1759,N1762,N1763);
and and817(N1771,N1775,R5);
and and818(N1772,N1776,R7);
and and826(N1784,R4,N1789);
and and827(N1785,R6,R7);
and and835(N1797,N1802,R4);
and and836(N1798,R6,R7);
and and844(N1810,N1813,N1814);
and and845(N1811,N1815,R7);
and and853(N1823,R3,R4);
and and854(N1824,N1827,N1828);
and and862(N1836,N1840,R5);
and and863(N1837,R6,N1841);
and and871(N1849,N1853,N1854);
and and872(N1850,R6,R7);
and and880(N1862,N1866,R5);
and and881(N1863,N1867,R7);
and and889(N1875,N1880,R5);
and and890(N1876,R6,R7);
and and898(N1888,R3,R4);
and and899(N1889,R6,R7);
and and907(N1901,N1904,N1905);
and and908(N1902,N1906,R7);
and and916(N1914,R4,R5);
and and917(N1915,N1918,N1919);
and and925(N1927,N1930,N1931);
and and926(N1928,N1932,R7);
and and934(N1940,R4,N1944);
and and935(N1941,N1945,R7);
and and943(N1953,N1956,N1957);
and and944(N1954,R6,N1958);
and and952(N1966,N1969,N1970);
and and953(N1967,R5,N1971);
and and961(N1979,N1983,R5);
and and962(N1980,R6,N1984);
and and970(N1992,R4,N1996);
and and971(N1993,R6,N1997);
and and979(N2005,R4,N2009);
and and980(N2006,R6,N2010);
and and988(N2018,R4,N2022);
and and989(N2019,R6,N2023);
and and997(N2031,R4,N2035);
and and998(N2032,N2036,R7);
and and1006(N2044,N2049,R4);
and and1007(N2045,R5,R6);
and and1015(N2057,R4,R5);
and and1016(N2058,R6,R7);
and and1024(N2070,R4,R5);
and and1025(N2071,N2075,R7);
and and1033(N2083,N2087,N2088);
and and1034(N2084,R6,R7);
and and1042(N2096,N2100,N2101);
and and1043(N2097,R6,R7);
and and1051(N2109,N2113,R4);
and and1052(N2110,R5,N2114);
and and1060(N2122,R4,R5);
and and1061(N2123,N2126,N2127);
and and1069(N2135,N2139,R4);
and and1070(N2136,R5,N2140);
and and1078(N2148,N2153,R5);
and and1079(N2149,R6,R7);
and and1087(N2161,R4,R5);
and and1088(N2162,N2166,R7);
and and1096(N2174,R3,R4);
and and1097(N2175,N2179,R7);
and and1105(N2187,R4,R5);
and and1106(N2188,N2192,R7);
and and1114(N2200,R3,R5);
and and1115(N2201,R6,R7);
and and1123(N2213,R3,N2217);
and and1124(N2214,N2218,R7);
and and1132(N2226,N2231,R5);
and and1133(N2227,R6,R7);
and and1141(N2239,N2243,R5);
and and1142(N2240,N2244,R7);
and and1150(N2252,R4,R5);
and and1151(N2253,R6,N2257);
and and1159(N2265,R3,R4);
and and1160(N2266,R5,R7);
and and1168(N2278,R3,N2283);
and and1169(N2279,R6,R7);
and and1177(N2291,R3,N2296);
and and1178(N2292,R6,R7);
and and1186(N2304,R3,R5);
and and1187(N2305,R6,N2309);
and and1195(N2317,R3,R5);
and and1196(N2318,R6,N2322);
and and1204(N2330,R3,N2334);
and and1205(N2331,R5,N2335);
and and1213(N2343,R4,R5);
and and1214(N2344,N2346,N2347);
and and1222(N2355,R4,N2359);
and and1223(N2356,R6,R7);
and and1231(N2367,R3,N2371);
and and1232(N2368,R6,R7);
and and1240(N2379,N2381,N2382);
and and1241(N2380,R6,N2383);
and and1249(N2391,R4,R5);
and and1250(N2392,R6,R7);
and and1258(N2403,R3,N2407);
and and1259(N2404,R6,R7);
and and1267(N2415,N2419,R5);
and and1268(N2416,R6,R7);
and and1276(N2427,R4,N2431);
and and1277(N2428,R6,R7);
and and1285(N2439,N2443,R5);
and and1286(N2440,R6,R7);
and and1294(N2451,R4,R5);
and and1295(N2452,N2455,R7);
and and1303(N2463,R4,N2467);
and and1304(N2464,R6,R7);
and and1312(N2475,N2477,N2478);
and and1313(N2476,R6,N2479);
and and1321(N2487,R3,R4);
and and1322(N2488,R5,N2491);
and and1330(N2499,R3,R4);
and and1331(N2500,N2502,N2503);
and and1339(N2511,N2514,N2515);
and and1340(N2512,R6,R7);
and and1348(N2523,R4,R5);
and and1349(N2524,N2527,R7);
and and1357(N2535,N2538,N2539);
and and1358(N2536,R6,R7);
and and1366(N2547,R3,R5);
and and1367(N2548,N2551,R7);
and and1375(N2559,R3,N2563);
and and1376(N2560,R6,R7);
and and1384(N2571,R4,R5);
and and1385(N2572,N2573,N2574);
and and1393(N2582,R4,R5);
and and1394(N2583,R6,N2585);
and and1402(N2593,N2595,R4);
and and1403(N2594,R5,N2596);
and and1411(N2604,R3,R4);
and and1412(N2605,N2607,R7);
and and1420(N2615,R4,R5);
and and1421(N2616,R6,R7);
and and1429(N2626,R3,N2629);
and and1430(N2627,R6,R7);
and and1438(N2637,R4,R5);
and and1439(N2638,N2640,R7);
and and1447(N2648,N2650,R5);
and and1448(N2649,N2651,R7);
and and1456(N2659,R3,R4);
and and1457(N2660,R5,R6);
and and1465(N2670,R3,R4);
and and1466(N2671,R5,N2673);
and and1474(N2681,R3,R4);
and and1475(N2682,N2683,N2684);
and and1483(N2692,R3,R4);
and and1484(N2693,R6,N2695);
and and1492(N2703,R3,R4);
and and1493(N2704,R5,R7);
and and1501(N2714,R4,N2717);
and and1502(N2715,R6,R7);
and and1510(N2725,R4,R5);
and and1511(N2726,N2728,R7);
and and1519(N2736,N2739,R5);
and and1520(N2737,R6,R7);
and and1528(N2747,N2750,R5);
and and1529(N2748,R6,R7);
and and1537(N2758,R3,R5);
and and1538(N2759,R6,R7);
and and1546(N2769,N2772,R4);
and and1547(N2770,R5,R6);
and and1555(N2780,N2782,N2783);
and and1556(N2781,R6,R7);
and and1564(N2791,R4,R5);
and and1565(N2792,R6,R7);
and and1573(N2800,R3,R4);
and and1574(N2801,R5,R7);
and and1582(N2809,R6,N2817);
and and1590(N2825,N2832,N2833);
and and1598(N2841,N2848,N2849);
and and1606(N2857,N2864,N2865);
and and1614(N2873,N2880,R7);
and and1622(N2888,N2894,N2895);
and and1630(N2903,N2909,N2910);
and and1638(N2918,N2924,N2925);
and and1646(N2933,R6,N2940);
and and1654(N2948,N2954,N2955);
and and1662(N2963,R6,N2970);
and and1670(N2978,N2983,N2984);
and and1678(N2992,N2998,R7);
and and1686(N3006,R5,N3012);
and and1694(N3020,N3025,N3026);
and and1702(N3034,N3039,N3040);
and and1710(N3048,N3053,N3054);
and and1718(N3062,N3068,R7);
and and1726(N3076,R6,N3082);
and and1734(N3090,R6,N3096);
and and1742(N3104,R6,N3110);
and and1750(N3118,N3124,R7);
and and1758(N3132,N3137,N3138);
and and1766(N3146,N3151,N3152);
and and1774(N3160,N3165,N3166);
and and1782(N3174,N3180,R7);
and and1790(N3188,R5,R6);
and and1798(N3202,N3207,N3208);
and and1806(N3216,N3221,N3222);
and and1814(N3230,N3235,N3236);
and and1822(N3244,N3249,N3250);
and and1830(N3258,R6,N3264);
and and1838(N3272,N3278,R6);
and and1846(N3286,N3291,N3292);
and and1854(N3300,R6,N3306);
and and1862(N3314,R6,N3320);
and and1870(N3328,N3333,N3334);
and and1878(N3342,N3347,N3348);
and and1886(N3356,N3362,R7);
and and1894(N3370,R5,N3376);
and and1902(N3384,N3389,N3390);
and and1910(N3398,N3404,R7);
and and1918(N3412,N3417,N3418);
and and1926(N3426,N3431,N3432);
and and1934(N3440,N3445,N3446);
and and1942(N3454,N3459,N3460);
and and1950(N3468,R6,R7);
and and1958(N3482,N3486,N3487);
and and1966(N3495,N3499,N3500);
and and1974(N3508,N3512,N3513);
and and1982(N3521,N3525,N3526);
and and1990(N3534,R5,N3539);
and and1998(N3547,N3551,N3552);
and and2006(N3560,N3564,N3565);
and and2014(N3573,N3578,R7);
and and2022(N3586,N3591,R7);
and and2030(N3599,N3604,R7);
and and2038(N3612,N3616,N3617);
and and2046(N3625,N3629,N3630);
and and2054(N3638,N3642,N3643);
and and2062(N3651,R6,N3656);
and and2070(N3664,N3668,N3669);
and and2078(N3677,N3682,R7);
and and2086(N3690,R5,R6);
and and2094(N3703,N3707,N3708);
and and2102(N3716,N3720,N3721);
and and2110(N3729,R5,R6);
and and2118(N3742,N3746,N3747);
and and2126(N3755,N3759,N3760);
and and2134(N3768,R5,N3773);
and and2142(N3781,R6,R7);
and and2150(N3794,R6,N3799);
and and2158(N3807,N3812,R7);
and and2166(N3820,R6,N3825);
and and2174(N3833,N3837,N3838);
and and2182(N3846,N3851,R6);
and and2190(N3859,R6,N3864);
and and2198(N3872,N3877,R7);
and and2206(N3885,N3890,R7);
and and2214(N3898,N3903,R7);
and and2222(N3911,N3915,N3916);
and and2230(N3924,R6,N3929);
and and2238(N3937,R6,N3942);
and and2246(N3950,N3954,N3955);
and and2254(N3963,N3968,R7);
and and2262(N3976,N3979,N3980);
and and2270(N3988,N3992,R7);
and and2278(N4000,N4003,N4004);
and and2286(N4012,R6,R7);
and and2294(N4024,R6,N4028);
and and2302(N4036,R6,R7);
and and2310(N4048,R6,N4052);
and and2318(N4060,R6,R7);
and and2326(N4072,N4075,N4076);
and and2334(N4084,N4087,N4088);
and and2342(N4096,N4100,R7);
and and2350(N4108,N4112,R7);
and and2358(N4120,N4123,N4124);
and and2366(N4132,N4136,R7);
and and2374(N4144,N4147,N4148);
and and2382(N4156,N4159,N4160);
and and2390(N4168,N4172,R7);
and and2398(N4180,R6,R7);
and and2406(N4192,R6,N4196);
and and2414(N4204,R6,N4208);
and and2422(N4216,N4220,R7);
and and2430(N4228,N4231,N4232);
and and2438(N4240,N4243,N4244);
and and2446(N4252,R6,R7);
and and2454(N4264,R6,R7);
and and2462(N4276,R6,N4280);
and and2470(N4288,N4292,R7);
and and2478(N4300,N4304,R7);
and and2486(N4312,N4315,N4316);
and and2494(N4324,N4327,N4328);
and and2502(N4336,R6,N4340);
and and2510(N4348,N4352,R7);
and and2518(N4360,N4364,R7);
and and2526(N4372,R6,N4376);
and and2534(N4384,N4388,R6);
and and2542(N4396,R6,N4400);
and and2550(N4408,N4412,R7);
and and2558(N4420,R6,N4424);
and and2566(N4432,N4436,R7);
and and2574(N4444,N4448,R7);
and and2582(N4456,N4459,N4460);
and and2590(N4468,N4471,N4472);
and and2598(N4480,R6,N4484);
and and2606(N4492,N4495,N4496);
and and2614(N4504,N4508,R7);
and and2622(N4516,N4519,N4520);
and and2630(N4528,N4532,R7);
and and2638(N4540,R6,N4544);
and and2646(N4552,N4555,N4556);
and and2654(N4564,N4568,R7);
and and2662(N4576,R6,N4580);
and and2670(N4588,N4592,R7);
and and2678(N4600,N4603,R7);
and and2686(N4611,R6,R7);
and and2694(N4622,R6,N4625);
and and2702(N4633,R6,N4636);
and and2710(N4644,N4647,R7);
and and2718(N4655,R5,N4658);
and and2726(N4666,R6,R7);
and and2734(N4677,R6,N4680);
and and2742(N4688,N4690,N4691);
and and2750(N4699,N4701,N4702);
and and2758(N4710,R6,N4713);
and and2766(N4721,R6,R7);
and and2774(N4732,R6,R7);
and and2782(N4743,R5,R6);
and and2790(N4754,R5,R6);
and and2798(N4765,N4768,R7);
and and2806(N4776,N4779,R7);
and and2814(N4787,N4790,R7);
and and2822(N4798,R6,N4801);
and and2830(N4809,R6,N4812);
and and2838(N4820,R6,R7);
and and2846(N4831,N4834,R7);
and and2854(N4842,R6,N4845);
and and2862(N4853,R6,N4856);
and and2870(N4864,N4867,R7);
and and2878(N4875,R6,R7);
and and2886(N4886,R5,N4889);
and and2894(N4897,R6,R7);
and and2902(N4907,R6,R7);
and and2910(N4917,R6,R7);
and and2918(N4927,R6,R7);
and and2926(N4937,R6,R7);
and and2934(N4947,R6,R7);
and and2942(N4957,R6,N4959);
and and2950(N4967,R6,N4969);
and and2958(N4977,R6,N4979);
and and2966(N4987,N4989,R7);
and and2974(N4997,N4999,R7);
and and2982(N5007,N5009,R7);
and and2990(N5017,N5019,R7);
and and2998(N5027,N5029,R7);
and and3006(N5037,R6,N5039);
and and3014(N5047,N5048,N5049);
and and3022(N5057,N5059,R7);
and and3030(N5067,N5069,R7);
and and3038(N5077,R6,R7);
and and3046(N5086,R6,R7);
and and3054(N5095,R6,R7);
and and3062(N5104,R6,R7);
and and3070(N5113,R6,R7);
and and3078(N5122,R6,N5123);
and and3422(N5844,N5845,N5846);
and and3432(N5860,N5861,N5862);
and and3442(N5875,N5876,N5877);
and and3451(N5892,N5893,N5894);
and and3460(N5909,N5910,N5911);
and and3469(N5926,N5927,N5928);
and and3478(N5943,N5944,N5945);
and and3487(N5960,N5961,N5962);
and and3496(N5977,N5978,N5979);
and and3505(N5994,N5995,N5996);
and and3514(N6011,N6012,N6013);
and and3523(N6028,N6029,N6030);
and and3532(N6045,N6046,N6047);
and and3541(N6062,N6063,N6064);
and and3550(N6078,N6079,N6080);
and and3559(N6094,N6095,N6096);
and and3568(N6110,N6111,N6112);
and and3577(N6126,N6127,N6128);
and and3586(N6142,N6143,N6144);
and and3595(N6158,N6159,N6160);
and and3604(N6174,N6175,N6176);
and and3613(N6190,N6191,N6192);
and and3622(N6206,N6207,N6208);
and and3631(N6222,N6223,N6224);
and and3640(N6238,N6239,N6240);
and and3649(N6254,N6255,N6256);
and and3658(N6270,N6271,N6272);
and and3667(N6286,N6287,N6288);
and and3676(N6301,N6302,N6303);
and and3685(N6316,N6317,N6318);
and and3694(N6331,N6332,N6333);
and and3703(N6346,N6347,N6348);
and and3712(N6361,N6362,N6363);
and and3721(N6376,N6377,N6378);
and and3730(N6391,N6392,N6393);
and and3739(N6406,N6407,N6408);
and and3748(N6421,N6422,N6423);
and and3757(N6436,N6437,N6438);
and and3766(N6451,N6452,N6453);
and and3775(N6466,N6467,N6468);
and and3784(N6481,N6482,N6483);
and and3793(N6496,N6497,N6498);
and and3802(N6511,N6512,N6513);
and and3811(N6526,N6527,N6528);
and and3820(N6541,N6542,N6543);
and and3829(N6556,N6557,N6558);
and and3838(N6571,N6572,N6573);
and and3847(N6586,N6587,N6588);
and and3856(N6601,N6602,N6603);
and and3865(N6616,N6617,N6618);
and and3874(N6631,N6632,N6633);
and and3883(N6646,N6647,N6648);
and and3892(N6661,N6662,N6663);
and and3901(N6676,N6677,N6678);
and and3910(N6691,N6692,N6693);
and and3919(N6706,N6707,N6708);
and and3928(N6721,N6722,N6723);
and and3937(N6736,N6737,N6738);
and and3946(N6751,N6752,N6753);
and and3955(N6766,N6767,N6768);
and and3964(N6781,N6782,N6783);
and and3973(N6796,N6797,N6798);
and and3982(N6811,N6812,N6813);
and and3991(N6826,N6827,N6828);
and and4000(N6841,N6842,N6843);
and and4009(N6856,N6857,N6858);
and and4018(N6871,N6872,N6873);
and and4027(N6886,N6887,N6888);
and and4036(N6901,N6902,N6903);
and and4045(N6916,N6917,N6918);
and and4054(N6931,N6932,N6933);
and and4063(N6946,N6947,N6948);
and and4072(N6960,N6961,N6962);
and and4081(N6974,N6975,N6976);
and and4090(N6988,N6989,N6990);
and and4099(N7002,N7003,N7004);
and and4108(N7016,N7017,N7018);
and and4117(N7030,N7031,N7032);
and and4126(N7044,N7045,N7046);
and and4135(N7058,N7059,N7060);
and and4144(N7072,N7073,N7074);
and and4153(N7086,N7087,N7088);
and and4162(N7100,N7101,N7102);
and and4171(N7114,N7115,N7116);
and and4180(N7128,N7129,N7130);
and and4189(N7142,N7143,N7144);
and and4198(N7156,N7157,N7158);
and and4207(N7170,N7171,N7172);
and and4216(N7184,N7185,N7186);
and and4225(N7198,N7199,N7200);
and and4234(N7212,N7213,N7214);
and and4243(N7226,N7227,N7228);
and and4252(N7240,N7241,N7242);
and and4261(N7254,N7255,N7256);
and and4270(N7268,N7269,N7270);
and and4279(N7281,N7282,N7283);
and and4288(N7294,N7295,N7296);
and and4297(N7307,N7308,N7309);
and and4306(N7320,N7321,N7322);
and and4315(N7333,N7334,N7335);
and and4324(N7346,N7347,N7348);
and and4333(N7359,N7360,N7361);
and and4342(N7372,N7373,N7374);
and and4351(N7385,N7386,N7387);
and and4360(N7398,N7399,N7400);
and and4369(N7411,N7412,N7413);
and and4378(N7424,N7425,N7426);
and and4387(N7437,N7438,N7439);
and and4396(N7450,N7451,N7452);
and and4405(N7463,N7464,N7465);
and and4414(N7476,N7477,N7478);
and and4423(N7489,N7490,N7491);
and and4432(N7502,N7503,N7504);
and and4441(N7515,N7516,N7517);
and and4450(N7528,N7529,N7530);
and and4459(N7541,N7542,N7543);
and and4468(N7554,N7555,N7556);
and and4477(N7567,N7568,N7569);
and and4486(N7580,N7581,N7582);
and and4495(N7593,N7594,N7595);
and and4504(N7606,N7607,N7608);
and and4513(N7619,N7620,N7621);
and and4522(N7632,N7633,N7634);
and and4531(N7645,N7646,N7647);
and and4540(N7658,N7659,N7660);
and and4549(N7671,N7672,N7673);
and and4558(N7684,N7685,N7686);
and and4567(N7697,N7698,N7699);
and and4576(N7710,N7711,N7712);
and and4585(N7723,N7724,N7725);
and and4594(N7736,N7737,N7738);
and and4603(N7749,N7750,N7751);
and and4612(N7762,N7763,N7764);
and and4621(N7775,N7776,N7777);
and and4630(N7788,N7789,N7790);
and and4639(N7801,N7802,N7803);
and and4648(N7814,N7815,N7816);
and and4657(N7826,N7827,N7828);
and and4666(N7838,N7839,N7840);
and and4675(N7850,N7851,N7852);
and and4684(N7862,N7863,N7864);
and and4693(N7874,N7875,N7876);
and and4702(N7886,N7887,N7888);
and and4711(N7898,N7899,N7900);
and and4720(N7910,N7911,N7912);
and and4729(N7922,N7923,N7924);
and and4738(N7934,N7935,N7936);
and and4747(N7946,N7947,N7948);
and and4756(N7958,N7959,N7960);
and and4765(N7970,N7971,N7972);
and and4774(N7981,N7982,N7983);
and and4783(N7992,N7993,N7994);
and and4792(N8003,N8004,N8005);
and and4801(N8014,N8015,N8016);
and and4810(N8025,N8026,N8027);
and and4819(N8036,N8037,N8038);
and and4828(N8047,N8048,N8049);
and and4837(N8058,N8059,N8060);
and and4846(N8068,N8069,N8070);
and and4854(N8084,N8085,N8086);
and and4862(N8100,N8101,N8102);
and and4870(N8116,N8117,N8118);
and and4878(N8132,N8133,N8134);
and and4886(N8147,N8148,N8149);
and and4894(N8162,N8163,N8164);
and and4902(N8177,N8178,N8179);
and and4910(N8192,N8193,N8194);
and and4918(N8206,N8207,N8208);
and and4926(N8220,N8221,N8222);
and and4934(N8234,N8235,N8236);
and and4942(N8248,N8249,N8250);
and and4950(N8262,N8263,N8264);
and and4958(N8275,N8276,N8277);
and and4966(N8288,N8289,N8290);
and and4974(N8301,N8302,N8303);
and and4982(N8314,N8315,N8316);
and and4990(N8327,N8328,N8329);
and and4998(N8340,N8341,N8342);
and and5006(N8353,N8354,N8355);
and and5014(N8365,N8366,N8367);
and and5022(N8377,N8378,N8379);
and and5030(N8389,N8390,N8391);
and and5038(N8401,N8402,N8403);
and and5046(N8413,N8414,N8415);
and and3423(N5845,N5847,N5848);
and and3424(N5846,N5849,N5850);
and and3433(N5861,N5863,N5864);
and and3434(N5862,N5865,N5866);
and and3443(N5876,N5878,N5879);
and and3444(N5877,N5880,N5881);
and and3452(N5893,N5895,N5896);
and and3453(N5894,N5897,N5898);
and and3461(N5910,N5912,N5913);
and and3462(N5911,N5914,N5915);
and and3470(N5927,N5929,N5930);
and and3471(N5928,N5931,N5932);
and and3479(N5944,N5946,N5947);
and and3480(N5945,N5948,N5949);
and and3488(N5961,N5963,N5964);
and and3489(N5962,N5965,N5966);
and and3497(N5978,N5980,N5981);
and and3498(N5979,N5982,N5983);
and and3506(N5995,N5997,N5998);
and and3507(N5996,N5999,N6000);
and and3515(N6012,N6014,N6015);
and and3516(N6013,N6016,N6017);
and and3524(N6029,N6031,N6032);
and and3525(N6030,N6033,N6034);
and and3533(N6046,N6048,N6049);
and and3534(N6047,N6050,N6051);
and and3542(N6063,N6065,N6066);
and and3543(N6064,N6067,N6068);
and and3551(N6079,N6081,N6082);
and and3552(N6080,N6083,N6084);
and and3560(N6095,N6097,N6098);
and and3561(N6096,N6099,N6100);
and and3569(N6111,N6113,N6114);
and and3570(N6112,N6115,N6116);
and and3578(N6127,N6129,N6130);
and and3579(N6128,N6131,N6132);
and and3587(N6143,N6145,N6146);
and and3588(N6144,N6147,N6148);
and and3596(N6159,N6161,N6162);
and and3597(N6160,N6163,N6164);
and and3605(N6175,N6177,N6178);
and and3606(N6176,N6179,N6180);
and and3614(N6191,N6193,N6194);
and and3615(N6192,N6195,N6196);
and and3623(N6207,N6209,N6210);
and and3624(N6208,N6211,N6212);
and and3632(N6223,N6225,N6226);
and and3633(N6224,N6227,N6228);
and and3641(N6239,N6241,N6242);
and and3642(N6240,N6243,N6244);
and and3650(N6255,N6257,N6258);
and and3651(N6256,N6259,N6260);
and and3659(N6271,N6273,N6274);
and and3660(N6272,N6275,N6276);
and and3668(N6287,N6289,N6290);
and and3669(N6288,N6291,N6292);
and and3677(N6302,N6304,N6305);
and and3678(N6303,N6306,N6307);
and and3686(N6317,N6319,N6320);
and and3687(N6318,N6321,N6322);
and and3695(N6332,N6334,N6335);
and and3696(N6333,N6336,N6337);
and and3704(N6347,N6349,N6350);
and and3705(N6348,N6351,N6352);
and and3713(N6362,N6364,N6365);
and and3714(N6363,N6366,N6367);
and and3722(N6377,N6379,N6380);
and and3723(N6378,N6381,N6382);
and and3731(N6392,N6394,N6395);
and and3732(N6393,N6396,N6397);
and and3740(N6407,N6409,N6410);
and and3741(N6408,N6411,N6412);
and and3749(N6422,N6424,N6425);
and and3750(N6423,N6426,N6427);
and and3758(N6437,N6439,N6440);
and and3759(N6438,N6441,N6442);
and and3767(N6452,N6454,N6455);
and and3768(N6453,N6456,N6457);
and and3776(N6467,N6469,N6470);
and and3777(N6468,N6471,N6472);
and and3785(N6482,N6484,N6485);
and and3786(N6483,N6486,N6487);
and and3794(N6497,N6499,N6500);
and and3795(N6498,N6501,N6502);
and and3803(N6512,N6514,N6515);
and and3804(N6513,N6516,N6517);
and and3812(N6527,N6529,N6530);
and and3813(N6528,N6531,N6532);
and and3821(N6542,N6544,N6545);
and and3822(N6543,N6546,N6547);
and and3830(N6557,N6559,N6560);
and and3831(N6558,N6561,N6562);
and and3839(N6572,N6574,N6575);
and and3840(N6573,N6576,N6577);
and and3848(N6587,N6589,N6590);
and and3849(N6588,N6591,N6592);
and and3857(N6602,N6604,N6605);
and and3858(N6603,N6606,N6607);
and and3866(N6617,N6619,N6620);
and and3867(N6618,N6621,N6622);
and and3875(N6632,N6634,N6635);
and and3876(N6633,N6636,N6637);
and and3884(N6647,N6649,N6650);
and and3885(N6648,N6651,N6652);
and and3893(N6662,N6664,N6665);
and and3894(N6663,N6666,N6667);
and and3902(N6677,N6679,N6680);
and and3903(N6678,N6681,N6682);
and and3911(N6692,N6694,N6695);
and and3912(N6693,N6696,N6697);
and and3920(N6707,N6709,N6710);
and and3921(N6708,N6711,N6712);
and and3929(N6722,N6724,N6725);
and and3930(N6723,N6726,N6727);
and and3938(N6737,N6739,N6740);
and and3939(N6738,N6741,N6742);
and and3947(N6752,N6754,N6755);
and and3948(N6753,N6756,N6757);
and and3956(N6767,N6769,N6770);
and and3957(N6768,N6771,N6772);
and and3965(N6782,N6784,N6785);
and and3966(N6783,N6786,N6787);
and and3974(N6797,N6799,N6800);
and and3975(N6798,N6801,N6802);
and and3983(N6812,N6814,N6815);
and and3984(N6813,N6816,N6817);
and and3992(N6827,N6829,N6830);
and and3993(N6828,N6831,N6832);
and and4001(N6842,N6844,N6845);
and and4002(N6843,N6846,N6847);
and and4010(N6857,N6859,N6860);
and and4011(N6858,N6861,N6862);
and and4019(N6872,N6874,N6875);
and and4020(N6873,N6876,N6877);
and and4028(N6887,N6889,N6890);
and and4029(N6888,N6891,N6892);
and and4037(N6902,N6904,N6905);
and and4038(N6903,N6906,N6907);
and and4046(N6917,N6919,N6920);
and and4047(N6918,N6921,N6922);
and and4055(N6932,N6934,N6935);
and and4056(N6933,N6936,N6937);
and and4064(N6947,N6949,N6950);
and and4065(N6948,N6951,N6952);
and and4073(N6961,N6963,N6964);
and and4074(N6962,N6965,N6966);
and and4082(N6975,N6977,N6978);
and and4083(N6976,N6979,N6980);
and and4091(N6989,N6991,N6992);
and and4092(N6990,N6993,N6994);
and and4100(N7003,N7005,N7006);
and and4101(N7004,N7007,N7008);
and and4109(N7017,N7019,N7020);
and and4110(N7018,N7021,N7022);
and and4118(N7031,N7033,N7034);
and and4119(N7032,N7035,N7036);
and and4127(N7045,N7047,N7048);
and and4128(N7046,N7049,N7050);
and and4136(N7059,N7061,N7062);
and and4137(N7060,N7063,N7064);
and and4145(N7073,N7075,N7076);
and and4146(N7074,N7077,N7078);
and and4154(N7087,N7089,N7090);
and and4155(N7088,N7091,N7092);
and and4163(N7101,N7103,N7104);
and and4164(N7102,N7105,N7106);
and and4172(N7115,N7117,N7118);
and and4173(N7116,N7119,N7120);
and and4181(N7129,N7131,N7132);
and and4182(N7130,N7133,N7134);
and and4190(N7143,N7145,N7146);
and and4191(N7144,N7147,N7148);
and and4199(N7157,N7159,N7160);
and and4200(N7158,N7161,N7162);
and and4208(N7171,N7173,N7174);
and and4209(N7172,N7175,N7176);
and and4217(N7185,N7187,N7188);
and and4218(N7186,N7189,N7190);
and and4226(N7199,N7201,N7202);
and and4227(N7200,N7203,N7204);
and and4235(N7213,N7215,N7216);
and and4236(N7214,N7217,N7218);
and and4244(N7227,N7229,N7230);
and and4245(N7228,N7231,N7232);
and and4253(N7241,N7243,N7244);
and and4254(N7242,N7245,N7246);
and and4262(N7255,N7257,N7258);
and and4263(N7256,N7259,N7260);
and and4271(N7269,N7271,N7272);
and and4272(N7270,N7273,N7274);
and and4280(N7282,N7284,N7285);
and and4281(N7283,N7286,N7287);
and and4289(N7295,N7297,N7298);
and and4290(N7296,N7299,N7300);
and and4298(N7308,N7310,N7311);
and and4299(N7309,N7312,N7313);
and and4307(N7321,N7323,N7324);
and and4308(N7322,N7325,N7326);
and and4316(N7334,N7336,N7337);
and and4317(N7335,N7338,N7339);
and and4325(N7347,N7349,N7350);
and and4326(N7348,N7351,N7352);
and and4334(N7360,N7362,N7363);
and and4335(N7361,N7364,N7365);
and and4343(N7373,N7375,N7376);
and and4344(N7374,N7377,N7378);
and and4352(N7386,N7388,N7389);
and and4353(N7387,N7390,N7391);
and and4361(N7399,N7401,N7402);
and and4362(N7400,N7403,N7404);
and and4370(N7412,N7414,N7415);
and and4371(N7413,N7416,N7417);
and and4379(N7425,N7427,N7428);
and and4380(N7426,N7429,N7430);
and and4388(N7438,N7440,N7441);
and and4389(N7439,N7442,N7443);
and and4397(N7451,N7453,N7454);
and and4398(N7452,N7455,N7456);
and and4406(N7464,N7466,N7467);
and and4407(N7465,N7468,N7469);
and and4415(N7477,N7479,N7480);
and and4416(N7478,N7481,N7482);
and and4424(N7490,N7492,N7493);
and and4425(N7491,N7494,N7495);
and and4433(N7503,N7505,N7506);
and and4434(N7504,N7507,N7508);
and and4442(N7516,N7518,N7519);
and and4443(N7517,N7520,N7521);
and and4451(N7529,N7531,N7532);
and and4452(N7530,N7533,N7534);
and and4460(N7542,N7544,N7545);
and and4461(N7543,N7546,N7547);
and and4469(N7555,N7557,N7558);
and and4470(N7556,N7559,N7560);
and and4478(N7568,N7570,N7571);
and and4479(N7569,N7572,N7573);
and and4487(N7581,N7583,N7584);
and and4488(N7582,N7585,N7586);
and and4496(N7594,N7596,N7597);
and and4497(N7595,N7598,N7599);
and and4505(N7607,N7609,N7610);
and and4506(N7608,N7611,N7612);
and and4514(N7620,N7622,N7623);
and and4515(N7621,N7624,N7625);
and and4523(N7633,N7635,N7636);
and and4524(N7634,N7637,N7638);
and and4532(N7646,N7648,N7649);
and and4533(N7647,N7650,N7651);
and and4541(N7659,N7661,N7662);
and and4542(N7660,N7663,N7664);
and and4550(N7672,N7674,N7675);
and and4551(N7673,N7676,N7677);
and and4559(N7685,N7687,N7688);
and and4560(N7686,N7689,N7690);
and and4568(N7698,N7700,N7701);
and and4569(N7699,N7702,N7703);
and and4577(N7711,N7713,N7714);
and and4578(N7712,N7715,N7716);
and and4586(N7724,N7726,N7727);
and and4587(N7725,N7728,N7729);
and and4595(N7737,N7739,N7740);
and and4596(N7738,N7741,N7742);
and and4604(N7750,N7752,N7753);
and and4605(N7751,N7754,N7755);
and and4613(N7763,N7765,N7766);
and and4614(N7764,N7767,N7768);
and and4622(N7776,N7778,N7779);
and and4623(N7777,N7780,N7781);
and and4631(N7789,N7791,N7792);
and and4632(N7790,N7793,N7794);
and and4640(N7802,N7804,N7805);
and and4641(N7803,N7806,N7807);
and and4649(N7815,N7817,N7818);
and and4650(N7816,N7819,N7820);
and and4658(N7827,N7829,N7830);
and and4659(N7828,N7831,N7832);
and and4667(N7839,N7841,N7842);
and and4668(N7840,N7843,N7844);
and and4676(N7851,N7853,N7854);
and and4677(N7852,N7855,N7856);
and and4685(N7863,N7865,N7866);
and and4686(N7864,N7867,N7868);
and and4694(N7875,N7877,N7878);
and and4695(N7876,N7879,N7880);
and and4703(N7887,N7889,N7890);
and and4704(N7888,N7891,N7892);
and and4712(N7899,N7901,N7902);
and and4713(N7900,N7903,N7904);
and and4721(N7911,N7913,N7914);
and and4722(N7912,N7915,N7916);
and and4730(N7923,N7925,N7926);
and and4731(N7924,N7927,N7928);
and and4739(N7935,N7937,N7938);
and and4740(N7936,N7939,N7940);
and and4748(N7947,N7949,N7950);
and and4749(N7948,N7951,N7952);
and and4757(N7959,N7961,N7962);
and and4758(N7960,N7963,N7964);
and and4766(N7971,N7973,N7974);
and and4767(N7972,N7975,N7976);
and and4775(N7982,N7984,N7985);
and and4776(N7983,N7986,N7987);
and and4784(N7993,N7995,N7996);
and and4785(N7994,N7997,N7998);
and and4793(N8004,N8006,N8007);
and and4794(N8005,N8008,N8009);
and and4802(N8015,N8017,N8018);
and and4803(N8016,N8019,N8020);
and and4811(N8026,N8028,N8029);
and and4812(N8027,N8030,N8031);
and and4820(N8037,N8039,N8040);
and and4821(N8038,N8041,N8042);
and and4829(N8048,N8050,N8051);
and and4830(N8049,N8052,N8053);
and and4838(N8059,N8061,N8062);
and and4839(N8060,N8063,N8064);
and and4847(N8069,N8071,N8072);
and and4848(N8070,N8073,N8074);
and and4855(N8085,N8087,N8088);
and and4856(N8086,N8089,N8090);
and and4863(N8101,N8103,N8104);
and and4864(N8102,N8105,N8106);
and and4871(N8117,N8119,N8120);
and and4872(N8118,N8121,N8122);
and and4879(N8133,N8135,N8136);
and and4880(N8134,N8137,N8138);
and and4887(N8148,N8150,N8151);
and and4888(N8149,N8152,N8153);
and and4895(N8163,N8165,N8166);
and and4896(N8164,N8167,N8168);
and and4903(N8178,N8180,N8181);
and and4904(N8179,N8182,N8183);
and and4911(N8193,N8195,N8196);
and and4912(N8194,N8197,N8198);
and and4919(N8207,N8209,N8210);
and and4920(N8208,N8211,N8212);
and and4927(N8221,N8223,N8224);
and and4928(N8222,N8225,N8226);
and and4935(N8235,N8237,N8238);
and and4936(N8236,N8239,N8240);
and and4943(N8249,N8251,N8252);
and and4944(N8250,N8253,N8254);
and and4951(N8263,N8265,N8266);
and and4952(N8264,N8267,N8268);
and and4959(N8276,N8278,N8279);
and and4960(N8277,N8280,N8281);
and and4967(N8289,N8291,N8292);
and and4968(N8290,N8293,N8294);
and and4975(N8302,N8304,N8305);
and and4976(N8303,N8306,N8307);
and and4983(N8315,N8317,N8318);
and and4984(N8316,N8319,N8320);
and and4991(N8328,N8330,N8331);
and and4992(N8329,N8332,N8333);
and and4999(N8341,N8343,N8344);
and and5000(N8342,N8345,N8346);
and and5007(N8354,N8356,N8357);
and and5008(N8355,N8358,N8359);
and and5015(N8366,N8368,N8369);
and and5016(N8367,N8370,N8371);
and and5023(N8378,N8380,N8381);
and and5024(N8379,N8382,N8383);
and and5031(N8390,N8392,N8393);
and and5032(N8391,N8394,N8395);
and and5039(N8402,N8404,N8405);
and and5040(N8403,N8406,N8407);
and and5047(N8414,N8416,N8417);
and and5048(N8415,N8418,N8419);
and and3425(N5847,N5851,N5852);
and and3426(N5848,N5853,N5854);
and and3427(N5849,in1,in2);
and and3428(N5850,N5855,N5856);
and and3435(N5863,N5867,N5868);
and and3436(N5864,N5869,N5870);
and and3437(N5865,N5871,in2);
and and3438(N5866,R0,R1);
and and3445(N5878,N5882,N5883);
and and3446(N5879,N5884,N5885);
and and3447(N5880,in2,N5886);
and and3448(N5881,R1,N5887);
and and3454(N5895,N5899,N5900);
and and3455(N5896,N5901,in1);
and and3456(N5897,N5902,N5903);
and and3457(N5898,N5904,N5905);
and and3463(N5912,N5916,N5917);
and and3464(N5913,N5918,in1);
and and3465(N5914,in2,N5919);
and and3466(N5915,N5920,N5921);
and and3472(N5929,N5933,N5934);
and and3473(N5930,N5935,N5936);
and and3474(N5931,in2,N5937);
and and3475(N5932,N5938,R2);
and and3481(N5946,N5950,N5951);
and and3482(N5947,N5952,in1);
and and3483(N5948,N5953,N5954);
and and3484(N5949,N5955,R2);
and and3490(N5963,N5967,N5968);
and and3491(N5964,N5969,N5970);
and and3492(N5965,in2,N5971);
and and3493(N5966,N5972,N5973);
and and3499(N5980,N5984,N5985);
and and3500(N5981,N5986,in1);
and and3501(N5982,N5987,N5988);
and and3502(N5983,N5989,N5990);
and and3508(N5997,N6001,N6002);
and and3509(N5998,N6003,N6004);
and and3510(N5999,N6005,R0);
and and3511(N6000,N6006,N6007);
and and3517(N6014,N6018,N6019);
and and3518(N6015,N6020,N6021);
and and3519(N6016,N6022,N6023);
and and3520(N6017,R1,N6024);
and and3526(N6031,N6035,N6036);
and and3527(N6032,N6037,N6038);
and and3528(N6033,N6039,N6040);
and and3529(N6034,N6041,R3);
and and3535(N6048,N6052,N6053);
and and3536(N6049,N6054,N6055);
and and3537(N6050,N6056,N6057);
and and3538(N6051,N6058,R2);
and and3544(N6065,N6069,N6070);
and and3545(N6066,N6071,in1);
and and3546(N6067,in2,N6072);
and and3547(N6068,N6073,N6074);
and and3553(N6081,N6085,N6086);
and and3554(N6082,N6087,in1);
and and3555(N6083,N6088,R0);
and and3556(N6084,N6089,N6090);
and and3562(N6097,N6101,N6102);
and and3563(N6098,N6103,N6104);
and and3564(N6099,in2,R0);
and and3565(N6100,N6105,N6106);
and and3571(N6113,N6117,N6118);
and and3572(N6114,N6119,N6120);
and and3573(N6115,N6121,R1);
and and3574(N6116,R2,R3);
and and3580(N6129,N6133,N6134);
and and3581(N6130,N6135,N6136);
and and3582(N6131,N6137,N6138);
and and3583(N6132,R2,R3);
and and3589(N6145,N6149,N6150);
and and3590(N6146,N6151,in1);
and and3591(N6147,N6152,N6153);
and and3592(N6148,N6154,R2);
and and3598(N6161,N6165,N6166);
and and3599(N6162,N6167,N6168);
and and3600(N6163,N6169,R1);
and and3601(N6164,N6170,R3);
and and3607(N6177,N6181,N6182);
and and3608(N6178,N6183,N6184);
and and3609(N6179,in2,R0);
and and3610(N6180,N6185,N6186);
and and3616(N6193,N6197,N6198);
and and3617(N6194,N6199,N6200);
and and3618(N6195,N6201,R0);
and and3619(N6196,N6202,N6203);
and and3625(N6209,N6213,N6214);
and and3626(N6210,N6215,N6216);
and and3627(N6211,N6217,R1);
and and3628(N6212,N6218,R3);
and and3634(N6225,N6229,N6230);
and and3635(N6226,N6231,N6232);
and and3636(N6227,in2,N6233);
and and3637(N6228,N6234,N6235);
and and3643(N6241,N6245,N6246);
and and3644(N6242,N6247,N6248);
and and3645(N6243,N6249,R0);
and and3646(N6244,R1,N6250);
and and3652(N6257,N6261,N6262);
and and3653(N6258,N6263,in1);
and and3654(N6259,N6264,N6265);
and and3655(N6260,R1,N6266);
and and3661(N6273,N6277,N6278);
and and3662(N6274,N6279,N6280);
and and3663(N6275,N6281,N6282);
and and3664(N6276,R1,N6283);
and and3670(N6289,N6293,N6294);
and and3671(N6290,N6295,N6296);
and and3672(N6291,in2,N6297);
and and3673(N6292,N6298,R2);
and and3679(N6304,N6308,N6309);
and and3680(N6305,N6310,N6311);
and and3681(N6306,N6312,N6313);
and and3682(N6307,R2,N6314);
and and3688(N6319,N6323,N6324);
and and3689(N6320,N6325,in1);
and and3690(N6321,in2,R1);
and and3691(N6322,N6326,N6327);
and and3697(N6334,N6338,N6339);
and and3698(N6335,N6340,N6341);
and and3699(N6336,N6342,R1);
and and3700(N6337,R2,N6343);
and and3706(N6349,N6353,N6354);
and and3707(N6350,N6355,N6356);
and and3708(N6351,R0,N6357);
and and3709(N6352,R2,R3);
and and3715(N6364,N6368,N6369);
and and3716(N6365,N6370,in1);
and and3717(N6366,in2,R0);
and and3718(N6367,N6371,N6372);
and and3724(N6379,N6383,N6384);
and and3725(N6380,N6385,N6386);
and and3726(N6381,N6387,R0);
and and3727(N6382,R1,R2);
and and3733(N6394,N6398,N6399);
and and3734(N6395,N6400,in2);
and and3735(N6396,N6401,R1);
and and3736(N6397,N6402,R3);
and and3742(N6409,N6413,N6414);
and and3743(N6410,N6415,in1);
and and3744(N6411,N6416,N6417);
and and3745(N6412,R2,R3);
and and3751(N6424,N6428,N6429);
and and3752(N6425,N6430,N6431);
and and3753(N6426,N6432,N6433);
and and3754(N6427,N6434,R3);
and and3760(N6439,N6443,N6444);
and and3761(N6440,N6445,N6446);
and and3762(N6441,in2,N6447);
and and3763(N6442,R2,N6448);
and and3769(N6454,N6458,N6459);
and and3770(N6455,N6460,in1);
and and3771(N6456,N6461,N6462);
and and3772(N6457,N6463,R2);
and and3778(N6469,N6473,N6474);
and and3779(N6470,N6475,N6476);
and and3780(N6471,N6477,R1);
and and3781(N6472,R2,N6478);
and and3787(N6484,N6488,N6489);
and and3788(N6485,N6490,N6491);
and and3789(N6486,N6492,N6493);
and and3790(N6487,R1,R2);
and and3796(N6499,N6503,N6504);
and and3797(N6500,N6505,in1);
and and3798(N6501,N6506,R0);
and and3799(N6502,R1,N6507);
and and3805(N6514,N6518,N6519);
and and3806(N6515,N6520,in1);
and and3807(N6516,N6521,R0);
and and3808(N6517,N6522,R2);
and and3814(N6529,N6533,N6534);
and and3815(N6530,N6535,N6536);
and and3816(N6531,in2,R0);
and and3817(N6532,N6537,R2);
and and3823(N6544,N6548,N6549);
and and3824(N6545,N6550,in2);
and and3825(N6546,N6551,R1);
and and3826(N6547,N6552,N6553);
and and3832(N6559,N6563,N6564);
and and3833(N6560,N6565,in1);
and and3834(N6561,in2,N6566);
and and3835(N6562,R2,N6567);
and and3841(N6574,N6578,N6579);
and and3842(N6575,N6580,N6581);
and and3843(N6576,N6582,R0);
and and3844(N6577,N6583,R2);
and and3850(N6589,N6593,N6594);
and and3851(N6590,N6595,N6596);
and and3852(N6591,N6597,R1);
and and3853(N6592,R2,N6598);
and and3859(N6604,N6608,N6609);
and and3860(N6605,N6610,in1);
and and3861(N6606,in2,N6611);
and and3862(N6607,N6612,N6613);
and and3868(N6619,N6623,N6624);
and and3869(N6620,N6625,N6626);
and and3870(N6621,R0,N6627);
and and3871(N6622,N6628,N6629);
and and3877(N6634,N6638,N6639);
and and3878(N6635,N6640,N6641);
and and3879(N6636,N6642,R0);
and and3880(N6637,N6643,R2);
and and3886(N6649,N6653,N6654);
and and3887(N6650,N6655,in1);
and and3888(N6651,N6656,N6657);
and and3889(N6652,N6658,R3);
and and3895(N6664,N6668,N6669);
and and3896(N6665,N6670,in1);
and and3897(N6666,R0,N6671);
and and3898(N6667,R2,N6672);
and and3904(N6679,N6683,N6684);
and and3905(N6680,N6685,N6686);
and and3906(N6681,in2,R0);
and and3907(N6682,N6687,R3);
and and3913(N6694,N6698,N6699);
and and3914(N6695,N6700,N6701);
and and3915(N6696,in2,N6702);
and and3916(N6697,N6703,R2);
and and3922(N6709,N6713,N6714);
and and3923(N6710,N6715,in1);
and and3924(N6711,N6716,N6717);
and and3925(N6712,N6718,R2);
and and3931(N6724,N6728,N6729);
and and3932(N6725,N6730,N6731);
and and3933(N6726,N6732,N6733);
and and3934(N6727,R1,R2);
and and3940(N6739,N6743,N6744);
and and3941(N6740,N6745,N6746);
and and3942(N6741,in2,R0);
and and3943(N6742,N6747,N6748);
and and3949(N6754,N6758,N6759);
and and3950(N6755,N6760,N6761);
and and3951(N6756,in2,N6762);
and and3952(N6757,N6763,R3);
and and3958(N6769,N6773,N6774);
and and3959(N6770,N6775,N6776);
and and3960(N6771,in2,R0);
and and3961(N6772,N6777,N6778);
and and3967(N6784,N6788,N6789);
and and3968(N6785,N6790,in1);
and and3969(N6786,N6791,R0);
and and3970(N6787,R1,N6792);
and and3976(N6799,N6803,N6804);
and and3977(N6800,N6805,N6806);
and and3978(N6801,N6807,R1);
and and3979(N6802,R2,R3);
and and3985(N6814,N6818,N6819);
and and3986(N6815,N6820,in1);
and and3987(N6816,N6821,N6822);
and and3988(N6817,R2,N6823);
and and3994(N6829,N6833,N6834);
and and3995(N6830,N6835,N6836);
and and3996(N6831,N6837,N6838);
and and3997(N6832,N6839,R3);
and and4003(N6844,N6848,N6849);
and and4004(N6845,N6850,in1);
and and4005(N6846,N6851,R0);
and and4006(N6847,N6852,N6853);
and and4012(N6859,N6863,N6864);
and and4013(N6860,N6865,in1);
and and4014(N6861,in2,N6866);
and and4015(N6862,N6867,N6868);
and and4021(N6874,N6878,N6879);
and and4022(N6875,N6880,N6881);
and and4023(N6876,in2,N6882);
and and4024(N6877,N6883,R2);
and and4030(N6889,N6893,N6894);
and and4031(N6890,N6895,N6896);
and and4032(N6891,N6897,N6898);
and and4033(N6892,R2,R3);
and and4039(N6904,N6908,N6909);
and and4040(N6905,N6910,N6911);
and and4041(N6906,N6912,N6913);
and and4042(N6907,R1,R2);
and and4048(N6919,N6923,N6924);
and and4049(N6920,N6925,N6926);
and and4050(N6921,in2,R1);
and and4051(N6922,R2,R3);
and and4057(N6934,N6938,N6939);
and and4058(N6935,N6940,in1);
and and4059(N6936,N6941,R1);
and and4060(N6937,N6942,R3);
and and4066(N6949,N6953,N6954);
and and4067(N6950,N6955,in1);
and and4068(N6951,N6956,N6957);
and and4069(N6952,N6958,R2);
and and4075(N6963,N6967,N6968);
and and4076(N6964,N6969,in1);
and and4077(N6965,in2,R0);
and and4078(N6966,R1,R2);
and and4084(N6977,N6981,N6982);
and and4085(N6978,N6983,in1);
and and4086(N6979,in2,N6984);
and and4087(N6980,R1,R2);
and and4093(N6991,N6995,N6996);
and and4094(N6992,N6997,in1);
and and4095(N6993,in2,N6998);
and and4096(N6994,R2,R3);
and and4102(N7005,N7009,N7010);
and and4103(N7006,N7011,in1);
and and4104(N7007,N7012,R1);
and and4105(N7008,R2,R3);
and and4111(N7019,N7023,N7024);
and and4112(N7020,N7025,N7026);
and and4113(N7021,N7027,N7028);
and and4114(N7022,R2,N7029);
and and4120(N7033,N7037,N7038);
and and4121(N7034,N7039,in1);
and and4122(N7035,in2,R0);
and and4123(N7036,N7040,N7041);
and and4129(N7047,N7051,N7052);
and and4130(N7048,N7053,N7054);
and and4131(N7049,N7055,R0);
and and4132(N7050,R1,R2);
and and4138(N7061,N7065,N7066);
and and4139(N7062,N7067,N7068);
and and4140(N7063,N7069,R0);
and and4141(N7064,N7070,R3);
and and4147(N7075,N7079,N7080);
and and4148(N7076,N7081,in1);
and and4149(N7077,in2,R0);
and and4150(N7078,N7082,N7083);
and and4156(N7089,N7093,N7094);
and and4157(N7090,N7095,N7096);
and and4158(N7091,R0,N7097);
and and4159(N7092,R2,R3);
and and4165(N7103,N7107,N7108);
and and4166(N7104,N7109,in1);
and and4167(N7105,N7110,R0);
and and4168(N7106,R1,R2);
and and4174(N7117,N7121,N7122);
and and4175(N7118,N7123,N7124);
and and4176(N7119,in2,R0);
and and4177(N7120,R1,R2);
and and4183(N7131,N7135,N7136);
and and4184(N7132,N7137,in1);
and and4185(N7133,in2,R0);
and and4186(N7134,N7138,R2);
and and4192(N7145,N7149,N7150);
and and4193(N7146,N7151,N7152);
and and4194(N7147,N7153,R0);
and and4195(N7148,R1,N7154);
and and4201(N7159,N7163,N7164);
and and4202(N7160,N7165,in1);
and and4203(N7161,N7166,R0);
and and4204(N7162,N7167,N7168);
and and4210(N7173,N7177,N7178);
and and4211(N7174,N7179,in1);
and and4212(N7175,in2,R0);
and and4213(N7176,R2,N7180);
and and4219(N7187,N7191,N7192);
and and4220(N7188,N7193,N7194);
and and4221(N7189,in2,R0);
and and4222(N7190,R1,N7195);
and and4228(N7201,N7205,N7206);
and and4229(N7202,N7207,N7208);
and and4230(N7203,N7209,N7210);
and and4231(N7204,N7211,R2);
and and4237(N7215,N7219,N7220);
and and4238(N7216,N7221,in1);
and and4239(N7217,in2,N7222);
and and4240(N7218,N7223,R3);
and and4246(N7229,N7233,N7234);
and and4247(N7230,N7235,N7236);
and and4248(N7231,N7237,R0);
and and4249(N7232,R2,R3);
and and4255(N7243,N7247,N7248);
and and4256(N7244,N7249,in1);
and and4257(N7245,in2,R0);
and and4258(N7246,R1,N7250);
and and4264(N7257,N7261,N7262);
and and4265(N7258,N7263,in1);
and and4266(N7259,in2,R0);
and and4267(N7260,N7264,R2);
and and4273(N7271,N7275,N7276);
and and4274(N7272,N7277,N7278);
and and4275(N7273,R0,R1);
and and4276(N7274,R2,R3);
and and4282(N7284,N7288,N7289);
and and4283(N7285,N7290,N7291);
and and4284(N7286,N7292,R1);
and and4285(N7287,R2,R3);
and and4291(N7297,N7301,N7302);
and and4292(N7298,N7303,N7304);
and and4293(N7299,N7305,R1);
and and4294(N7300,N7306,R3);
and and4300(N7310,N7314,N7315);
and and4301(N7311,N7316,in1);
and and4302(N7312,in2,N7317);
and and4303(N7313,N7318,R2);
and and4309(N7323,N7327,N7328);
and and4310(N7324,N7329,in2);
and and4311(N7325,R0,R1);
and and4312(N7326,R2,N7330);
and and4318(N7336,N7340,N7341);
and and4319(N7337,N7342,in1);
and and4320(N7338,in2,N7343);
and and4321(N7339,R1,R2);
and and4327(N7349,N7353,N7354);
and and4328(N7350,N7355,in1);
and and4329(N7351,in2,R0);
and and4330(N7352,R1,N7356);
and and4336(N7362,N7366,N7367);
and and4337(N7363,N7368,N7369);
and and4338(N7364,in2,N7370);
and and4339(N7365,R1,R2);
and and4345(N7375,N7379,N7380);
and and4346(N7376,N7381,in1);
and and4347(N7377,N7382,R0);
and and4348(N7378,N7383,R2);
and and4354(N7388,N7392,N7393);
and and4355(N7389,N7394,N7395);
and and4356(N7390,in2,R1);
and and4357(N7391,R2,R3);
and and4363(N7401,N7405,N7406);
and and4364(N7402,N7407,in1);
and and4365(N7403,N7408,R1);
and and4366(N7404,R2,R3);
and and4372(N7414,N7418,N7419);
and and4373(N7415,N7420,N7421);
and and4374(N7416,R0,R1);
and and4375(N7417,R2,R3);
and and4381(N7427,N7431,N7432);
and and4382(N7428,N7433,in1);
and and4383(N7429,in2,N7434);
and and4384(N7430,N7435,N7436);
and and4390(N7440,N7444,N7445);
and and4391(N7441,N7446,in1);
and and4392(N7442,in2,R0);
and and4393(N7443,N7447,N7448);
and and4399(N7453,N7457,N7458);
and and4400(N7454,N7459,N7460);
and and4401(N7455,N7461,R0);
and and4402(N7456,R1,R2);
and and4408(N7466,N7470,N7471);
and and4409(N7467,N7472,N7473);
and and4410(N7468,R0,N7474);
and and4411(N7469,R2,R3);
and and4417(N7479,N7483,N7484);
and and4418(N7480,N7485,in2);
and and4419(N7481,R0,R1);
and and4420(N7482,N7486,R3);
and and4426(N7492,N7496,N7497);
and and4427(N7493,N7498,in1);
and and4428(N7494,R0,R1);
and and4429(N7495,N7499,R3);
and and4435(N7505,N7509,N7510);
and and4436(N7506,N7511,N7512);
and and4437(N7507,N7513,R1);
and and4438(N7508,R2,R3);
and and4444(N7518,N7522,N7523);
and and4445(N7519,N7524,in1);
and and4446(N7520,in2,R1);
and and4447(N7521,R2,N7525);
and and4453(N7531,N7535,N7536);
and and4454(N7532,N7537,in1);
and and4455(N7533,N7538,N7539);
and and4456(N7534,R2,N7540);
and and4462(N7544,N7548,N7549);
and and4463(N7545,N7550,in2);
and and4464(N7546,N7551,N7552);
and and4465(N7547,R2,N7553);
and and4471(N7557,N7561,N7562);
and and4472(N7558,N7563,in1);
and and4473(N7559,R0,R1);
and and4474(N7560,R2,R3);
and and4480(N7570,N7574,N7575);
and and4481(N7571,N7576,N7577);
and and4482(N7572,in2,R0);
and and4483(N7573,N7578,R2);
and and4489(N7583,N7587,N7588);
and and4490(N7584,N7589,N7590);
and and4491(N7585,in2,N7591);
and and4492(N7586,R1,R2);
and and4498(N7596,N7600,N7601);
and and4499(N7597,N7602,in1);
and and4500(N7598,N7603,R1);
and and4501(N7599,R2,R3);
and and4507(N7609,N7613,N7614);
and and4508(N7610,N7615,in1);
and and4509(N7611,R0,R1);
and and4510(N7612,R2,R3);
and and4516(N7622,N7626,N7627);
and and4517(N7623,N7628,N7629);
and and4518(N7624,in2,R0);
and and4519(N7625,R2,N7630);
and and4525(N7635,N7639,N7640);
and and4526(N7636,N7641,in1);
and and4527(N7637,N7642,N7643);
and and4528(N7638,R1,N7644);
and and4534(N7648,N7652,N7653);
and and4535(N7649,N7654,in1);
and and4536(N7650,in2,N7655);
and and4537(N7651,R2,N7656);
and and4543(N7661,N7665,N7666);
and and4544(N7662,N7667,N7668);
and and4545(N7663,R0,R1);
and and4546(N7664,R2,N7669);
and and4552(N7674,N7678,N7679);
and and4553(N7675,N7680,N7681);
and and4554(N7676,in2,N7682);
and and4555(N7677,R1,R2);
and and4561(N7687,N7691,N7692);
and and4562(N7688,N7693,in1);
and and4563(N7689,N7694,N7695);
and and4564(N7690,R1,R2);
and and4570(N7700,N7704,N7705);
and and4571(N7701,N7706,in1);
and and4572(N7702,in2,N7707);
and and4573(N7703,R2,R3);
and and4579(N7713,N7717,N7718);
and and4580(N7714,N7719,N7720);
and and4581(N7715,in2,R0);
and and4582(N7716,N7721,R3);
and and4588(N7726,N7730,N7731);
and and4589(N7727,N7732,N7733);
and and4590(N7728,in2,N7734);
and and4591(N7729,R2,R3);
and and4597(N7739,N7743,N7744);
and and4598(N7740,N7745,N7746);
and and4599(N7741,in2,N7747);
and and4600(N7742,R2,R3);
and and4606(N7752,N7756,N7757);
and and4607(N7753,N7758,in1);
and and4608(N7754,in2,N7759);
and and4609(N7755,N7760,R3);
and and4615(N7765,N7769,N7770);
and and4616(N7766,N7771,in1);
and and4617(N7767,in2,R0);
and and4618(N7768,N7772,R3);
and and4624(N7778,N7782,N7783);
and and4625(N7779,N7784,in2);
and and4626(N7780,R0,N7785);
and and4627(N7781,R2,N7786);
and and4633(N7791,N7795,N7796);
and and4634(N7792,N7797,N7798);
and and4635(N7793,in2,R0);
and and4636(N7794,R1,R3);
and and4642(N7804,N7808,N7809);
and and4643(N7805,N7810,in1);
and and4644(N7806,in2,N7811);
and and4645(N7807,N7812,R3);
and and4651(N7817,N7821,N7822);
and and4652(N7818,N7823,N7824);
and and4653(N7819,in2,N7825);
and and4654(N7820,R1,R3);
and and4660(N7829,N7833,N7834);
and and4661(N7830,N7835,in1);
and and4662(N7831,in2,R1);
and and4663(N7832,R2,R3);
and and4669(N7841,N7845,N7846);
and and4670(N7842,N7847,in2);
and and4671(N7843,R0,N7848);
and and4672(N7844,R2,R3);
and and4678(N7853,N7857,N7858);
and and4679(N7854,N7859,in1);
and and4680(N7855,R0,R1);
and and4681(N7856,R2,N7860);
and and4687(N7865,N7869,N7870);
and and4688(N7866,N7871,in1);
and and4689(N7867,N7872,R0);
and and4690(N7868,R1,R3);
and and4696(N7877,N7881,N7882);
and and4697(N7878,N7883,in1);
and and4698(N7879,in2,R0);
and and4699(N7880,R1,R2);
and and4705(N7889,N7893,N7894);
and and4706(N7890,N7895,in1);
and and4707(N7891,R0,R1);
and and4708(N7892,R2,N7896);
and and4714(N7901,N7905,N7906);
and and4715(N7902,N7907,N7908);
and and4716(N7903,in2,R0);
and and4717(N7904,R1,R2);
and and4723(N7913,N7917,N7918);
and and4724(N7914,N7919,in1);
and and4725(N7915,N7920,R0);
and and4726(N7916,R1,R2);
and and4732(N7925,N7929,N7930);
and and4733(N7926,N7931,in1);
and and4734(N7927,in2,R1);
and and4735(N7928,R2,R3);
and and4741(N7937,N7941,N7942);
and and4742(N7938,N7943,in1);
and and4743(N7939,N7944,R0);
and and4744(N7940,R1,R2);
and and4750(N7949,N7953,N7954);
and and4751(N7950,N7955,in1);
and and4752(N7951,N7956,R0);
and and4753(N7952,R1,R2);
and and4759(N7961,N7965,N7966);
and and4760(N7962,N7967,in2);
and and4761(N7963,R0,R1);
and and4762(N7964,R2,N7968);
and and4768(N7973,N7977,N7978);
and and4769(N7974,N7979,in1);
and and4770(N7975,in2,R0);
and and4771(N7976,N7980,R2);
and and4777(N7984,N7988,N7989);
and and4778(N7985,N7990,in1);
and and4779(N7986,in2,R0);
and and4780(N7987,N7991,R2);
and and4786(N7995,N7999,N8000);
and and4787(N7996,N8001,in1);
and and4788(N7997,in2,R0);
and and4789(N7998,N8002,R2);
and and4795(N8006,N8010,N8011);
and and4796(N8007,N8012,in1);
and and4797(N8008,in2,R0);
and and4798(N8009,N8013,R3);
and and4804(N8017,N8021,N8022);
and and4805(N8018,N8023,in1);
and and4806(N8019,in2,N8024);
and and4807(N8020,R2,R3);
and and4813(N8028,N8032,N8033);
and and4814(N8029,N8034,in1);
and and4815(N8030,in2,N8035);
and and4816(N8031,R1,R2);
and and4822(N8039,N8043,N8044);
and and4823(N8040,N8045,in1);
and and4824(N8041,in2,R0);
and and4825(N8042,N8046,R2);
and and4831(N8050,N8054,N8055);
and and4832(N8051,N8056,in1);
and and4833(N8052,R0,R1);
and and4834(N8053,N8057,R3);
and and4840(N8061,N8065,N8066);
and and4841(N8062,N8067,in2);
and and4842(N8063,R0,R1);
and and4843(N8064,R2,R3);
and and4849(N8071,N8075,N8076);
and and4850(N8072,N8077,R0);
and and4851(N8073,N8078,N8079);
and and4852(N8074,N8080,N8081);
and and4857(N8087,N8091,N8092);
and and4858(N8088,N8093,N8094);
and and4859(N8089,N8095,R3);
and and4860(N8090,N8096,N8097);
and and4865(N8103,N8107,N8108);
and and4866(N8104,N8109,N8110);
and and4867(N8105,N8111,N8112);
and and4868(N8106,N8113,N8114);
and and4873(N8119,N8123,N8124);
and and4874(N8120,N8125,N8126);
and and4875(N8121,N8127,N8128);
and and4876(N8122,N8129,N8130);
and and4881(N8135,N8139,N8140);
and and4882(N8136,N8141,N8142);
and and4883(N8137,R0,R1);
and and4884(N8138,N8143,N8144);
and and4889(N8150,N8154,N8155);
and and4890(N8151,N8156,N8157);
and and4891(N8152,N8158,N8159);
and and4892(N8153,R4,R5);
and and4897(N8165,N8169,N8170);
and and4898(N8166,in2,N8171);
and and4899(N8167,N8172,R3);
and and4900(N8168,N8173,N8174);
and and4905(N8180,N8184,N8185);
and and4906(N8181,in2,N8186);
and and4907(N8182,N8187,R3);
and and4908(N8183,N8188,N8189);
and and4913(N8195,N8199,N8200);
and and4914(N8196,in1,N8201);
and and4915(N8197,N8202,R1);
and and4916(N8198,R3,N8203);
and and4921(N8209,N8213,N8214);
and and4922(N8210,N8215,in2);
and and4923(N8211,N8216,R1);
and and4924(N8212,R2,N8217);
and and4929(N8223,N8227,N8228);
and and4930(N8224,N8229,N8230);
and and4931(N8225,R0,N8231);
and and4932(N8226,R2,N8232);
and and4937(N8237,N8241,N8242);
and and4938(N8238,N8243,N8244);
and and4939(N8239,N8245,N8246);
and and4940(N8240,R2,R4);
and and4945(N8251,N8255,N8256);
and and4946(N8252,in1,N8257);
and and4947(N8253,N8258,R1);
and and4948(N8254,R3,N8259);
and and4953(N8265,N8269,N8270);
and and4954(N8266,in1,N8271);
and and4955(N8267,N8272,R3);
and and4956(N8268,R4,R5);
and and4961(N8278,N8282,N8283);
and and4962(N8279,in1,N8284);
and and4963(N8280,R0,N8285);
and and4964(N8281,N8286,N8287);
and and4969(N8291,N8295,N8296);
and and4970(N8292,in1,in2);
and and4971(N8293,R0,N8297);
and and4972(N8294,N8298,R5);
and and4977(N8304,N8308,N8309);
and and4978(N8305,in1,N8310);
and and4979(N8306,R0,N8311);
and and4980(N8307,R3,N8312);
and and4985(N8317,N8321,N8322);
and and4986(N8318,in1,in2);
and and4987(N8319,N8323,R3);
and and4988(N8320,R4,N8324);
and and4993(N8330,N8334,N8335);
and and4994(N8331,N8336,N8337);
and and4995(N8332,N8338,R2);
and and4996(N8333,R3,N8339);
and and5001(N8343,N8347,N8348);
and and5002(N8344,in1,in2);
and and5003(N8345,R0,N8349);
and and5004(N8346,N8350,R5);
and and5009(N8356,N8360,N8361);
and and5010(N8357,N8362,in2);
and and5011(N8358,N8363,R1);
and and5012(N8359,R2,R3);
and and5017(N8368,N8372,N8373);
and and5018(N8369,N8374,in2);
and and5019(N8370,R0,R1);
and and5020(N8371,N8375,R4);
and and5025(N8380,N8384,N8385);
and and5026(N8381,in2,R0);
and and5027(N8382,N8386,N8387);
and and5028(N8383,R3,N8388);
and and5033(N8392,N8396,N8397);
and and5034(N8393,in1,N8398);
and and5035(N8394,N8399,N8400);
and and5036(N8395,R3,R4);
and and5041(N8404,N8408,N8409);
and and5042(N8405,in1,N8410);
and and5043(N8406,N8411,R2);
and and5044(N8407,N8412,R5);
and and5049(N8416,N8420,N8421);
and and5050(N8417,in1,R0);
and and5051(N8418,N8422,N8423);
and and5052(N8419,R3,R4);
and and3429(N5851,R2,N5857);
and and3430(N5852,N5858,N5859);
and and3431(N5853,R6,R7);
and and3439(N5867,R2,N5872);
and and3440(N5868,R4,N5873);
and and3441(N5869,R6,N5874);
and and3449(N5882,N5888,N5889);
and and3450(N5883,N5890,N5891);
and and3458(N5899,R4,N5906);
and and3459(N5900,N5907,N5908);
and and3467(N5916,N5922,N5923);
and and3468(N5917,N5924,N5925);
and and3476(N5933,N5939,N5940);
and and3477(N5934,N5941,N5942);
and and3485(N5950,N5956,N5957);
and and3486(N5951,N5958,N5959);
and and3494(N5967,N5974,R5);
and and3495(N5968,N5975,N5976);
and and3503(N5984,N5991,R5);
and and3504(N5985,N5992,N5993);
and and3512(N6001,N6008,N6009);
and and3513(N6002,R5,N6010);
and and3521(N6018,N6025,R5);
and and3522(N6019,N6026,N6027);
and and3530(N6035,N6042,N6043);
and and3531(N6036,N6044,R7);
and and3539(N6052,R4,N6059);
and and3540(N6053,N6060,N6061);
and and3548(N6069,N6075,N6076);
and and3549(N6070,R6,N6077);
and and3557(N6085,R4,N6091);
and and3558(N6086,N6092,N6093);
and and3566(N6101,R4,N6107);
and and3567(N6102,N6108,N6109);
and and3575(N6117,N6122,N6123);
and and3576(N6118,N6124,N6125);
and and3584(N6133,N6139,N6140);
and and3585(N6134,R6,N6141);
and and3593(N6149,R3,N6155);
and and3594(N6150,N6156,N6157);
and and3602(N6165,R4,N6171);
and and3603(N6166,N6172,N6173);
and and3611(N6181,N6187,N6188);
and and3612(N6182,N6189,R6);
and and3620(N6197,R4,N6204);
and and3621(N6198,R6,N6205);
and and3629(N6213,N6219,N6220);
and and3630(N6214,R6,N6221);
and and3638(N6229,R3,N6236);
and and3639(N6230,N6237,R6);
and and3647(N6245,R3,N6251);
and and3648(N6246,N6252,N6253);
and and3656(N6261,R3,N6267);
and and3657(N6262,N6268,N6269);
and and3665(N6277,R3,R4);
and and3666(N6278,N6284,N6285);
and and3674(N6293,N6299,R5);
and and3675(N6294,N6300,R7);
and and3683(N6308,R4,R5);
and and3684(N6309,N6315,R7);
and and3692(N6323,N6328,N6329);
and and3693(N6324,N6330,R7);
and and3701(N6338,R4,R5);
and and3702(N6339,N6344,N6345);
and and3710(N6353,R4,N6358);
and and3711(N6354,N6359,N6360);
and and3719(N6368,N6373,N6374);
and and3720(N6369,N6375,R7);
and and3728(N6383,N6388,N6389);
and and3729(N6384,R6,N6390);
and and3737(N6398,N6403,R5);
and and3738(N6399,N6404,N6405);
and and3746(N6413,N6418,N6419);
and and3747(N6414,N6420,R7);
and and3755(N6428,N6435,R5);
and and3756(N6429,R6,R7);
and and3764(N6443,N6449,R5);
and and3765(N6444,R6,N6450);
and and3773(N6458,N6464,R5);
and and3774(N6459,R6,N6465);
and and3782(N6473,N6479,R5);
and and3783(N6474,N6480,R7);
and and3791(N6488,N6494,R5);
and and3792(N6489,R6,N6495);
and and3800(N6503,N6508,N6509);
and and3801(N6504,N6510,R7);
and and3809(N6518,N6523,N6524);
and and3810(N6519,N6525,R7);
and and3818(N6533,N6538,N6539);
and and3819(N6534,N6540,R7);
and and3827(N6548,N6554,R5);
and and3828(N6549,N6555,R7);
and and3836(N6563,N6568,R5);
and and3837(N6564,N6569,N6570);
and and3845(N6578,N6584,R4);
and and3846(N6579,R5,N6585);
and and3854(N6593,R4,N6599);
and and3855(N6594,N6600,R7);
and and3863(N6608,N6614,R5);
and and3864(N6609,N6615,R7);
and and3872(N6623,N6630,R5);
and and3873(N6624,R6,R7);
and and3881(N6638,N6644,R5);
and and3882(N6639,R6,N6645);
and and3890(N6653,N6659,N6660);
and and3891(N6654,R6,R7);
and and3899(N6668,N6673,R5);
and and3900(N6669,N6674,N6675);
and and3908(N6683,N6688,N6689);
and and3909(N6684,N6690,R7);
and and3917(N6698,R3,R4);
and and3918(N6699,N6704,N6705);
and and3926(N6713,R3,R4);
and and3927(N6714,N6719,N6720);
and and3935(N6728,R3,N6734);
and and3936(N6729,R5,N6735);
and and3944(N6743,R3,R4);
and and3945(N6744,N6749,N6750);
and and3953(N6758,R4,N6764);
and and3954(N6759,R6,N6765);
and and3962(N6773,N6779,R4);
and and3963(N6774,R5,N6780);
and and3971(N6788,N6793,R5);
and and3972(N6789,N6794,N6795);
and and3980(N6803,N6808,N6809);
and and3981(N6804,N6810,R7);
and and3989(N6818,R4,N6824);
and and3990(N6819,R6,N6825);
and and3998(N6833,R4,R5);
and and3999(N6834,N6840,R7);
and and4007(N6848,R3,N6854);
and and4008(N6849,R6,N6855);
and and4016(N6863,R3,R5);
and and4017(N6864,N6869,N6870);
and and4025(N6878,N6884,R4);
and and4026(N6879,N6885,R7);
and and4034(N6893,N6899,R5);
and and4035(N6894,R6,N6900);
and and4043(N6908,N6914,R4);
and and4044(N6909,N6915,R7);
and and4052(N6923,N6927,N6928);
and and4053(N6924,N6929,N6930);
and and4061(N6938,N6943,R5);
and and4062(N6939,N6944,N6945);
and and4070(N6953,R4,R5);
and and4071(N6954,N6959,R7);
and and4079(N6967,N6970,N6971);
and and4080(N6968,N6972,N6973);
and and4088(N6981,R3,N6985);
and and4089(N6982,N6986,N6987);
and and4097(N6995,N6999,N7000);
and and4098(N6996,R6,N7001);
and and4106(N7009,N7013,N7014);
and and4107(N7010,R6,N7015);
and and4115(N7023,R4,R5);
and and4116(N7024,R6,R7);
and and4124(N7037,N7042,R4);
and and4125(N7038,N7043,R7);
and and4133(N7051,R3,N7056);
and and4134(N7052,R6,N7057);
and and4142(N7065,R4,R5);
and and4143(N7066,R6,N7071);
and and4151(N7079,N7084,N7085);
and and4152(N7080,R5,R6);
and and4160(N7093,R4,N7098);
and and4161(N7094,R6,N7099);
and and4169(N7107,N7111,R4);
and and4170(N7108,N7112,N7113);
and and4178(N7121,N7125,R5);
and and4179(N7122,N7126,N7127);
and and4187(N7135,N7139,R4);
and and4188(N7136,N7140,N7141);
and and4196(N7149,R3,N7155);
and and4197(N7150,R6,R7);
and and4205(N7163,R3,N7169);
and and4206(N7164,R6,R7);
and and4214(N7177,N7181,N7182);
and and4215(N7178,R6,N7183);
and and4223(N7191,R3,N7196);
and and4224(N7192,N7197,R7);
and and4232(N7205,R3,R4);
and and4233(N7206,R5,R7);
and and4241(N7219,R4,R5);
and and4242(N7220,N7224,N7225);
and and4250(N7233,N7238,R5);
and and4251(N7234,R6,N7239);
and and4259(N7247,N7251,N7252);
and and4260(N7248,N7253,R7);
and and4268(N7261,N7265,N7266);
and and4269(N7262,N7267,R7);
and and4277(N7275,R4,R5);
and and4278(N7276,N7279,N7280);
and and4286(N7288,R4,R5);
and and4287(N7289,R6,N7293);
and and4295(N7301,R4,R5);
and and4296(N7302,R6,R7);
and and4304(N7314,R3,R5);
and and4305(N7315,N7319,R7);
and and4313(N7327,N7331,R5);
and and4314(N7328,R6,N7332);
and and4322(N7340,N7344,R4);
and and4323(N7341,R5,N7345);
and and4331(N7353,R3,R4);
and and4332(N7354,N7357,N7358);
and and4340(N7366,R3,R4);
and and4341(N7367,N7371,R7);
and and4349(N7379,N7384,R4);
and and4350(N7380,R6,R7);
and and4358(N7392,N7396,R5);
and and4359(N7393,N7397,R7);
and and4367(N7405,N7409,R5);
and and4368(N7406,N7410,R7);
and and4376(N7418,N7422,R5);
and and4377(N7419,N7423,R7);
and and4385(N7431,R3,R5);
and and4386(N7432,R6,R7);
and and4394(N7444,R3,R4);
and and4395(N7445,N7449,R6);
and and4403(N7457,N7462,R4);
and and4404(N7458,R5,R6);
and and4412(N7470,N7475,R5);
and and4413(N7471,R6,R7);
and and4421(N7483,R4,N7487);
and and4422(N7484,R6,N7488);
and and4430(N7496,R4,N7500);
and and4431(N7497,R6,N7501);
and and4439(N7509,N7514,R5);
and and4440(N7510,R6,R7);
and and4448(N7522,N7526,R5);
and and4449(N7523,R6,N7527);
and and4457(N7535,R4,R5);
and and4458(N7536,R6,R7);
and and4466(N7548,R4,R5);
and and4467(N7549,R6,R7);
and and4475(N7561,N7564,N7565);
and and4476(N7562,N7566,R7);
and and4484(N7574,R3,R4);
and and4485(N7575,N7579,R7);
and and4493(N7587,R3,R4);
and and4494(N7588,R5,N7592);
and and4502(N7600,R4,R5);
and and4503(N7601,N7604,N7605);
and and4511(N7613,R4,N7616);
and and4512(N7614,N7617,N7618);
and and4520(N7626,R4,R5);
and and4521(N7627,N7631,R7);
and and4529(N7639,R3,R4);
and and4530(N7640,R5,R7);
and and4538(N7652,R4,R5);
and and4539(N7653,R6,N7657);
and and4547(N7665,N7670,R5);
and and4548(N7666,R6,R7);
and and4556(N7678,R4,R5);
and and4557(N7679,N7683,R7);
and and4565(N7691,N7696,R4);
and and4566(N7692,R5,R7);
and and4574(N7704,R4,N7708);
and and4575(N7705,N7709,R7);
and and4583(N7717,R4,R5);
and and4584(N7718,N7722,R7);
and and4592(N7730,N7735,R5);
and and4593(N7731,R6,R7);
and and4601(N7743,R4,R5);
and and4602(N7744,R6,N7748);
and and4610(N7756,R4,R5);
and and4611(N7757,N7761,R7);
and and4619(N7769,N7773,R5);
and and4620(N7770,R6,N7774);
and and4628(N7782,R4,R5);
and and4629(N7783,R6,N7787);
and and4637(N7795,N7799,R5);
and and4638(N7796,N7800,R7);
and and4646(N7808,N7813,R5);
and and4647(N7809,R6,R7);
and and4655(N7821,R4,R5);
and and4656(N7822,R6,R7);
and and4664(N7833,N7836,N7837);
and and4665(N7834,R6,R7);
and and4673(N7845,R4,N7849);
and and4674(N7846,R6,R7);
and and4682(N7857,R4,R5);
and and4683(N7858,R6,N7861);
and and4691(N7869,N7873,R5);
and and4692(N7870,R6,R7);
and and4700(N7881,R3,N7884);
and and4701(N7882,R6,N7885);
and and4709(N7893,R4,N7897);
and and4710(N7894,R6,R7);
and and4718(N7905,R3,N7909);
and and4719(N7906,R6,R7);
and and4727(N7917,R3,R4);
and and4728(N7918,R5,N7921);
and and4736(N7929,R4,N7932);
and and4737(N7930,N7933,R7);
and and4745(N7941,R3,R4);
and and4746(N7942,R5,N7945);
and and4754(N7953,R4,N7957);
and and4755(N7954,R6,R7);
and and4763(N7965,R4,R5);
and and4764(N7966,N7969,R7);
and and4772(N7977,R4,R5);
and and4773(N7978,R6,R7);
and and4781(N7988,R3,R4);
and and4782(N7989,R5,R6);
and and4790(N7999,R3,R4);
and and4791(N8000,R5,R7);
and and4799(N8010,R4,R5);
and and4800(N8011,R6,R7);
and and4808(N8021,R4,R5);
and and4809(N8022,R6,R7);
and and4817(N8032,R3,R4);
and and4818(N8033,R5,R7);
and and4826(N8043,R3,R5);
and and4827(N8044,R6,R7);
and and4835(N8054,R4,R5);
and and4836(N8055,R6,R7);
and and4844(N8065,R4,R5);
and and4845(N8066,R6,R7);
and and4853(N8075,N8082,N8083);
and and4861(N8091,N8098,N8099);
and and4869(N8107,N8115,R7);
and and4877(N8123,N8131,R7);
and and4885(N8139,N8145,N8146);
and and4893(N8154,N8160,N8161);
and and4901(N8169,N8175,N8176);
and and4909(N8184,N8190,N8191);
and and4917(N8199,N8204,N8205);
and and4925(N8213,N8218,N8219);
and and4933(N8227,N8233,R7);
and and4941(N8241,N8247,R6);
and and4949(N8255,N8260,N8261);
and and4957(N8269,N8273,N8274);
and and4965(N8282,R5,R7);
and and4973(N8295,N8299,N8300);
and and4981(N8308,N8313,R7);
and and4989(N8321,N8325,N8326);
and and4997(N8334,R6,R7);
and and5005(N8347,N8351,N8352);
and and5013(N8360,R6,N8364);
and and5021(N8372,N8376,R7);
and and5029(N8384,R6,R7);
and and5037(N8396,R5,R6);
and and5045(N8408,R6,R7);
and and5053(N8420,R5,N8424);
and and5054(N8885,N8886,N8887);
and and5063(N8903,N8904,N8905);
and and5072(N8920,N8921,N8922);
and and5081(N8937,N8938,N8939);
and and5090(N8954,N8955,N8956);
and and5099(N8971,N8972,N8973);
and and5108(N8988,N8989,N8990);
and and5117(N9004,N9005,N9006);
and and5126(N9020,N9021,N9022);
and and5135(N9036,N9037,N9038);
and and5144(N9052,N9053,N9054);
and and5153(N9068,N9069,N9070);
and and5162(N9084,N9085,N9086);
and and5171(N9100,N9101,N9102);
and and5180(N9116,N9117,N9118);
and and5189(N9132,N9133,N9134);
and and5198(N9148,N9149,N9150);
and and5207(N9164,N9165,N9166);
and and5216(N9180,N9181,N9182);
and and5225(N9196,N9197,N9198);
and and5234(N9212,N9213,N9214);
and and5243(N9228,N9229,N9230);
and and5252(N9243,N9244,N9245);
and and5261(N9258,N9259,N9260);
and and5270(N9273,N9274,N9275);
and and5279(N9288,N9289,N9290);
and and5288(N9303,N9304,N9305);
and and5297(N9318,N9319,N9320);
and and5306(N9333,N9334,N9335);
and and5315(N9348,N9349,N9350);
and and5324(N9363,N9364,N9365);
and and5333(N9378,N9379,N9380);
and and5342(N9393,N9394,N9395);
and and5351(N9408,N9409,N9410);
and and5360(N9423,N9424,N9425);
and and5369(N9438,N9439,N9440);
and and5378(N9453,N9454,N9455);
and and5387(N9468,N9469,N9470);
and and5396(N9483,N9484,N9485);
and and5405(N9498,N9499,N9500);
and and5414(N9513,N9514,N9515);
and and5423(N9528,N9529,N9530);
and and5432(N9543,N9544,N9545);
and and5441(N9558,N9559,N9560);
and and5450(N9573,N9574,N9575);
and and5459(N9588,N9589,N9590);
and and5468(N9603,N9604,N9605);
and and5477(N9618,N9619,N9620);
and and5486(N9633,N9634,N9635);
and and5495(N9648,N9649,N9650);
and and5504(N9663,N9664,N9665);
and and5513(N9678,N9679,N9680);
and and5522(N9693,N9694,N9695);
and and5531(N9708,N9709,N9710);
and and5540(N9723,N9724,N9725);
and and5549(N9738,N9739,N9740);
and and5558(N9752,N9753,N9754);
and and5567(N9766,N9767,N9768);
and and5576(N9780,N9781,N9782);
and and5585(N9794,N9795,N9796);
and and5594(N9808,N9809,N9810);
and and5603(N9822,N9823,N9824);
and and5612(N9836,N9837,N9838);
and and5621(N9850,N9851,N9852);
and and5630(N9864,N9865,N9866);
and and5639(N9878,N9879,N9880);
and and5648(N9892,N9893,N9894);
and and5657(N9906,N9907,N9908);
and and5666(N9920,N9921,N9922);
and and5675(N9934,N9935,N9936);
and and5684(N9948,N9949,N9950);
and and5693(N9962,N9963,N9964);
and and5702(N9976,N9977,N9978);
and and5711(N9990,N9991,N9992);
and and5720(N10004,N10005,N10006);
and and5729(N10018,N10019,N10020);
and and5738(N10032,N10033,N10034);
and and5747(N10046,N10047,N10048);
and and5756(N10060,N10061,N10062);
and and5765(N10074,N10075,N10076);
and and5774(N10088,N10089,N10090);
and and5783(N10102,N10103,N10104);
and and5792(N10116,N10117,N10118);
and and5801(N10130,N10131,N10132);
and and5810(N10144,N10145,N10146);
and and5819(N10158,N10159,N10160);
and and5828(N10172,N10173,N10174);
and and5837(N10186,N10187,N10188);
and and5846(N10200,N10201,N10202);
and and5855(N10214,N10215,N10216);
and and5864(N10228,N10229,N10230);
and and5873(N10242,N10243,N10244);
and and5882(N10256,N10257,N10258);
and and5891(N10270,N10271,N10272);
and and5900(N10284,N10285,N10286);
and and5909(N10298,N10299,N10300);
and and5918(N10311,N10312,N10313);
and and5927(N10324,N10325,N10326);
and and5936(N10337,N10338,N10339);
and and5945(N10350,N10351,N10352);
and and5954(N10363,N10364,N10365);
and and5963(N10376,N10377,N10378);
and and5972(N10389,N10390,N10391);
and and5981(N10402,N10403,N10404);
and and5990(N10415,N10416,N10417);
and and5999(N10428,N10429,N10430);
and and6008(N10441,N10442,N10443);
and and6017(N10454,N10455,N10456);
and and6026(N10467,N10468,N10469);
and and6035(N10480,N10481,N10482);
and and6044(N10493,N10494,N10495);
and and6053(N10506,N10507,N10508);
and and6062(N10519,N10520,N10521);
and and6071(N10532,N10533,N10534);
and and6080(N10545,N10546,N10547);
and and6089(N10558,N10559,N10560);
and and6098(N10571,N10572,N10573);
and and6107(N10584,N10585,N10586);
and and6116(N10597,N10598,N10599);
and and6125(N10610,N10611,N10612);
and and6134(N10623,N10624,N10625);
and and6143(N10636,N10637,N10638);
and and6152(N10649,N10650,N10651);
and and6161(N10662,N10663,N10664);
and and6170(N10675,N10676,N10677);
and and6179(N10688,N10689,N10690);
and and6188(N10701,N10702,N10703);
and and6197(N10714,N10715,N10716);
and and6206(N10727,N10728,N10729);
and and6215(N10740,N10741,N10742);
and and6224(N10753,N10754,N10755);
and and6233(N10766,N10767,N10768);
and and6242(N10779,N10780,N10781);
and and6251(N10792,N10793,N10794);
and and6260(N10805,N10806,N10807);
and and6269(N10818,N10819,N10820);
and and6278(N10830,N10831,N10832);
and and6287(N10842,N10843,N10844);
and and6296(N10854,N10855,N10856);
and and6305(N10866,N10867,N10868);
and and6314(N10878,N10879,N10880);
and and6323(N10890,N10891,N10892);
and and6332(N10902,N10903,N10904);
and and6341(N10914,N10915,N10916);
and and6350(N10926,N10927,N10928);
and and6359(N10938,N10939,N10940);
and and6368(N10950,N10951,N10952);
and and6377(N10962,N10963,N10964);
and and6386(N10974,N10975,N10976);
and and6395(N10986,N10987,N10988);
and and6404(N10998,N10999,N11000);
and and6413(N11010,N11011,N11012);
and and6422(N11022,N11023,N11024);
and and6431(N11034,N11035,N11036);
and and6440(N11046,N11047,N11048);
and and6449(N11058,N11059,N11060);
and and6458(N11070,N11071,N11072);
and and6467(N11082,N11083,N11084);
and and6476(N11094,N11095,N11096);
and and6485(N11106,N11107,N11108);
and and6494(N11118,N11119,N11120);
and and6503(N11130,N11131,N11132);
and and6512(N11142,N11143,N11144);
and and6521(N11153,N11154,N11155);
and and6530(N11164,N11165,N11166);
and and6539(N11175,N11176,N11177);
and and6548(N11186,N11187,N11188);
and and6557(N11197,N11198,N11199);
and and6566(N11208,N11209,N11210);
and and6575(N11219,N11220,N11221);
and and6584(N11230,N11231,N11232);
and and6593(N11241,N11242,N11243);
and and6602(N11252,N11253,N11254);
and and6611(N11263,N11264,N11265);
and and6620(N11274,N11275,N11276);
and and6629(N11285,N11286,N11287);
and and6638(N11296,N11297,N11298);
and and6647(N11307,N11308,N11309);
and and6656(N11318,N11319,N11320);
and and6665(N11328,N11329,N11330);
and and6674(N11338,N11339,N11340);
and and6683(N11348,N11349,N11350);
and and6692(N11358,N11359,N11360);
and and6701(N11368,N11369,N11370);
and and6709(N11384,N11385,N11386);
and and6717(N11400,N11401,N11402);
and and6725(N11416,N11417,N11418);
and and6733(N11432,N11433,N11434);
and and6741(N11448,N11449,N11450);
and and6749(N11464,N11465,N11466);
and and6757(N11480,N11481,N11482);
and and6765(N11495,N11496,N11497);
and and6773(N11510,N11511,N11512);
and and6781(N11525,N11526,N11527);
and and6789(N11540,N11541,N11542);
and and6797(N11555,N11556,N11557);
and and6805(N11570,N11571,N11572);
and and6813(N11585,N11586,N11587);
and and6821(N11599,N11600,N11601);
and and6829(N11613,N11614,N11615);
and and6837(N11627,N11628,N11629);
and and6845(N11641,N11642,N11643);
and and6853(N11655,N11656,N11657);
and and6861(N11669,N11670,N11671);
and and6869(N11683,N11684,N11685);
and and6877(N11697,N11698,N11699);
and and6885(N11711,N11712,N11713);
and and6893(N11725,N11726,N11727);
and and6901(N11739,N11740,N11741);
and and6909(N11753,N11754,N11755);
and and6917(N11767,N11768,N11769);
and and6925(N11781,N11782,N11783);
and and6933(N11795,N11796,N11797);
and and6941(N11809,N11810,N11811);
and and6949(N11823,N11824,N11825);
and and6957(N11837,N11838,N11839);
and and6965(N11851,N11852,N11853);
and and6973(N11865,N11866,N11867);
and and6981(N11879,N11880,N11881);
and and6989(N11893,N11894,N11895);
and and6997(N11907,N11908,N11909);
and and7005(N11921,N11922,N11923);
and and7013(N11935,N11936,N11937);
and and7021(N11949,N11950,N11951);
and and7029(N11963,N11964,N11965);
and and7037(N11977,N11978,N11979);
and and7045(N11991,N11992,N11993);
and and7053(N12005,N12006,N12007);
and and7061(N12019,N12020,N12021);
and and7069(N12033,N12034,N12035);
and and7077(N12047,N12048,N12049);
and and7085(N12061,N12062,N12063);
and and7093(N12075,N12076,N12077);
and and7101(N12088,N12089,N12090);
and and7109(N12101,N12102,N12103);
and and7117(N12114,N12115,N12116);
and and7125(N12127,N12128,N12129);
and and7133(N12140,N12141,N12142);
and and7141(N12153,N12154,N12155);
and and7149(N12166,N12167,N12168);
and and7157(N12179,N12180,N12181);
and and7165(N12192,N12193,N12194);
and and7173(N12205,N12206,N12207);
and and7181(N12218,N12219,N12220);
and and7189(N12231,N12232,N12233);
and and7197(N12244,N12245,N12246);
and and7205(N12257,N12258,N12259);
and and7213(N12270,N12271,N12272);
and and7221(N12283,N12284,N12285);
and and7229(N12296,N12297,N12298);
and and7237(N12309,N12310,N12311);
and and7245(N12322,N12323,N12324);
and and7253(N12335,N12336,N12337);
and and7261(N12348,N12349,N12350);
and and7269(N12361,N12362,N12363);
and and7277(N12374,N12375,N12376);
and and7285(N12387,N12388,N12389);
and and7293(N12400,N12401,N12402);
and and7301(N12413,N12414,N12415);
and and7309(N12426,N12427,N12428);
and and7317(N12439,N12440,N12441);
and and7325(N12452,N12453,N12454);
and and7333(N12465,N12466,N12467);
and and7341(N12478,N12479,N12480);
and and7349(N12491,N12492,N12493);
and and7357(N12504,N12505,N12506);
and and7365(N12517,N12518,N12519);
and and7373(N12530,N12531,N12532);
and and7381(N12543,N12544,N12545);
and and7389(N12556,N12557,N12558);
and and7397(N12569,N12570,N12571);
and and7405(N12582,N12583,N12584);
and and7413(N12595,N12596,N12597);
and and7421(N12608,N12609,N12610);
and and7429(N12621,N12622,N12623);
and and7437(N12634,N12635,N12636);
and and7445(N12647,N12648,N12649);
and and7453(N12660,N12661,N12662);
and and7461(N12673,N12674,N12675);
and and7469(N12685,N12686,N12687);
and and7477(N12697,N12698,N12699);
and and7485(N12709,N12710,N12711);
and and7493(N12721,N12722,N12723);
and and7501(N12733,N12734,N12735);
and and7509(N12745,N12746,N12747);
and and7517(N12757,N12758,N12759);
and and7525(N12769,N12770,N12771);
and and7533(N12781,N12782,N12783);
and and7541(N12793,N12794,N12795);
and and7549(N12805,N12806,N12807);
and and7557(N12817,N12818,N12819);
and and7565(N12829,N12830,N12831);
and and7573(N12841,N12842,N12843);
and and7581(N12853,N12854,N12855);
and and7589(N12865,N12866,N12867);
and and7597(N12877,N12878,N12879);
and and7605(N12889,N12890,N12891);
and and7613(N12901,N12902,N12903);
and and7621(N12913,N12914,N12915);
and and7629(N12925,N12926,N12927);
and and7637(N12937,N12938,N12939);
and and7645(N12949,N12950,N12951);
and and7653(N12961,N12962,N12963);
and and7661(N12973,N12974,N12975);
and and7669(N12985,N12986,N12987);
and and7677(N12997,N12998,N12999);
and and7685(N13009,N13010,N13011);
and and7693(N13021,N13022,N13023);
and and7701(N13033,N13034,N13035);
and and7709(N13045,N13046,N13047);
and and7717(N13057,N13058,N13059);
and and7725(N13069,N13070,N13071);
and and7733(N13081,N13082,N13083);
and and7741(N13093,N13094,N13095);
and and7749(N13105,N13106,N13107);
and and7757(N13117,N13118,N13119);
and and7765(N13129,N13130,N13131);
and and7773(N13141,N13142,N13143);
and and7781(N13153,N13154,N13155);
and and7789(N13165,N13166,N13167);
and and7797(N13177,N13178,N13179);
and and7805(N13189,N13190,N13191);
and and7813(N13201,N13202,N13203);
and and7821(N13213,N13214,N13215);
and and7829(N13225,N13226,N13227);
and and7837(N13237,N13238,N13239);
and and7845(N13249,N13250,N13251);
and and7853(N13261,N13262,N13263);
and and7861(N13273,N13274,N13275);
and and7869(N13285,N13286,N13287);
and and7877(N13297,N13298,N13299);
and and7885(N13309,N13310,N13311);
and and7893(N13321,N13322,N13323);
and and7901(N13333,N13334,N13335);
and and7909(N13345,N13346,N13347);
and and7917(N13357,N13358,N13359);
and and7925(N13369,N13370,N13371);
and and7933(N13381,N13382,N13383);
and and7941(N13393,N13394,N13395);
and and7949(N13404,N13405,N13406);
and and7957(N13415,N13416,N13417);
and and7965(N13426,N13427,N13428);
and and7973(N13437,N13438,N13439);
and and7981(N13448,N13449,N13450);
and and7989(N13459,N13460,N13461);
and and7997(N13470,N13471,N13472);
and and8005(N13481,N13482,N13483);
and and8013(N13492,N13493,N13494);
and and8021(N13503,N13504,N13505);
and and8029(N13514,N13515,N13516);
and and8037(N13525,N13526,N13527);
and and8045(N13536,N13537,N13538);
and and8053(N13547,N13548,N13549);
and and8061(N13558,N13559,N13560);
and and8069(N13569,N13570,N13571);
and and8077(N13580,N13581,N13582);
and and8085(N13591,N13592,N13593);
and and8093(N13602,N13603,N13604);
and and8101(N13613,N13614,N13615);
and and8109(N13624,N13625,N13626);
and and8117(N13635,N13636,N13637);
and and8125(N13646,N13647,N13648);
and and8133(N13657,N13658,N13659);
and and8141(N13668,N13669,N13670);
and and8149(N13679,N13680,N13681);
and and8157(N13690,N13691,N13692);
and and8165(N13701,N13702,N13703);
and and8173(N13712,N13713,N13714);
and and8181(N13723,N13724,N13725);
and and8189(N13734,N13735,N13736);
and and8197(N13745,N13746,N13747);
and and8205(N13756,N13757,N13758);
and and8213(N13767,N13768,N13769);
and and8221(N13778,N13779,N13780);
and and8229(N13789,N13790,N13791);
and and8237(N13800,N13801,N13802);
and and8245(N13811,N13812,N13813);
and and8253(N13822,N13823,N13824);
and and8261(N13833,N13834,N13835);
and and8269(N13844,N13845,N13846);
and and8277(N13855,N13856,N13857);
and and8285(N13866,N13867,N13868);
and and8293(N13877,N13878,N13879);
and and8301(N13888,N13889,N13890);
and and8309(N13899,N13900,N13901);
and and8317(N13910,N13911,N13912);
and and8325(N13921,N13922,N13923);
and and8333(N13932,N13933,N13934);
and and8341(N13943,N13944,N13945);
and and8349(N13954,N13955,N13956);
and and8357(N13964,N13965,N13966);
and and8365(N13974,N13975,N13976);
and and8373(N13984,N13985,N13986);
and and8381(N13994,N13995,N13996);
and and8389(N14004,N14005,N14006);
and and8397(N14014,N14015,N14016);
and and8405(N14024,N14025,N14026);
and and8413(N14034,N14035,N14036);
and and8421(N14044,N14045,N14046);
and and8429(N14054,N14055,N14056);
and and8437(N14064,N14065,N14066);
and and8445(N14074,N14075,N14076);
and and8453(N14084,N14085,N14086);
and and8461(N14094,N14095,N14096);
and and8469(N14104,N14105,N14106);
and and8477(N14114,N14115,N14116);
and and8485(N14123,N14124,N14125);
and and8493(N14132,N14133,N14134);
and and8501(N14141,N14142,N14143);
and and8509(N14150,N14151,N14152);
and and8517(N14159,N14160,N14161);
and and8525(N14168,N14169,N14170);
and and8533(N14177,N14178,N14179);
and and8541(N14186,N14187,N14188);
and and8549(N14195,N14196,N14197);
and and8557(N14204,N14205,N14206);
and and8564(N14218,N14219,N14220);
and and8571(N14232,N14233,N14234);
and and8578(N14246,N14247,N14248);
and and8585(N14260,N14261,N14262);
and and8592(N14273,N14274,N14275);
and and8599(N14286,N14287,N14288);
and and8606(N14299,N14300,N14301);
and and8613(N14312,N14313,N14314);
and and8620(N14325,N14326,N14327);
and and8627(N14338,N14339,N14340);
and and8634(N14351,N14352,N14353);
and and8641(N14363,N14364,N14365);
and and8648(N14375,N14376,N14377);
and and8655(N14387,N14388,N14389);
and and8662(N14399,N14400,N14401);
and and8669(N14411,N14412,N14413);
and and8676(N14423,N14424,N14425);
and and8683(N14435,N14436,N14437);
and and8690(N14447,N14448,N14449);
and and8697(N14459,N14460,N14461);
and and8704(N14471,N14472,N14473);
and and8711(N14483,N14484,N14485);
and and8718(N14495,N14496,N14497);
and and8725(N14507,N14508,N14509);
and and8732(N14518,N14519,N14520);
and and8739(N14529,N14530,N14531);
and and8746(N14540,N14541,N14542);
and and8753(N14551,N14552,N14553);
and and8760(N14562,N14563,N14564);
and and8767(N14573,N14574,N14575);
and and8774(N14584,N14585,N14586);
and and8781(N14595,N14596,N14597);
and and8788(N14606,N14607,N14608);
and and8795(N14616,N14617,N14618);
and and8802(N14626,N14627,N14628);
and and8809(N14636,N14637,N14638);
and and8816(N14646,N14647,N14648);
and and8823(N14656,N14657,N14658);
and and8830(N14665,N14666,N14667);
and and8837(N14674,N14675,N14676);
and and8844(N14683,N14684,N14685);
and and8851(N14692,N14693,N14694);
and and8858(N14701,N14702,N14703);
and and8865(N14708,N14709,N14710);
and and8871(N14718,N14719,N14720);
and and5055(N8886,N8888,N8889);
and and5056(N8887,N8890,N8891);
and and5064(N8904,N8906,N8907);
and and5065(N8905,N8908,N8909);
and and5073(N8921,N8923,N8924);
and and5074(N8922,N8925,N8926);
and and5082(N8938,N8940,N8941);
and and5083(N8939,N8942,N8943);
and and5091(N8955,N8957,N8958);
and and5092(N8956,N8959,N8960);
and and5100(N8972,N8974,N8975);
and and5101(N8973,N8976,N8977);
and and5109(N8989,N8991,N8992);
and and5110(N8990,N8993,N8994);
and and5118(N9005,N9007,N9008);
and and5119(N9006,N9009,N9010);
and and5127(N9021,N9023,N9024);
and and5128(N9022,N9025,N9026);
and and5136(N9037,N9039,N9040);
and and5137(N9038,N9041,N9042);
and and5145(N9053,N9055,N9056);
and and5146(N9054,N9057,N9058);
and and5154(N9069,N9071,N9072);
and and5155(N9070,N9073,N9074);
and and5163(N9085,N9087,N9088);
and and5164(N9086,N9089,N9090);
and and5172(N9101,N9103,N9104);
and and5173(N9102,N9105,N9106);
and and5181(N9117,N9119,N9120);
and and5182(N9118,N9121,N9122);
and and5190(N9133,N9135,N9136);
and and5191(N9134,N9137,N9138);
and and5199(N9149,N9151,N9152);
and and5200(N9150,N9153,N9154);
and and5208(N9165,N9167,N9168);
and and5209(N9166,N9169,N9170);
and and5217(N9181,N9183,N9184);
and and5218(N9182,N9185,N9186);
and and5226(N9197,N9199,N9200);
and and5227(N9198,N9201,N9202);
and and5235(N9213,N9215,N9216);
and and5236(N9214,N9217,N9218);
and and5244(N9229,N9231,N9232);
and and5245(N9230,N9233,N9234);
and and5253(N9244,N9246,N9247);
and and5254(N9245,N9248,N9249);
and and5262(N9259,N9261,N9262);
and and5263(N9260,N9263,N9264);
and and5271(N9274,N9276,N9277);
and and5272(N9275,N9278,N9279);
and and5280(N9289,N9291,N9292);
and and5281(N9290,N9293,N9294);
and and5289(N9304,N9306,N9307);
and and5290(N9305,N9308,N9309);
and and5298(N9319,N9321,N9322);
and and5299(N9320,N9323,N9324);
and and5307(N9334,N9336,N9337);
and and5308(N9335,N9338,N9339);
and and5316(N9349,N9351,N9352);
and and5317(N9350,N9353,N9354);
and and5325(N9364,N9366,N9367);
and and5326(N9365,N9368,N9369);
and and5334(N9379,N9381,N9382);
and and5335(N9380,N9383,N9384);
and and5343(N9394,N9396,N9397);
and and5344(N9395,N9398,N9399);
and and5352(N9409,N9411,N9412);
and and5353(N9410,N9413,N9414);
and and5361(N9424,N9426,N9427);
and and5362(N9425,N9428,N9429);
and and5370(N9439,N9441,N9442);
and and5371(N9440,N9443,N9444);
and and5379(N9454,N9456,N9457);
and and5380(N9455,N9458,N9459);
and and5388(N9469,N9471,N9472);
and and5389(N9470,N9473,N9474);
and and5397(N9484,N9486,N9487);
and and5398(N9485,N9488,N9489);
and and5406(N9499,N9501,N9502);
and and5407(N9500,N9503,N9504);
and and5415(N9514,N9516,N9517);
and and5416(N9515,N9518,N9519);
and and5424(N9529,N9531,N9532);
and and5425(N9530,N9533,N9534);
and and5433(N9544,N9546,N9547);
and and5434(N9545,N9548,N9549);
and and5442(N9559,N9561,N9562);
and and5443(N9560,N9563,N9564);
and and5451(N9574,N9576,N9577);
and and5452(N9575,N9578,N9579);
and and5460(N9589,N9591,N9592);
and and5461(N9590,N9593,N9594);
and and5469(N9604,N9606,N9607);
and and5470(N9605,N9608,N9609);
and and5478(N9619,N9621,N9622);
and and5479(N9620,N9623,N9624);
and and5487(N9634,N9636,N9637);
and and5488(N9635,N9638,N9639);
and and5496(N9649,N9651,N9652);
and and5497(N9650,N9653,N9654);
and and5505(N9664,N9666,N9667);
and and5506(N9665,N9668,N9669);
and and5514(N9679,N9681,N9682);
and and5515(N9680,N9683,N9684);
and and5523(N9694,N9696,N9697);
and and5524(N9695,N9698,N9699);
and and5532(N9709,N9711,N9712);
and and5533(N9710,N9713,N9714);
and and5541(N9724,N9726,N9727);
and and5542(N9725,N9728,N9729);
and and5550(N9739,N9741,N9742);
and and5551(N9740,N9743,N9744);
and and5559(N9753,N9755,N9756);
and and5560(N9754,N9757,N9758);
and and5568(N9767,N9769,N9770);
and and5569(N9768,N9771,N9772);
and and5577(N9781,N9783,N9784);
and and5578(N9782,N9785,N9786);
and and5586(N9795,N9797,N9798);
and and5587(N9796,N9799,N9800);
and and5595(N9809,N9811,N9812);
and and5596(N9810,N9813,N9814);
and and5604(N9823,N9825,N9826);
and and5605(N9824,N9827,N9828);
and and5613(N9837,N9839,N9840);
and and5614(N9838,N9841,N9842);
and and5622(N9851,N9853,N9854);
and and5623(N9852,N9855,N9856);
and and5631(N9865,N9867,N9868);
and and5632(N9866,N9869,N9870);
and and5640(N9879,N9881,N9882);
and and5641(N9880,N9883,N9884);
and and5649(N9893,N9895,N9896);
and and5650(N9894,N9897,N9898);
and and5658(N9907,N9909,N9910);
and and5659(N9908,N9911,N9912);
and and5667(N9921,N9923,N9924);
and and5668(N9922,N9925,N9926);
and and5676(N9935,N9937,N9938);
and and5677(N9936,N9939,N9940);
and and5685(N9949,N9951,N9952);
and and5686(N9950,N9953,N9954);
and and5694(N9963,N9965,N9966);
and and5695(N9964,N9967,N9968);
and and5703(N9977,N9979,N9980);
and and5704(N9978,N9981,N9982);
and and5712(N9991,N9993,N9994);
and and5713(N9992,N9995,N9996);
and and5721(N10005,N10007,N10008);
and and5722(N10006,N10009,N10010);
and and5730(N10019,N10021,N10022);
and and5731(N10020,N10023,N10024);
and and5739(N10033,N10035,N10036);
and and5740(N10034,N10037,N10038);
and and5748(N10047,N10049,N10050);
and and5749(N10048,N10051,N10052);
and and5757(N10061,N10063,N10064);
and and5758(N10062,N10065,N10066);
and and5766(N10075,N10077,N10078);
and and5767(N10076,N10079,N10080);
and and5775(N10089,N10091,N10092);
and and5776(N10090,N10093,N10094);
and and5784(N10103,N10105,N10106);
and and5785(N10104,N10107,N10108);
and and5793(N10117,N10119,N10120);
and and5794(N10118,N10121,N10122);
and and5802(N10131,N10133,N10134);
and and5803(N10132,N10135,N10136);
and and5811(N10145,N10147,N10148);
and and5812(N10146,N10149,N10150);
and and5820(N10159,N10161,N10162);
and and5821(N10160,N10163,N10164);
and and5829(N10173,N10175,N10176);
and and5830(N10174,N10177,N10178);
and and5838(N10187,N10189,N10190);
and and5839(N10188,N10191,N10192);
and and5847(N10201,N10203,N10204);
and and5848(N10202,N10205,N10206);
and and5856(N10215,N10217,N10218);
and and5857(N10216,N10219,N10220);
and and5865(N10229,N10231,N10232);
and and5866(N10230,N10233,N10234);
and and5874(N10243,N10245,N10246);
and and5875(N10244,N10247,N10248);
and and5883(N10257,N10259,N10260);
and and5884(N10258,N10261,N10262);
and and5892(N10271,N10273,N10274);
and and5893(N10272,N10275,N10276);
and and5901(N10285,N10287,N10288);
and and5902(N10286,N10289,N10290);
and and5910(N10299,N10301,N10302);
and and5911(N10300,N10303,N10304);
and and5919(N10312,N10314,N10315);
and and5920(N10313,N10316,N10317);
and and5928(N10325,N10327,N10328);
and and5929(N10326,N10329,N10330);
and and5937(N10338,N10340,N10341);
and and5938(N10339,N10342,N10343);
and and5946(N10351,N10353,N10354);
and and5947(N10352,N10355,N10356);
and and5955(N10364,N10366,N10367);
and and5956(N10365,N10368,N10369);
and and5964(N10377,N10379,N10380);
and and5965(N10378,N10381,N10382);
and and5973(N10390,N10392,N10393);
and and5974(N10391,N10394,N10395);
and and5982(N10403,N10405,N10406);
and and5983(N10404,N10407,N10408);
and and5991(N10416,N10418,N10419);
and and5992(N10417,N10420,N10421);
and and6000(N10429,N10431,N10432);
and and6001(N10430,N10433,N10434);
and and6009(N10442,N10444,N10445);
and and6010(N10443,N10446,N10447);
and and6018(N10455,N10457,N10458);
and and6019(N10456,N10459,N10460);
and and6027(N10468,N10470,N10471);
and and6028(N10469,N10472,N10473);
and and6036(N10481,N10483,N10484);
and and6037(N10482,N10485,N10486);
and and6045(N10494,N10496,N10497);
and and6046(N10495,N10498,N10499);
and and6054(N10507,N10509,N10510);
and and6055(N10508,N10511,N10512);
and and6063(N10520,N10522,N10523);
and and6064(N10521,N10524,N10525);
and and6072(N10533,N10535,N10536);
and and6073(N10534,N10537,N10538);
and and6081(N10546,N10548,N10549);
and and6082(N10547,N10550,N10551);
and and6090(N10559,N10561,N10562);
and and6091(N10560,N10563,N10564);
and and6099(N10572,N10574,N10575);
and and6100(N10573,N10576,N10577);
and and6108(N10585,N10587,N10588);
and and6109(N10586,N10589,N10590);
and and6117(N10598,N10600,N10601);
and and6118(N10599,N10602,N10603);
and and6126(N10611,N10613,N10614);
and and6127(N10612,N10615,N10616);
and and6135(N10624,N10626,N10627);
and and6136(N10625,N10628,N10629);
and and6144(N10637,N10639,N10640);
and and6145(N10638,N10641,N10642);
and and6153(N10650,N10652,N10653);
and and6154(N10651,N10654,N10655);
and and6162(N10663,N10665,N10666);
and and6163(N10664,N10667,N10668);
and and6171(N10676,N10678,N10679);
and and6172(N10677,N10680,N10681);
and and6180(N10689,N10691,N10692);
and and6181(N10690,N10693,N10694);
and and6189(N10702,N10704,N10705);
and and6190(N10703,N10706,N10707);
and and6198(N10715,N10717,N10718);
and and6199(N10716,N10719,N10720);
and and6207(N10728,N10730,N10731);
and and6208(N10729,N10732,N10733);
and and6216(N10741,N10743,N10744);
and and6217(N10742,N10745,N10746);
and and6225(N10754,N10756,N10757);
and and6226(N10755,N10758,N10759);
and and6234(N10767,N10769,N10770);
and and6235(N10768,N10771,N10772);
and and6243(N10780,N10782,N10783);
and and6244(N10781,N10784,N10785);
and and6252(N10793,N10795,N10796);
and and6253(N10794,N10797,N10798);
and and6261(N10806,N10808,N10809);
and and6262(N10807,N10810,N10811);
and and6270(N10819,N10821,N10822);
and and6271(N10820,N10823,N10824);
and and6279(N10831,N10833,N10834);
and and6280(N10832,N10835,N10836);
and and6288(N10843,N10845,N10846);
and and6289(N10844,N10847,N10848);
and and6297(N10855,N10857,N10858);
and and6298(N10856,N10859,N10860);
and and6306(N10867,N10869,N10870);
and and6307(N10868,N10871,N10872);
and and6315(N10879,N10881,N10882);
and and6316(N10880,N10883,N10884);
and and6324(N10891,N10893,N10894);
and and6325(N10892,N10895,N10896);
and and6333(N10903,N10905,N10906);
and and6334(N10904,N10907,N10908);
and and6342(N10915,N10917,N10918);
and and6343(N10916,N10919,N10920);
and and6351(N10927,N10929,N10930);
and and6352(N10928,N10931,N10932);
and and6360(N10939,N10941,N10942);
and and6361(N10940,N10943,N10944);
and and6369(N10951,N10953,N10954);
and and6370(N10952,N10955,N10956);
and and6378(N10963,N10965,N10966);
and and6379(N10964,N10967,N10968);
and and6387(N10975,N10977,N10978);
and and6388(N10976,N10979,N10980);
and and6396(N10987,N10989,N10990);
and and6397(N10988,N10991,N10992);
and and6405(N10999,N11001,N11002);
and and6406(N11000,N11003,N11004);
and and6414(N11011,N11013,N11014);
and and6415(N11012,N11015,N11016);
and and6423(N11023,N11025,N11026);
and and6424(N11024,N11027,N11028);
and and6432(N11035,N11037,N11038);
and and6433(N11036,N11039,N11040);
and and6441(N11047,N11049,N11050);
and and6442(N11048,N11051,N11052);
and and6450(N11059,N11061,N11062);
and and6451(N11060,N11063,N11064);
and and6459(N11071,N11073,N11074);
and and6460(N11072,N11075,N11076);
and and6468(N11083,N11085,N11086);
and and6469(N11084,N11087,N11088);
and and6477(N11095,N11097,N11098);
and and6478(N11096,N11099,N11100);
and and6486(N11107,N11109,N11110);
and and6487(N11108,N11111,N11112);
and and6495(N11119,N11121,N11122);
and and6496(N11120,N11123,N11124);
and and6504(N11131,N11133,N11134);
and and6505(N11132,N11135,N11136);
and and6513(N11143,N11145,N11146);
and and6514(N11144,N11147,N11148);
and and6522(N11154,N11156,N11157);
and and6523(N11155,N11158,N11159);
and and6531(N11165,N11167,N11168);
and and6532(N11166,N11169,N11170);
and and6540(N11176,N11178,N11179);
and and6541(N11177,N11180,N11181);
and and6549(N11187,N11189,N11190);
and and6550(N11188,N11191,N11192);
and and6558(N11198,N11200,N11201);
and and6559(N11199,N11202,N11203);
and and6567(N11209,N11211,N11212);
and and6568(N11210,N11213,N11214);
and and6576(N11220,N11222,N11223);
and and6577(N11221,N11224,N11225);
and and6585(N11231,N11233,N11234);
and and6586(N11232,N11235,N11236);
and and6594(N11242,N11244,N11245);
and and6595(N11243,N11246,N11247);
and and6603(N11253,N11255,N11256);
and and6604(N11254,N11257,N11258);
and and6612(N11264,N11266,N11267);
and and6613(N11265,N11268,N11269);
and and6621(N11275,N11277,N11278);
and and6622(N11276,N11279,N11280);
and and6630(N11286,N11288,N11289);
and and6631(N11287,N11290,N11291);
and and6639(N11297,N11299,N11300);
and and6640(N11298,N11301,N11302);
and and6648(N11308,N11310,N11311);
and and6649(N11309,N11312,N11313);
and and6657(N11319,N11321,N11322);
and and6658(N11320,N11323,N11324);
and and6666(N11329,N11331,N11332);
and and6667(N11330,N11333,N11334);
and and6675(N11339,N11341,N11342);
and and6676(N11340,N11343,N11344);
and and6684(N11349,N11351,N11352);
and and6685(N11350,N11353,N11354);
and and6693(N11359,N11361,N11362);
and and6694(N11360,N11363,N11364);
and and6702(N11369,N11371,N11372);
and and6703(N11370,N11373,N11374);
and and6710(N11385,N11387,N11388);
and and6711(N11386,N11389,N11390);
and and6718(N11401,N11403,N11404);
and and6719(N11402,N11405,N11406);
and and6726(N11417,N11419,N11420);
and and6727(N11418,N11421,N11422);
and and6734(N11433,N11435,N11436);
and and6735(N11434,N11437,N11438);
and and6742(N11449,N11451,N11452);
and and6743(N11450,N11453,N11454);
and and6750(N11465,N11467,N11468);
and and6751(N11466,N11469,N11470);
and and6758(N11481,N11483,N11484);
and and6759(N11482,N11485,N11486);
and and6766(N11496,N11498,N11499);
and and6767(N11497,N11500,N11501);
and and6774(N11511,N11513,N11514);
and and6775(N11512,N11515,N11516);
and and6782(N11526,N11528,N11529);
and and6783(N11527,N11530,N11531);
and and6790(N11541,N11543,N11544);
and and6791(N11542,N11545,N11546);
and and6798(N11556,N11558,N11559);
and and6799(N11557,N11560,N11561);
and and6806(N11571,N11573,N11574);
and and6807(N11572,N11575,N11576);
and and6814(N11586,N11588,N11589);
and and6815(N11587,N11590,N11591);
and and6822(N11600,N11602,N11603);
and and6823(N11601,N11604,N11605);
and and6830(N11614,N11616,N11617);
and and6831(N11615,N11618,N11619);
and and6838(N11628,N11630,N11631);
and and6839(N11629,N11632,N11633);
and and6846(N11642,N11644,N11645);
and and6847(N11643,N11646,N11647);
and and6854(N11656,N11658,N11659);
and and6855(N11657,N11660,N11661);
and and6862(N11670,N11672,N11673);
and and6863(N11671,N11674,N11675);
and and6870(N11684,N11686,N11687);
and and6871(N11685,N11688,N11689);
and and6878(N11698,N11700,N11701);
and and6879(N11699,N11702,N11703);
and and6886(N11712,N11714,N11715);
and and6887(N11713,N11716,N11717);
and and6894(N11726,N11728,N11729);
and and6895(N11727,N11730,N11731);
and and6902(N11740,N11742,N11743);
and and6903(N11741,N11744,N11745);
and and6910(N11754,N11756,N11757);
and and6911(N11755,N11758,N11759);
and and6918(N11768,N11770,N11771);
and and6919(N11769,N11772,N11773);
and and6926(N11782,N11784,N11785);
and and6927(N11783,N11786,N11787);
and and6934(N11796,N11798,N11799);
and and6935(N11797,N11800,N11801);
and and6942(N11810,N11812,N11813);
and and6943(N11811,N11814,N11815);
and and6950(N11824,N11826,N11827);
and and6951(N11825,N11828,N11829);
and and6958(N11838,N11840,N11841);
and and6959(N11839,N11842,N11843);
and and6966(N11852,N11854,N11855);
and and6967(N11853,N11856,N11857);
and and6974(N11866,N11868,N11869);
and and6975(N11867,N11870,N11871);
and and6982(N11880,N11882,N11883);
and and6983(N11881,N11884,N11885);
and and6990(N11894,N11896,N11897);
and and6991(N11895,N11898,N11899);
and and6998(N11908,N11910,N11911);
and and6999(N11909,N11912,N11913);
and and7006(N11922,N11924,N11925);
and and7007(N11923,N11926,N11927);
and and7014(N11936,N11938,N11939);
and and7015(N11937,N11940,N11941);
and and7022(N11950,N11952,N11953);
and and7023(N11951,N11954,N11955);
and and7030(N11964,N11966,N11967);
and and7031(N11965,N11968,N11969);
and and7038(N11978,N11980,N11981);
and and7039(N11979,N11982,N11983);
and and7046(N11992,N11994,N11995);
and and7047(N11993,N11996,N11997);
and and7054(N12006,N12008,N12009);
and and7055(N12007,N12010,N12011);
and and7062(N12020,N12022,N12023);
and and7063(N12021,N12024,N12025);
and and7070(N12034,N12036,N12037);
and and7071(N12035,N12038,N12039);
and and7078(N12048,N12050,N12051);
and and7079(N12049,N12052,N12053);
and and7086(N12062,N12064,N12065);
and and7087(N12063,N12066,N12067);
and and7094(N12076,N12078,N12079);
and and7095(N12077,N12080,N12081);
and and7102(N12089,N12091,N12092);
and and7103(N12090,N12093,N12094);
and and7110(N12102,N12104,N12105);
and and7111(N12103,N12106,N12107);
and and7118(N12115,N12117,N12118);
and and7119(N12116,N12119,N12120);
and and7126(N12128,N12130,N12131);
and and7127(N12129,N12132,N12133);
and and7134(N12141,N12143,N12144);
and and7135(N12142,N12145,N12146);
and and7142(N12154,N12156,N12157);
and and7143(N12155,N12158,N12159);
and and7150(N12167,N12169,N12170);
and and7151(N12168,N12171,N12172);
and and7158(N12180,N12182,N12183);
and and7159(N12181,N12184,N12185);
and and7166(N12193,N12195,N12196);
and and7167(N12194,N12197,N12198);
and and7174(N12206,N12208,N12209);
and and7175(N12207,N12210,N12211);
and and7182(N12219,N12221,N12222);
and and7183(N12220,N12223,N12224);
and and7190(N12232,N12234,N12235);
and and7191(N12233,N12236,N12237);
and and7198(N12245,N12247,N12248);
and and7199(N12246,N12249,N12250);
and and7206(N12258,N12260,N12261);
and and7207(N12259,N12262,N12263);
and and7214(N12271,N12273,N12274);
and and7215(N12272,N12275,N12276);
and and7222(N12284,N12286,N12287);
and and7223(N12285,N12288,N12289);
and and7230(N12297,N12299,N12300);
and and7231(N12298,N12301,N12302);
and and7238(N12310,N12312,N12313);
and and7239(N12311,N12314,N12315);
and and7246(N12323,N12325,N12326);
and and7247(N12324,N12327,N12328);
and and7254(N12336,N12338,N12339);
and and7255(N12337,N12340,N12341);
and and7262(N12349,N12351,N12352);
and and7263(N12350,N12353,N12354);
and and7270(N12362,N12364,N12365);
and and7271(N12363,N12366,N12367);
and and7278(N12375,N12377,N12378);
and and7279(N12376,N12379,N12380);
and and7286(N12388,N12390,N12391);
and and7287(N12389,N12392,N12393);
and and7294(N12401,N12403,N12404);
and and7295(N12402,N12405,N12406);
and and7302(N12414,N12416,N12417);
and and7303(N12415,N12418,N12419);
and and7310(N12427,N12429,N12430);
and and7311(N12428,N12431,N12432);
and and7318(N12440,N12442,N12443);
and and7319(N12441,N12444,N12445);
and and7326(N12453,N12455,N12456);
and and7327(N12454,N12457,N12458);
and and7334(N12466,N12468,N12469);
and and7335(N12467,N12470,N12471);
and and7342(N12479,N12481,N12482);
and and7343(N12480,N12483,N12484);
and and7350(N12492,N12494,N12495);
and and7351(N12493,N12496,N12497);
and and7358(N12505,N12507,N12508);
and and7359(N12506,N12509,N12510);
and and7366(N12518,N12520,N12521);
and and7367(N12519,N12522,N12523);
and and7374(N12531,N12533,N12534);
and and7375(N12532,N12535,N12536);
and and7382(N12544,N12546,N12547);
and and7383(N12545,N12548,N12549);
and and7390(N12557,N12559,N12560);
and and7391(N12558,N12561,N12562);
and and7398(N12570,N12572,N12573);
and and7399(N12571,N12574,N12575);
and and7406(N12583,N12585,N12586);
and and7407(N12584,N12587,N12588);
and and7414(N12596,N12598,N12599);
and and7415(N12597,N12600,N12601);
and and7422(N12609,N12611,N12612);
and and7423(N12610,N12613,N12614);
and and7430(N12622,N12624,N12625);
and and7431(N12623,N12626,N12627);
and and7438(N12635,N12637,N12638);
and and7439(N12636,N12639,N12640);
and and7446(N12648,N12650,N12651);
and and7447(N12649,N12652,N12653);
and and7454(N12661,N12663,N12664);
and and7455(N12662,N12665,N12666);
and and7462(N12674,N12676,N12677);
and and7463(N12675,N12678,N12679);
and and7470(N12686,N12688,N12689);
and and7471(N12687,N12690,N12691);
and and7478(N12698,N12700,N12701);
and and7479(N12699,N12702,N12703);
and and7486(N12710,N12712,N12713);
and and7487(N12711,N12714,N12715);
and and7494(N12722,N12724,N12725);
and and7495(N12723,N12726,N12727);
and and7502(N12734,N12736,N12737);
and and7503(N12735,N12738,N12739);
and and7510(N12746,N12748,N12749);
and and7511(N12747,N12750,N12751);
and and7518(N12758,N12760,N12761);
and and7519(N12759,N12762,N12763);
and and7526(N12770,N12772,N12773);
and and7527(N12771,N12774,N12775);
and and7534(N12782,N12784,N12785);
and and7535(N12783,N12786,N12787);
and and7542(N12794,N12796,N12797);
and and7543(N12795,N12798,N12799);
and and7550(N12806,N12808,N12809);
and and7551(N12807,N12810,N12811);
and and7558(N12818,N12820,N12821);
and and7559(N12819,N12822,N12823);
and and7566(N12830,N12832,N12833);
and and7567(N12831,N12834,N12835);
and and7574(N12842,N12844,N12845);
and and7575(N12843,N12846,N12847);
and and7582(N12854,N12856,N12857);
and and7583(N12855,N12858,N12859);
and and7590(N12866,N12868,N12869);
and and7591(N12867,N12870,N12871);
and and7598(N12878,N12880,N12881);
and and7599(N12879,N12882,N12883);
and and7606(N12890,N12892,N12893);
and and7607(N12891,N12894,N12895);
and and7614(N12902,N12904,N12905);
and and7615(N12903,N12906,N12907);
and and7622(N12914,N12916,N12917);
and and7623(N12915,N12918,N12919);
and and7630(N12926,N12928,N12929);
and and7631(N12927,N12930,N12931);
and and7638(N12938,N12940,N12941);
and and7639(N12939,N12942,N12943);
and and7646(N12950,N12952,N12953);
and and7647(N12951,N12954,N12955);
and and7654(N12962,N12964,N12965);
and and7655(N12963,N12966,N12967);
and and7662(N12974,N12976,N12977);
and and7663(N12975,N12978,N12979);
and and7670(N12986,N12988,N12989);
and and7671(N12987,N12990,N12991);
and and7678(N12998,N13000,N13001);
and and7679(N12999,N13002,N13003);
and and7686(N13010,N13012,N13013);
and and7687(N13011,N13014,N13015);
and and7694(N13022,N13024,N13025);
and and7695(N13023,N13026,N13027);
and and7702(N13034,N13036,N13037);
and and7703(N13035,N13038,N13039);
and and7710(N13046,N13048,N13049);
and and7711(N13047,N13050,N13051);
and and7718(N13058,N13060,N13061);
and and7719(N13059,N13062,N13063);
and and7726(N13070,N13072,N13073);
and and7727(N13071,N13074,N13075);
and and7734(N13082,N13084,N13085);
and and7735(N13083,N13086,N13087);
and and7742(N13094,N13096,N13097);
and and7743(N13095,N13098,N13099);
and and7750(N13106,N13108,N13109);
and and7751(N13107,N13110,N13111);
and and7758(N13118,N13120,N13121);
and and7759(N13119,N13122,N13123);
and and7766(N13130,N13132,N13133);
and and7767(N13131,N13134,N13135);
and and7774(N13142,N13144,N13145);
and and7775(N13143,N13146,N13147);
and and7782(N13154,N13156,N13157);
and and7783(N13155,N13158,N13159);
and and7790(N13166,N13168,N13169);
and and7791(N13167,N13170,N13171);
and and7798(N13178,N13180,N13181);
and and7799(N13179,N13182,N13183);
and and7806(N13190,N13192,N13193);
and and7807(N13191,N13194,N13195);
and and7814(N13202,N13204,N13205);
and and7815(N13203,N13206,N13207);
and and7822(N13214,N13216,N13217);
and and7823(N13215,N13218,N13219);
and and7830(N13226,N13228,N13229);
and and7831(N13227,N13230,N13231);
and and7838(N13238,N13240,N13241);
and and7839(N13239,N13242,N13243);
and and7846(N13250,N13252,N13253);
and and7847(N13251,N13254,N13255);
and and7854(N13262,N13264,N13265);
and and7855(N13263,N13266,N13267);
and and7862(N13274,N13276,N13277);
and and7863(N13275,N13278,N13279);
and and7870(N13286,N13288,N13289);
and and7871(N13287,N13290,N13291);
and and7878(N13298,N13300,N13301);
and and7879(N13299,N13302,N13303);
and and7886(N13310,N13312,N13313);
and and7887(N13311,N13314,N13315);
and and7894(N13322,N13324,N13325);
and and7895(N13323,N13326,N13327);
and and7902(N13334,N13336,N13337);
and and7903(N13335,N13338,N13339);
and and7910(N13346,N13348,N13349);
and and7911(N13347,N13350,N13351);
and and7918(N13358,N13360,N13361);
and and7919(N13359,N13362,N13363);
and and7926(N13370,N13372,N13373);
and and7927(N13371,N13374,N13375);
and and7934(N13382,N13384,N13385);
and and7935(N13383,N13386,N13387);
and and7942(N13394,N13396,N13397);
and and7943(N13395,N13398,N13399);
and and7950(N13405,N13407,N13408);
and and7951(N13406,N13409,N13410);
and and7958(N13416,N13418,N13419);
and and7959(N13417,N13420,N13421);
and and7966(N13427,N13429,N13430);
and and7967(N13428,N13431,N13432);
and and7974(N13438,N13440,N13441);
and and7975(N13439,N13442,N13443);
and and7982(N13449,N13451,N13452);
and and7983(N13450,N13453,N13454);
and and7990(N13460,N13462,N13463);
and and7991(N13461,N13464,N13465);
and and7998(N13471,N13473,N13474);
and and7999(N13472,N13475,N13476);
and and8006(N13482,N13484,N13485);
and and8007(N13483,N13486,N13487);
and and8014(N13493,N13495,N13496);
and and8015(N13494,N13497,N13498);
and and8022(N13504,N13506,N13507);
and and8023(N13505,N13508,N13509);
and and8030(N13515,N13517,N13518);
and and8031(N13516,N13519,N13520);
and and8038(N13526,N13528,N13529);
and and8039(N13527,N13530,N13531);
and and8046(N13537,N13539,N13540);
and and8047(N13538,N13541,N13542);
and and8054(N13548,N13550,N13551);
and and8055(N13549,N13552,N13553);
and and8062(N13559,N13561,N13562);
and and8063(N13560,N13563,N13564);
and and8070(N13570,N13572,N13573);
and and8071(N13571,N13574,N13575);
and and8078(N13581,N13583,N13584);
and and8079(N13582,N13585,N13586);
and and8086(N13592,N13594,N13595);
and and8087(N13593,N13596,N13597);
and and8094(N13603,N13605,N13606);
and and8095(N13604,N13607,N13608);
and and8102(N13614,N13616,N13617);
and and8103(N13615,N13618,N13619);
and and8110(N13625,N13627,N13628);
and and8111(N13626,N13629,N13630);
and and8118(N13636,N13638,N13639);
and and8119(N13637,N13640,N13641);
and and8126(N13647,N13649,N13650);
and and8127(N13648,N13651,N13652);
and and8134(N13658,N13660,N13661);
and and8135(N13659,N13662,N13663);
and and8142(N13669,N13671,N13672);
and and8143(N13670,N13673,N13674);
and and8150(N13680,N13682,N13683);
and and8151(N13681,N13684,N13685);
and and8158(N13691,N13693,N13694);
and and8159(N13692,N13695,N13696);
and and8166(N13702,N13704,N13705);
and and8167(N13703,N13706,N13707);
and and8174(N13713,N13715,N13716);
and and8175(N13714,N13717,N13718);
and and8182(N13724,N13726,N13727);
and and8183(N13725,N13728,N13729);
and and8190(N13735,N13737,N13738);
and and8191(N13736,N13739,N13740);
and and8198(N13746,N13748,N13749);
and and8199(N13747,N13750,N13751);
and and8206(N13757,N13759,N13760);
and and8207(N13758,N13761,N13762);
and and8214(N13768,N13770,N13771);
and and8215(N13769,N13772,N13773);
and and8222(N13779,N13781,N13782);
and and8223(N13780,N13783,N13784);
and and8230(N13790,N13792,N13793);
and and8231(N13791,N13794,N13795);
and and8238(N13801,N13803,N13804);
and and8239(N13802,N13805,N13806);
and and8246(N13812,N13814,N13815);
and and8247(N13813,N13816,N13817);
and and8254(N13823,N13825,N13826);
and and8255(N13824,N13827,N13828);
and and8262(N13834,N13836,N13837);
and and8263(N13835,N13838,N13839);
and and8270(N13845,N13847,N13848);
and and8271(N13846,N13849,N13850);
and and8278(N13856,N13858,N13859);
and and8279(N13857,N13860,N13861);
and and8286(N13867,N13869,N13870);
and and8287(N13868,N13871,N13872);
and and8294(N13878,N13880,N13881);
and and8295(N13879,N13882,N13883);
and and8302(N13889,N13891,N13892);
and and8303(N13890,N13893,N13894);
and and8310(N13900,N13902,N13903);
and and8311(N13901,N13904,N13905);
and and8318(N13911,N13913,N13914);
and and8319(N13912,N13915,N13916);
and and8326(N13922,N13924,N13925);
and and8327(N13923,N13926,N13927);
and and8334(N13933,N13935,N13936);
and and8335(N13934,N13937,N13938);
and and8342(N13944,N13946,N13947);
and and8343(N13945,N13948,N13949);
and and8350(N13955,N13957,N13958);
and and8351(N13956,N13959,N13960);
and and8358(N13965,N13967,N13968);
and and8359(N13966,N13969,N13970);
and and8366(N13975,N13977,N13978);
and and8367(N13976,N13979,N13980);
and and8374(N13985,N13987,N13988);
and and8375(N13986,N13989,N13990);
and and8382(N13995,N13997,N13998);
and and8383(N13996,N13999,N14000);
and and8390(N14005,N14007,N14008);
and and8391(N14006,N14009,N14010);
and and8398(N14015,N14017,N14018);
and and8399(N14016,N14019,N14020);
and and8406(N14025,N14027,N14028);
and and8407(N14026,N14029,N14030);
and and8414(N14035,N14037,N14038);
and and8415(N14036,N14039,N14040);
and and8422(N14045,N14047,N14048);
and and8423(N14046,N14049,N14050);
and and8430(N14055,N14057,N14058);
and and8431(N14056,N14059,N14060);
and and8438(N14065,N14067,N14068);
and and8439(N14066,N14069,N14070);
and and8446(N14075,N14077,N14078);
and and8447(N14076,N14079,N14080);
and and8454(N14085,N14087,N14088);
and and8455(N14086,N14089,N14090);
and and8462(N14095,N14097,N14098);
and and8463(N14096,N14099,N14100);
and and8470(N14105,N14107,N14108);
and and8471(N14106,N14109,N14110);
and and8478(N14115,N14117,N14118);
and and8479(N14116,N14119,N14120);
and and8486(N14124,N14126,N14127);
and and8487(N14125,N14128,N14129);
and and8494(N14133,N14135,N14136);
and and8495(N14134,N14137,N14138);
and and8502(N14142,N14144,N14145);
and and8503(N14143,N14146,N14147);
and and8510(N14151,N14153,N14154);
and and8511(N14152,N14155,N14156);
and and8518(N14160,N14162,N14163);
and and8519(N14161,N14164,N14165);
and and8526(N14169,N14171,N14172);
and and8527(N14170,N14173,N14174);
and and8534(N14178,N14180,N14181);
and and8535(N14179,N14182,N14183);
and and8542(N14187,N14189,N14190);
and and8543(N14188,N14191,N14192);
and and8550(N14196,N14198,N14199);
and and8551(N14197,N14200,N14201);
and and8558(N14205,N14207,N14208);
and and8559(N14206,N14209,N14210);
and and8565(N14219,N14221,N14222);
and and8566(N14220,N14223,N14224);
and and8572(N14233,N14235,N14236);
and and8573(N14234,N14237,N14238);
and and8579(N14247,N14249,N14250);
and and8580(N14248,N14251,N14252);
and and8586(N14261,N14263,N14264);
and and8587(N14262,N14265,N14266);
and and8593(N14274,N14276,N14277);
and and8594(N14275,N14278,N14279);
and and8600(N14287,N14289,N14290);
and and8601(N14288,N14291,N14292);
and and8607(N14300,N14302,N14303);
and and8608(N14301,N14304,N14305);
and and8614(N14313,N14315,N14316);
and and8615(N14314,N14317,N14318);
and and8621(N14326,N14328,N14329);
and and8622(N14327,N14330,N14331);
and and8628(N14339,N14341,N14342);
and and8629(N14340,N14343,N14344);
and and8635(N14352,N14354,N14355);
and and8636(N14353,N14356,N14357);
and and8642(N14364,N14366,N14367);
and and8643(N14365,N14368,N14369);
and and8649(N14376,N14378,N14379);
and and8650(N14377,N14380,N14381);
and and8656(N14388,N14390,N14391);
and and8657(N14389,N14392,N14393);
and and8663(N14400,N14402,N14403);
and and8664(N14401,N14404,N14405);
and and8670(N14412,N14414,N14415);
and and8671(N14413,N14416,N14417);
and and8677(N14424,N14426,N14427);
and and8678(N14425,N14428,N14429);
and and8684(N14436,N14438,N14439);
and and8685(N14437,N14440,N14441);
and and8691(N14448,N14450,N14451);
and and8692(N14449,N14452,N14453);
and and8698(N14460,N14462,N14463);
and and8699(N14461,N14464,N14465);
and and8705(N14472,N14474,N14475);
and and8706(N14473,N14476,N14477);
and and8712(N14484,N14486,N14487);
and and8713(N14485,N14488,N14489);
and and8719(N14496,N14498,N14499);
and and8720(N14497,N14500,N14501);
and and8726(N14508,N14510,N14511);
and and8727(N14509,N14512,N14513);
and and8733(N14519,N14521,N14522);
and and8734(N14520,N14523,N14524);
and and8740(N14530,N14532,N14533);
and and8741(N14531,N14534,N14535);
and and8747(N14541,N14543,N14544);
and and8748(N14542,N14545,N14546);
and and8754(N14552,N14554,N14555);
and and8755(N14553,N14556,N14557);
and and8761(N14563,N14565,N14566);
and and8762(N14564,N14567,N14568);
and and8768(N14574,N14576,N14577);
and and8769(N14575,N14578,N14579);
and and8775(N14585,N14587,N14588);
and and8776(N14586,N14589,N14590);
and and8782(N14596,N14598,N14599);
and and8783(N14597,N14600,N14601);
and and8789(N14607,N14609,N14610);
and and8790(N14608,N14611,N14612);
and and8796(N14617,N14619,N14620);
and and8797(N14618,N14621,N14622);
and and8803(N14627,N14629,N14630);
and and8804(N14628,N14631,N14632);
and and8810(N14637,N14639,N14640);
and and8811(N14638,N14641,N14642);
and and8817(N14647,N14649,N14650);
and and8818(N14648,N14651,N14652);
and and8824(N14657,N14659,N14660);
and and8825(N14658,N14661,N14662);
and and8831(N14666,N14668,N14669);
and and8832(N14667,N14670,N14671);
and and8838(N14675,N14677,N14678);
and and8839(N14676,N14679,N14680);
and and8845(N14684,N14686,N14687);
and and8846(N14685,N14688,N14689);
and and8852(N14693,N14695,N14696);
and and8853(N14694,N14697,N14698);
and and8859(N14702,N14704,N14705);
and and8860(N14703,N14706,N14707);
and and8866(N14709,N14711,N14712);
and and8867(N14710,N14713,R0);
and and8872(N14719,N14721,N14722);
and and8873(N14720,N14723,in0);
and and5057(N8888,N8892,N8893);
and and5058(N8889,N8894,N8895);
and and5059(N8890,N8896,N8897);
and and5060(N8891,N8898,N8899);
and and5066(N8906,N8910,N8911);
and and5067(N8907,N8912,N8913);
and and5068(N8908,R0,N8914);
and and5069(N8909,N8915,R3);
and and5075(N8923,N8927,N8928);
and and5076(N8924,N8929,N8930);
and and5077(N8925,N8931,N8932);
and and5078(N8926,N8933,R2);
and and5084(N8940,N8944,N8945);
and and5085(N8941,N8946,N8947);
and and5086(N8942,in2,N8948);
and and5087(N8943,N8949,N8950);
and and5093(N8957,N8961,N8962);
and and5094(N8958,N8963,N8964);
and and5095(N8959,N8965,N8966);
and and5096(N8960,N8967,N8968);
and and5102(N8974,N8978,N8979);
and and5103(N8975,N8980,N8981);
and and5104(N8976,N8982,N8983);
and and5105(N8977,R2,N8984);
and and5111(N8991,N8995,N8996);
and and5112(N8992,in0,N8997);
and and5113(N8993,N8998,R1);
and and5114(N8994,N8999,R3);
and and5120(N9007,N9011,N9012);
and and5121(N9008,in1,in2);
and and5122(N9009,N9013,R1);
and and5123(N9010,N9014,N9015);
and and5129(N9023,N9027,N9028);
and and5130(N9024,N9029,N9030);
and and5131(N9025,N9031,N9032);
and and5132(N9026,R2,N9033);
and and5138(N9039,N9043,N9044);
and and5139(N9040,in0,in1);
and and5140(N9041,N9045,N9046);
and and5141(N9042,N9047,N9048);
and and5147(N9055,N9059,N9060);
and and5148(N9056,in0,N9061);
and and5149(N9057,R0,N9062);
and and5150(N9058,N9063,N9064);
and and5156(N9071,N9075,N9076);
and and5157(N9072,in0,in1);
and and5158(N9073,in2,N9077);
and and5159(N9074,N9078,N9079);
and and5165(N9087,N9091,N9092);
and and5166(N9088,in1,in2);
and and5167(N9089,N9093,N9094);
and and5168(N9090,N9095,N9096);
and and5174(N9103,N9107,N9108);
and and5175(N9104,in0,N9109);
and and5176(N9105,R0,R1);
and and5177(N9106,N9110,N9111);
and and5183(N9119,N9123,N9124);
and and5184(N9120,N9125,in2);
and and5185(N9121,R0,R1);
and and5186(N9122,N9126,N9127);
and and5192(N9135,N9139,N9140);
and and5193(N9136,N9141,N9142);
and and5194(N9137,in2,N9143);
and and5195(N9138,N9144,R2);
and and5201(N9151,N9155,N9156);
and and5202(N9152,N9157,in2);
and and5203(N9153,R0,N9158);
and and5204(N9154,N9159,N9160);
and and5210(N9167,N9171,N9172);
and and5211(N9168,N9173,N9174);
and and5212(N9169,N9175,R0);
and and5213(N9170,N9176,N9177);
and and5219(N9183,N9187,N9188);
and and5220(N9184,N9189,N9190);
and and5221(N9185,in2,N9191);
and and5222(N9186,N9192,N9193);
and and5228(N9199,N9203,N9204);
and and5229(N9200,N9205,N9206);
and and5230(N9201,R0,R1);
and and5231(N9202,N9207,N9208);
and and5237(N9215,N9219,N9220);
and and5238(N9216,N9221,N9222);
and and5239(N9217,N9223,N9224);
and and5240(N9218,N9225,R2);
and and5246(N9231,N9235,N9236);
and and5247(N9232,N9237,N9238);
and and5248(N9233,N9239,R0);
and and5249(N9234,N9240,R2);
and and5255(N9246,N9250,N9251);
and and5256(N9247,N9252,N9253);
and and5257(N9248,N9254,R0);
and and5258(N9249,N9255,R2);
and and5264(N9261,N9265,N9266);
and and5265(N9262,in1,N9267);
and and5266(N9263,N9268,R1);
and and5267(N9264,N9269,R3);
and and5273(N9276,N9280,N9281);
and and5274(N9277,N9282,N9283);
and and5275(N9278,N9284,N9285);
and and5276(N9279,N9286,R3);
and and5282(N9291,N9295,N9296);
and and5283(N9292,in0,N9297);
and and5284(N9293,N9298,N9299);
and and5285(N9294,R2,N9300);
and and5291(N9306,N9310,N9311);
and and5292(N9307,N9312,N9313);
and and5293(N9308,N9314,N9315);
and and5294(N9309,R1,R2);
and and5300(N9321,N9325,N9326);
and and5301(N9322,N9327,in2);
and and5302(N9323,R0,R1);
and and5303(N9324,N9328,N9329);
and and5309(N9336,N9340,N9341);
and and5310(N9337,N9342,in2);
and and5311(N9338,N9343,N9344);
and and5312(N9339,R2,R3);
and and5318(N9351,N9355,N9356);
and and5319(N9352,N9357,in1);
and and5320(N9353,N9358,N9359);
and and5321(N9354,R2,R3);
and and5327(N9366,N9370,N9371);
and and5328(N9367,N9372,in1);
and and5329(N9368,in2,N9373);
and and5330(N9369,R2,R3);
and and5336(N9381,N9385,N9386);
and and5337(N9382,in1,N9387);
and and5338(N9383,N9388,R1);
and and5339(N9384,N9389,N9390);
and and5345(N9396,N9400,N9401);
and and5346(N9397,N9402,N9403);
and and5347(N9398,N9404,R0);
and and5348(N9399,R2,N9405);
and and5354(N9411,N9415,N9416);
and and5355(N9412,N9417,N9418);
and and5356(N9413,N9419,R0);
and and5357(N9414,N9420,N9421);
and and5363(N9426,N9430,N9431);
and and5364(N9427,N9432,N9433);
and and5365(N9428,N9434,R0);
and and5366(N9429,R2,N9435);
and and5372(N9441,N9445,N9446);
and and5373(N9442,N9447,in2);
and and5374(N9443,N9448,N9449);
and and5375(N9444,N9450,R3);
and and5381(N9456,N9460,N9461);
and and5382(N9457,in1,N9462);
and and5383(N9458,N9463,N9464);
and and5384(N9459,N9465,R3);
and and5390(N9471,N9475,N9476);
and and5391(N9472,in1,N9477);
and and5392(N9473,R0,N9478);
and and5393(N9474,R2,N9479);
and and5399(N9486,N9490,N9491);
and and5400(N9487,N9492,N9493);
and and5401(N9488,R0,R1);
and and5402(N9489,N9494,N9495);
and and5408(N9501,N9505,N9506);
and and5409(N9502,N9507,N9508);
and and5410(N9503,N9509,R0);
and and5411(N9504,N9510,R2);
and and5417(N9516,N9520,N9521);
and and5418(N9517,N9522,N9523);
and and5419(N9518,N9524,R0);
and and5420(N9519,R1,R2);
and and5426(N9531,N9535,N9536);
and and5427(N9532,N9537,in2);
and and5428(N9533,N9538,N9539);
and and5429(N9534,R2,R3);
and and5435(N9546,N9550,N9551);
and and5436(N9547,N9552,N9553);
and and5437(N9548,in2,R0);
and and5438(N9549,N9554,N9555);
and and5444(N9561,N9565,N9566);
and and5445(N9562,N9567,in1);
and and5446(N9563,N9568,R0);
and and5447(N9564,N9569,R3);
and and5453(N9576,N9580,N9581);
and and5454(N9577,N9582,N9583);
and and5455(N9578,in2,R0);
and and5456(N9579,N9584,N9585);
and and5462(N9591,N9595,N9596);
and and5463(N9592,N9597,N9598);
and and5464(N9593,N9599,R0);
and and5465(N9594,N9600,N9601);
and and5471(N9606,N9610,N9611);
and and5472(N9607,N9612,in1);
and and5473(N9608,N9613,N9614);
and and5474(N9609,N9615,R3);
and and5480(N9621,N9625,N9626);
and and5481(N9622,N9627,N9628);
and and5482(N9623,in2,R0);
and and5483(N9624,N9629,N9630);
and and5489(N9636,N9640,N9641);
and and5490(N9637,N9642,N9643);
and and5491(N9638,N9644,N9645);
and and5492(N9639,R1,R2);
and and5498(N9651,N9655,N9656);
and and5499(N9652,N9657,N9658);
and and5500(N9653,in2,N9659);
and and5501(N9654,N9660,R2);
and and5507(N9666,N9670,N9671);
and and5508(N9667,N9672,in1);
and and5509(N9668,N9673,R0);
and and5510(N9669,R2,N9674);
and and5516(N9681,N9685,N9686);
and and5517(N9682,N9687,N9688);
and and5518(N9683,N9689,R0);
and and5519(N9684,N9690,N9691);
and and5525(N9696,N9700,N9701);
and and5526(N9697,N9702,N9703);
and and5527(N9698,R0,N9704);
and and5528(N9699,N9705,R3);
and and5534(N9711,N9715,N9716);
and and5535(N9712,N9717,in1);
and and5536(N9713,N9718,N9719);
and and5537(N9714,R1,R3);
and and5543(N9726,N9730,N9731);
and and5544(N9727,N9732,in1);
and and5545(N9728,in2,N9733);
and and5546(N9729,N9734,R3);
and and5552(N9741,N9745,N9746);
and and5553(N9742,N9747,in2);
and and5554(N9743,N9748,N9749);
and and5555(N9744,R2,N9750);
and and5561(N9755,N9759,N9760);
and and5562(N9756,in1,N9761);
and and5563(N9757,N9762,N9763);
and and5564(N9758,R2,N9764);
and and5570(N9769,N9773,N9774);
and and5571(N9770,N9775,N9776);
and and5572(N9771,N9777,N9778);
and and5573(N9772,R2,R3);
and and5579(N9783,N9787,N9788);
and and5580(N9784,N9789,N9790);
and and5581(N9785,N9791,R0);
and and5582(N9786,N9792,R2);
and and5588(N9797,N9801,N9802);
and and5589(N9798,N9803,in1);
and and5590(N9799,in2,N9804);
and and5591(N9800,R1,R2);
and and5597(N9811,N9815,N9816);
and and5598(N9812,N9817,N9818);
and and5599(N9813,in2,R0);
and and5600(N9814,R1,R2);
and and5606(N9825,N9829,N9830);
and and5607(N9826,in1,N9831);
and and5608(N9827,R0,R1);
and and5609(N9828,R2,N9832);
and and5615(N9839,N9843,N9844);
and and5616(N9840,N9845,in1);
and and5617(N9841,N9846,N9847);
and and5618(N9842,R1,R2);
and and5624(N9853,N9857,N9858);
and and5625(N9854,in1,in2);
and and5626(N9855,N9859,N9860);
and and5627(N9856,R2,N9861);
and and5633(N9867,N9871,N9872);
and and5634(N9868,in0,in1);
and and5635(N9869,N9873,N9874);
and and5636(N9870,R2,N9875);
and and5642(N9881,N9885,N9886);
and and5643(N9882,in0,N9887);
and and5644(N9883,in2,R0);
and and5645(N9884,R1,N9888);
and and5651(N9895,N9899,N9900);
and and5652(N9896,in0,in1);
and and5653(N9897,N9901,R0);
and and5654(N9898,R1,N9902);
and and5660(N9909,N9913,N9914);
and and5661(N9910,in0,in1);
and and5662(N9911,in2,N9915);
and and5663(N9912,N9916,R2);
and and5669(N9923,N9927,N9928);
and and5670(N9924,N9929,N9930);
and and5671(N9925,N9931,N9932);
and and5672(N9926,R2,N9933);
and and5678(N9937,N9941,N9942);
and and5679(N9938,in1,in2);
and and5680(N9939,N9943,R1);
and and5681(N9940,N9944,R3);
and and5687(N9951,N9955,N9956);
and and5688(N9952,in1,N9957);
and and5689(N9953,N9958,R1);
and and5690(N9954,R2,N9959);
and and5696(N9965,N9969,N9970);
and and5697(N9966,in1,in2);
and and5698(N9967,N9971,N9972);
and and5699(N9968,R2,N9973);
and and5705(N9979,N9983,N9984);
and and5706(N9980,N9985,N9986);
and and5707(N9981,in2,R0);
and and5708(N9982,N9987,R2);
and and5714(N9993,N9997,N9998);
and and5715(N9994,N9999,in1);
and and5716(N9995,in2,R0);
and and5717(N9996,N10000,N10001);
and and5723(N10007,N10011,N10012);
and and5724(N10008,N10013,in1);
and and5725(N10009,R0,R1);
and and5726(N10010,N10014,N10015);
and and5732(N10021,N10025,N10026);
and and5733(N10022,N10027,N10028);
and and5734(N10023,in2,R0);
and and5735(N10024,R1,N10029);
and and5741(N10035,N10039,N10040);
and and5742(N10036,N10041,N10042);
and and5743(N10037,N10043,R0);
and and5744(N10038,N10044,N10045);
and and5750(N10049,N10053,N10054);
and and5751(N10050,N10055,in1);
and and5752(N10051,N10056,R0);
and and5753(N10052,N10057,R2);
and and5759(N10063,N10067,N10068);
and and5760(N10064,N10069,N10070);
and and5761(N10065,in2,R0);
and and5762(N10066,R2,R3);
and and5768(N10077,N10081,N10082);
and and5769(N10078,in0,in1);
and and5770(N10079,in2,N10083);
and and5771(N10080,N10084,N10085);
and and5777(N10091,N10095,N10096);
and and5778(N10092,N10097,in1);
and and5779(N10093,in2,R0);
and and5780(N10094,N10098,R3);
and and5786(N10105,N10109,N10110);
and and5787(N10106,N10111,N10112);
and and5788(N10107,in2,R0);
and and5789(N10108,R1,R2);
and and5795(N10119,N10123,N10124);
and and5796(N10120,N10125,in1);
and and5797(N10121,N10126,R0);
and and5798(N10122,R1,R2);
and and5804(N10133,N10137,N10138);
and and5805(N10134,N10139,in1);
and and5806(N10135,in2,R0);
and and5807(N10136,N10140,N10141);
and and5813(N10147,N10151,N10152);
and and5814(N10148,N10153,in1);
and and5815(N10149,N10154,N10155);
and and5816(N10150,R2,N10156);
and and5822(N10161,N10165,N10166);
and and5823(N10162,N10167,in2);
and and5824(N10163,R0,R1);
and and5825(N10164,N10168,N10169);
and and5831(N10175,N10179,N10180);
and and5832(N10176,in0,in1);
and and5833(N10177,in2,N10181);
and and5834(N10178,N10182,N10183);
and and5840(N10189,N10193,N10194);
and and5841(N10190,N10195,in1);
and and5842(N10191,N10196,R0);
and and5843(N10192,N10197,N10198);
and and5849(N10203,N10207,N10208);
and and5850(N10204,N10209,in1);
and and5851(N10205,N10210,R0);
and and5852(N10206,R1,N10211);
and and5858(N10217,N10221,N10222);
and and5859(N10218,N10223,N10224);
and and5860(N10219,in2,N10225);
and and5861(N10220,R1,N10226);
and and5867(N10231,N10235,N10236);
and and5868(N10232,in0,in1);
and and5869(N10233,N10237,N10238);
and and5870(N10234,R1,N10239);
and and5876(N10245,N10249,N10250);
and and5877(N10246,in0,N10251);
and and5878(N10247,in2,N10252);
and and5879(N10248,R2,N10253);
and and5885(N10259,N10263,N10264);
and and5886(N10260,in0,in1);
and and5887(N10261,N10265,N10266);
and and5888(N10262,N10267,R2);
and and5894(N10273,N10277,N10278);
and and5895(N10274,N10279,N10280);
and and5896(N10275,in2,N10281);
and and5897(N10276,R2,R3);
and and5903(N10287,N10291,N10292);
and and5904(N10288,N10293,in2);
and and5905(N10289,R0,R1);
and and5906(N10290,N10294,R3);
and and5912(N10301,N10305,N10306);
and and5913(N10302,N10307,N10308);
and and5914(N10303,in2,R0);
and and5915(N10304,R1,R2);
and and5921(N10314,N10318,N10319);
and and5922(N10315,in0,in1);
and and5923(N10316,N10320,R0);
and and5924(N10317,N10321,R2);
and and5930(N10327,N10331,N10332);
and and5931(N10328,N10333,N10334);
and and5932(N10329,in2,N10335);
and and5933(N10330,R1,R2);
and and5939(N10340,N10344,N10345);
and and5940(N10341,N10346,in1);
and and5941(N10342,N10347,N10348);
and and5942(N10343,R1,R2);
and and5948(N10353,N10357,N10358);
and and5949(N10354,N10359,in1);
and and5950(N10355,in2,R0);
and and5951(N10356,R1,R2);
and and5957(N10366,N10370,N10371);
and and5958(N10367,in1,N10372);
and and5959(N10368,N10373,N10374);
and and5960(N10369,R2,R3);
and and5966(N10379,N10383,N10384);
and and5967(N10380,in1,N10385);
and and5968(N10381,R0,N10386);
and and5969(N10382,R2,N10387);
and and5975(N10392,N10396,N10397);
and and5976(N10393,N10398,in1);
and and5977(N10394,in2,R0);
and and5978(N10395,N10399,R2);
and and5984(N10405,N10409,N10410);
and and5985(N10406,in0,in2);
and and5986(N10407,N10411,N10412);
and and5987(N10408,N10413,R3);
and and5993(N10418,N10422,N10423);
and and5994(N10419,in0,in1);
and and5995(N10420,N10424,N10425);
and and5996(N10421,N10426,R3);
and and6002(N10431,N10435,N10436);
and and6003(N10432,N10437,N10438);
and and6004(N10433,R0,R1);
and and6005(N10434,R2,N10439);
and and6011(N10444,N10448,N10449);
and and6012(N10445,N10450,N10451);
and and6013(N10446,N10452,R1);
and and6014(N10447,R2,R3);
and and6020(N10457,N10461,N10462);
and and6021(N10458,N10463,in1);
and and6022(N10459,N10464,R0);
and and6023(N10460,N10465,N10466);
and and6029(N10470,N10474,N10475);
and and6030(N10471,in0,N10476);
and and6031(N10472,N10477,R0);
and and6032(N10473,N10478,N10479);
and and6038(N10483,N10487,N10488);
and and6039(N10484,N10489,N10490);
and and6040(N10485,in2,R0);
and and6041(N10486,N10491,N10492);
and and6047(N10496,N10500,N10501);
and and6048(N10497,N10502,N10503);
and and6049(N10498,R0,R1);
and and6050(N10499,N10504,R3);
and and6056(N10509,N10513,N10514);
and and6057(N10510,in0,N10515);
and and6058(N10511,in2,R0);
and and6059(N10512,R2,N10516);
and and6065(N10522,N10526,N10527);
and and6066(N10523,in0,in1);
and and6067(N10524,R0,N10528);
and and6068(N10525,R2,N10529);
and and6074(N10535,N10539,N10540);
and and6075(N10536,N10541,in1);
and and6076(N10537,in2,R0);
and and6077(N10538,N10542,N10543);
and and6083(N10548,N10552,N10553);
and and6084(N10549,N10554,in1);
and and6085(N10550,N10555,R0);
and and6086(N10551,R1,R2);
and and6092(N10561,N10565,N10566);
and and6093(N10562,N10567,in1);
and and6094(N10563,N10568,R0);
and and6095(N10564,R1,R2);
and and6101(N10574,N10578,N10579);
and and6102(N10575,in0,N10580);
and and6103(N10576,R0,N10581);
and and6104(N10577,N10582,N10583);
and and6110(N10587,N10591,N10592);
and and6111(N10588,N10593,N10594);
and and6112(N10589,in2,R0);
and and6113(N10590,N10595,N10596);
and and6119(N10600,N10604,N10605);
and and6120(N10601,in1,in2);
and and6121(N10602,R0,N10606);
and and6122(N10603,R2,R3);
and and6128(N10613,N10617,N10618);
and and6129(N10614,in0,in1);
and and6130(N10615,in2,N10619);
and and6131(N10616,R2,R3);
and and6137(N10626,N10630,N10631);
and and6138(N10627,N10632,in1);
and and6139(N10628,in2,N10633);
and and6140(N10629,N10634,R3);
and and6146(N10639,N10643,N10644);
and and6147(N10640,in0,N10645);
and and6148(N10641,R0,N10646);
and and6149(N10642,N10647,R3);
and and6155(N10652,N10656,N10657);
and and6156(N10653,N10658,N10659);
and and6157(N10654,in2,N10660);
and and6158(N10655,N10661,R2);
and and6164(N10665,N10669,N10670);
and and6165(N10666,in0,in1);
and and6166(N10667,N10671,N10672);
and and6167(N10668,R1,R2);
and and6173(N10678,N10682,N10683);
and and6174(N10679,N10684,in1);
and and6175(N10680,in2,N10685);
and and6176(N10681,R1,R2);
and and6182(N10691,N10695,N10696);
and and6183(N10692,in0,N10697);
and and6184(N10693,in2,N10698);
and and6185(N10694,N10699,N10700);
and and6191(N10704,N10708,N10709);
and and6192(N10705,in0,in1);
and and6193(N10706,in2,R0);
and and6194(N10707,R2,N10710);
and and6200(N10717,N10721,N10722);
and and6201(N10718,in0,in1);
and and6202(N10719,R0,N10723);
and and6203(N10720,N10724,R3);
and and6209(N10730,N10734,N10735);
and and6210(N10731,in0,in2);
and and6211(N10732,R0,N10736);
and and6212(N10733,N10737,R3);
and and6218(N10743,N10747,N10748);
and and6219(N10744,N10749,in1);
and and6220(N10745,in2,R0);
and and6221(N10746,N10750,N10751);
and and6227(N10756,N10760,N10761);
and and6228(N10757,in0,in1);
and and6229(N10758,N10762,N10763);
and and6230(N10759,N10764,R2);
and and6236(N10769,N10773,N10774);
and and6237(N10770,N10775,in1);
and and6238(N10771,in2,N10776);
and and6239(N10772,N10777,R2);
and and6245(N10782,N10786,N10787);
and and6246(N10783,in1,N10788);
and and6247(N10784,R0,N10789);
and and6248(N10785,R2,N10790);
and and6254(N10795,N10799,N10800);
and and6255(N10796,in0,N10801);
and and6256(N10797,R0,N10802);
and and6257(N10798,R2,N10803);
and and6263(N10808,N10812,N10813);
and and6264(N10809,in0,in1);
and and6265(N10810,N10814,N10815);
and and6266(N10811,N10816,R2);
and and6272(N10821,N10825,N10826);
and and6273(N10822,in0,in1);
and and6274(N10823,in2,N10827);
and and6275(N10824,R2,R3);
and and6281(N10833,N10837,N10838);
and and6282(N10834,in0,in1);
and and6283(N10835,in2,N10839);
and and6284(N10836,R1,R2);
and and6290(N10845,N10849,N10850);
and and6291(N10846,in1,in2);
and and6292(N10847,R0,N10851);
and and6293(N10848,R2,N10852);
and and6299(N10857,N10861,N10862);
and and6300(N10858,in0,N10863);
and and6301(N10859,in2,N10864);
and and6302(N10860,R1,R2);
and and6308(N10869,N10873,N10874);
and and6309(N10870,N10875,N10876);
and and6310(N10871,in2,R0);
and and6311(N10872,R1,R2);
and and6317(N10881,N10885,N10886);
and and6318(N10882,in0,N10887);
and and6319(N10883,in2,R0);
and and6320(N10884,R1,R2);
and and6326(N10893,N10897,N10898);
and and6327(N10894,in0,N10899);
and and6328(N10895,in2,R0);
and and6329(N10896,R1,R2);
and and6335(N10905,N10909,N10910);
and and6336(N10906,in0,in1);
and and6337(N10907,in2,N10911);
and and6338(N10908,R1,R2);
and and6344(N10917,N10921,N10922);
and and6345(N10918,in1,in2);
and and6346(N10919,R0,R1);
and and6347(N10920,R2,R3);
and and6353(N10929,N10933,N10934);
and and6354(N10930,N10935,N10936);
and and6355(N10931,N10937,R1);
and and6356(N10932,R2,R3);
and and6362(N10941,N10945,N10946);
and and6363(N10942,in0,in1);
and and6364(N10943,in2,N10947);
and and6365(N10944,R1,R2);
and and6371(N10953,N10957,N10958);
and and6372(N10954,in0,N10959);
and and6373(N10955,N10960,R1);
and and6374(N10956,R2,N10961);
and and6380(N10965,N10969,N10970);
and and6381(N10966,N10971,in2);
and and6382(N10967,R0,R1);
and and6383(N10968,R2,R3);
and and6389(N10977,N10981,N10982);
and and6390(N10978,in0,N10983);
and and6391(N10979,in2,N10984);
and and6392(N10980,R1,R2);
and and6398(N10989,N10993,N10994);
and and6399(N10990,N10995,in1);
and and6400(N10991,in2,R0);
and and6401(N10992,R1,R2);
and and6407(N11001,N11005,N11006);
and and6408(N11002,in0,N11007);
and and6409(N11003,in2,N11008);
and and6410(N11004,R1,R2);
and and6416(N11013,N11017,N11018);
and and6417(N11014,in0,in2);
and and6418(N11015,R0,N11019);
and and6419(N11016,R2,N11020);
and and6425(N11025,N11029,N11030);
and and6426(N11026,in0,in1);
and and6427(N11027,N11031,R0);
and and6428(N11028,R1,R2);
and and6434(N11037,N11041,N11042);
and and6435(N11038,in0,N11043);
and and6436(N11039,in2,N11044);
and and6437(N11040,R1,R3);
and and6443(N11049,N11053,N11054);
and and6444(N11050,in0,in1);
and and6445(N11051,in2,R0);
and and6446(N11052,R1,R2);
and and6452(N11061,N11065,N11066);
and and6453(N11062,N11067,in2);
and and6454(N11063,R0,R1);
and and6455(N11064,R2,N11068);
and and6461(N11073,N11077,N11078);
and and6462(N11074,in0,N11079);
and and6463(N11075,in2,R1);
and and6464(N11076,R2,N11080);
and and6470(N11085,N11089,N11090);
and and6471(N11086,in0,in1);
and and6472(N11087,in2,N11091);
and and6473(N11088,N11092,R2);
and and6479(N11097,N11101,N11102);
and and6480(N11098,in1,in2);
and and6481(N11099,R0,R1);
and and6482(N11100,R2,N11103);
and and6488(N11109,N11113,N11114);
and and6489(N11110,in0,in1);
and and6490(N11111,N11115,R0);
and and6491(N11112,R1,R2);
and and6497(N11121,N11125,N11126);
and and6498(N11122,in0,in1);
and and6499(N11123,in2,R0);
and and6500(N11124,R1,N11127);
and and6506(N11133,N11137,N11138);
and and6507(N11134,in0,N11139);
and and6508(N11135,in2,R0);
and and6509(N11136,R1,N11140);
and and6515(N11145,N11149,N11150);
and and6516(N11146,in0,in1);
and and6517(N11147,N11151,R1);
and and6518(N11148,R2,R3);
and and6524(N11156,N11160,N11161);
and and6525(N11157,in1,in2);
and and6526(N11158,R0,N11162);
and and6527(N11159,N11163,R3);
and and6533(N11167,N11171,N11172);
and and6534(N11168,in0,N11173);
and and6535(N11169,in2,R0);
and and6536(N11170,N11174,R3);
and and6542(N11178,N11182,N11183);
and and6543(N11179,N11184,in1);
and and6544(N11180,in2,N11185);
and and6545(N11181,R2,R3);
and and6551(N11189,N11193,N11194);
and and6552(N11190,in1,in2);
and and6553(N11191,R0,R1);
and and6554(N11192,R2,N11195);
and and6560(N11200,N11204,N11205);
and and6561(N11201,in0,N11206);
and and6562(N11202,in2,R0);
and and6563(N11203,R1,R2);
and and6569(N11211,N11215,N11216);
and and6570(N11212,in0,in1);
and and6571(N11213,N11217,R0);
and and6572(N11214,R1,R2);
and and6578(N11222,N11226,N11227);
and and6579(N11223,in0,in1);
and and6580(N11224,in2,R0);
and and6581(N11225,N11228,R3);
and and6587(N11233,N11237,N11238);
and and6588(N11234,in1,in2);
and and6589(N11235,R0,R1);
and and6590(N11236,N11239,R3);
and and6596(N11244,N11248,N11249);
and and6597(N11245,in0,N11250);
and and6598(N11246,in2,R0);
and and6599(N11247,R1,R3);
and and6605(N11255,N11259,N11260);
and and6606(N11256,in0,in1);
and and6607(N11257,in2,R0);
and and6608(N11258,R1,R2);
and and6614(N11266,N11270,N11271);
and and6615(N11267,in0,in1);
and and6616(N11268,in2,R0);
and and6617(N11269,N11272,N11273);
and and6623(N11277,N11281,N11282);
and and6624(N11278,in0,N11283);
and and6625(N11279,R0,R1);
and and6626(N11280,R2,R3);
and and6632(N11288,N11292,N11293);
and and6633(N11289,in0,in1);
and and6634(N11290,in2,R0);
and and6635(N11291,N11294,R3);
and and6641(N11299,N11303,N11304);
and and6642(N11300,in0,in1);
and and6643(N11301,in2,R0);
and and6644(N11302,N11305,R2);
and and6650(N11310,N11314,N11315);
and and6651(N11311,in0,in1);
and and6652(N11312,N11316,R0);
and and6653(N11313,R1,R2);
and and6659(N11321,N11325,N11326);
and and6660(N11322,in0,in2);
and and6661(N11323,N11327,R1);
and and6662(N11324,R2,R3);
and and6668(N11331,N11335,N11336);
and and6669(N11332,in0,in1);
and and6670(N11333,in2,R1);
and and6671(N11334,R2,N11337);
and and6677(N11341,N11345,N11346);
and and6678(N11342,in0,in1);
and and6679(N11343,in2,R0);
and and6680(N11344,R1,R2);
and and6686(N11351,N11355,N11356);
and and6687(N11352,N11357,in2);
and and6688(N11353,R0,R1);
and and6689(N11354,R2,R3);
and and6695(N11361,N11365,N11366);
and and6696(N11362,in0,in2);
and and6697(N11363,R0,N11367);
and and6698(N11364,R2,R3);
and and6704(N11371,N11375,N11376);
and and6705(N11372,N11377,N11378);
and and6706(N11373,N11379,R1);
and and6707(N11374,N11380,N11381);
and and6712(N11387,N11391,N11392);
and and6713(N11388,N11393,N11394);
and and6714(N11389,N11395,N11396);
and and6715(N11390,N11397,N11398);
and and6720(N11403,N11407,in0);
and and6721(N11404,N11408,N11409);
and and6722(N11405,N11410,N11411);
and and6723(N11406,N11412,N11413);
and and6728(N11419,N11423,N11424);
and and6729(N11420,in2,N11425);
and and6730(N11421,N11426,N11427);
and and6731(N11422,N11428,N11429);
and and6736(N11435,N11439,N11440);
and and6737(N11436,N11441,N11442);
and and6738(N11437,R2,N11443);
and and6739(N11438,N11444,N11445);
and and6744(N11451,N11455,N11456);
and and6745(N11452,N11457,N11458);
and and6746(N11453,N11459,R3);
and and6747(N11454,N11460,N11461);
and and6752(N11467,N11471,N11472);
and and6753(N11468,N11473,N11474);
and and6754(N11469,N11475,N11476);
and and6755(N11470,N11477,N11478);
and and6760(N11483,N11487,in0);
and and6761(N11484,N11488,N11489);
and and6762(N11485,N11490,N11491);
and and6763(N11486,R4,N11492);
and and6768(N11498,N11502,N11503);
and and6769(N11499,N11504,R0);
and and6770(N11500,N11505,R2);
and and6771(N11501,N11506,N11507);
and and6776(N11513,N11517,N11518);
and and6777(N11514,N11519,N11520);
and and6778(N11515,N11521,N11522);
and and6779(N11516,R3,R4);
and and6784(N11528,N11532,N11533);
and and6785(N11529,N11534,N11535);
and and6786(N11530,N11536,N11537);
and and6787(N11531,R3,N11538);
and and6792(N11543,N11547,N11548);
and and6793(N11544,N11549,N11550);
and and6794(N11545,N11551,N11552);
and and6795(N11546,R3,N11553);
and and6800(N11558,N11562,N11563);
and and6801(N11559,N11564,R0);
and and6802(N11560,N11565,N11566);
and and6803(N11561,N11567,N11568);
and and6808(N11573,N11577,in2);
and and6809(N11574,N11578,N11579);
and and6810(N11575,N11580,R3);
and and6811(N11576,N11581,N11582);
and and6816(N11588,N11592,N11593);
and and6817(N11589,in1,N11594);
and and6818(N11590,R1,N11595);
and and6819(N11591,N11596,N11597);
and and6824(N11602,N11606,in0);
and and6825(N11603,in1,N11607);
and and6826(N11604,N11608,N11609);
and and6827(N11605,N11610,N11611);
and and6832(N11616,N11620,N11621);
and and6833(N11617,in1,in2);
and and6834(N11618,N11622,N11623);
and and6835(N11619,N11624,N11625);
and and6840(N11630,N11634,in1);
and and6841(N11631,in2,N11635);
and and6842(N11632,N11636,N11637);
and and6843(N11633,R4,N11638);
and and6848(N11644,N11648,in0);
and and6849(N11645,N11649,in2);
and and6850(N11646,N11650,R2);
and and6851(N11647,N11651,N11652);
and and6856(N11658,N11662,in0);
and and6857(N11659,in1,N11663);
and and6858(N11660,N11664,N11665);
and and6859(N11661,N11666,N11667);
and and6864(N11672,N11676,N11677);
and and6865(N11673,N11678,in2);
and and6866(N11674,N11679,R2);
and and6867(N11675,N11680,N11681);
and and6872(N11686,N11690,in0);
and and6873(N11687,N11691,N11692);
and and6874(N11688,N11693,R2);
and and6875(N11689,N11694,N11695);
and and6880(N11700,N11704,N11705);
and and6881(N11701,in2,R1);
and and6882(N11702,R2,N11706);
and and6883(N11703,N11707,N11708);
and and6888(N11714,N11718,N11719);
and and6889(N11715,N11720,in2);
and and6890(N11716,R0,N11721);
and and6891(N11717,R3,N11722);
and and6896(N11728,N11732,in0);
and and6897(N11729,N11733,N11734);
and and6898(N11730,R2,R3);
and and6899(N11731,N11735,N11736);
and and6904(N11742,N11746,N11747);
and and6905(N11743,in2,N11748);
and and6906(N11744,R2,R3);
and and6907(N11745,N11749,N11750);
and and6912(N11756,N11760,in0);
and and6913(N11757,N11761,N11762);
and and6914(N11758,N11763,R2);
and and6915(N11759,N11764,R5);
and and6920(N11770,N11774,N11775);
and and6921(N11771,in1,N11776);
and and6922(N11772,N11777,R2);
and and6923(N11773,N11778,N11779);
and and6928(N11784,N11788,N11789);
and and6929(N11785,N11790,N11791);
and and6930(N11786,R1,N11792);
and and6931(N11787,R3,R4);
and and6936(N11798,N11802,in0);
and and6937(N11799,in2,N11803);
and and6938(N11800,N11804,N11805);
and and6939(N11801,N11806,N11807);
and and6944(N11812,N11816,in0);
and and6945(N11813,in1,N11817);
and and6946(N11814,N11818,N11819);
and and6947(N11815,N11820,N11821);
and and6952(N11826,N11830,N11831);
and and6953(N11827,N11832,in2);
and and6954(N11828,N11833,N11834);
and and6955(N11829,N11835,R5);
and and6960(N11840,N11844,in0);
and and6961(N11841,R0,N11845);
and and6962(N11842,N11846,N11847);
and and6963(N11843,N11848,N11849);
and and6968(N11854,N11858,in0);
and and6969(N11855,N11859,N11860);
and and6970(N11856,N11861,N11862);
and and6971(N11857,R3,R4);
and and6976(N11868,N11872,in1);
and and6977(N11869,N11873,N11874);
and and6978(N11870,N11875,N11876);
and and6979(N11871,N11877,R4);
and and6984(N11882,N11886,N11887);
and and6985(N11883,N11888,R0);
and and6986(N11884,N11889,R3);
and and6987(N11885,R4,N11890);
and and6992(N11896,N11900,N11901);
and and6993(N11897,N11902,N11903);
and and6994(N11898,R1,R3);
and and6995(N11899,N11904,N11905);
and and7000(N11910,N11914,N11915);
and and7001(N11911,N11916,N11917);
and and7002(N11912,N11918,R3);
and and7003(N11913,R4,N11919);
and and7008(N11924,N11928,N11929);
and and7009(N11925,N11930,R0);
and and7010(N11926,N11931,N11932);
and and7011(N11927,R4,R5);
and and7016(N11938,N11942,N11943);
and and7017(N11939,N11944,in2);
and and7018(N11940,N11945,R3);
and and7019(N11941,N11946,N11947);
and and7024(N11952,N11956,N11957);
and and7025(N11953,in2,N11958);
and and7026(N11954,N11959,R3);
and and7027(N11955,N11960,N11961);
and and7032(N11966,N11970,N11971);
and and7033(N11967,N11972,N11973);
and and7034(N11968,N11974,R2);
and and7035(N11969,N11975,R4);
and and7040(N11980,N11984,in0);
and and7041(N11981,N11985,N11986);
and and7042(N11982,R2,N11987);
and and7043(N11983,R4,N11988);
and and7048(N11994,N11998,in0);
and and7049(N11995,N11999,in2);
and and7050(N11996,N12000,N12001);
and and7051(N11997,R2,N12002);
and and7056(N12008,N12012,in0);
and and7057(N12009,N12013,N12014);
and and7058(N12010,N12015,N12016);
and and7059(N12011,N12017,R3);
and and7064(N12022,N12026,N12027);
and and7065(N12023,in1,N12028);
and and7066(N12024,N12029,N12030);
and and7067(N12025,R3,N12031);
and and7072(N12036,N12040,N12041);
and and7073(N12037,in1,N12042);
and and7074(N12038,N12043,N12044);
and and7075(N12039,N12045,R4);
and and7080(N12050,N12054,N12055);
and and7081(N12051,N12056,N12057);
and and7082(N12052,N12058,R1);
and and7083(N12053,R2,R5);
and and7088(N12064,N12068,N12069);
and and7089(N12065,N12070,N12071);
and and7090(N12066,R1,R3);
and and7091(N12067,N12072,N12073);
and and7096(N12078,N12082,in0);
and and7097(N12079,N12083,R0);
and and7098(N12080,R1,R2);
and and7099(N12081,N12084,N12085);
and and7104(N12091,N12095,in1);
and and7105(N12092,in2,N12096);
and and7106(N12093,N12097,R2);
and and7107(N12094,N12098,N12099);
and and7112(N12104,N12108,N12109);
and and7113(N12105,N12110,N12111);
and and7114(N12106,N12112,R1);
and and7115(N12107,R3,R5);
and and7120(N12117,N12121,in0);
and and7121(N12118,N12122,N12123);
and and7122(N12119,N12124,R3);
and and7123(N12120,R4,N12125);
and and7128(N12130,N12134,in0);
and and7129(N12131,in2,N12135);
and and7130(N12132,N12136,R2);
and and7131(N12133,N12137,N12138);
and and7136(N12143,N12147,N12148);
and and7137(N12144,N12149,R1);
and and7138(N12145,R2,N12150);
and and7139(N12146,N12151,R5);
and and7144(N12156,N12160,N12161);
and and7145(N12157,in2,N12162);
and and7146(N12158,N12163,N12164);
and and7147(N12159,R3,R5);
and and7152(N12169,N12173,in0);
and and7153(N12170,N12174,R0);
and and7154(N12171,R1,N12175);
and and7155(N12172,R4,N12176);
and and7160(N12182,N12186,in0);
and and7161(N12183,N12187,N12188);
and and7162(N12184,R1,N12189);
and and7163(N12185,N12190,R5);
and and7168(N12195,N12199,in0);
and and7169(N12196,N12200,N12201);
and and7170(N12197,R1,R3);
and and7171(N12198,R4,N12202);
and and7176(N12208,N12212,N12213);
and and7177(N12209,in1,N12214);
and and7178(N12210,N12215,R3);
and and7179(N12211,N12216,R5);
and and7184(N12221,N12225,in0);
and and7185(N12222,N12226,N12227);
and and7186(N12223,R2,N12228);
and and7187(N12224,N12229,N12230);
and and7192(N12234,N12238,in0);
and and7193(N12235,N12239,N12240);
and and7194(N12236,R0,N12241);
and and7195(N12237,R2,R5);
and and7200(N12247,N12251,N12252);
and and7201(N12248,in1,R0);
and and7202(N12249,N12253,N12254);
and and7203(N12250,N12255,R5);
and and7208(N12260,N12264,N12265);
and and7209(N12261,in2,R0);
and and7210(N12262,N12266,N12267);
and and7211(N12263,R4,N12268);
and and7216(N12273,N12277,in0);
and and7217(N12274,N12278,R0);
and and7218(N12275,N12279,N12280);
and and7219(N12276,R4,N12281);
and and7224(N12286,N12290,in1);
and and7225(N12287,in2,N12291);
and and7226(N12288,N12292,N12293);
and and7227(N12289,R3,R4);
and and7232(N12299,N12303,in0);
and and7233(N12300,in1,N12304);
and and7234(N12301,N12305,N12306);
and and7235(N12302,R3,R4);
and and7240(N12312,N12316,in0);
and and7241(N12313,N12317,N12318);
and and7242(N12314,N12319,N12320);
and and7243(N12315,R2,R3);
and and7248(N12325,N12329,in0);
and and7249(N12326,N12330,R0);
and and7250(N12327,N12331,R2);
and and7251(N12328,N12332,R4);
and and7256(N12338,N12342,in0);
and and7257(N12339,N12343,N12344);
and and7258(N12340,R1,N12345);
and and7259(N12341,R3,N12346);
and and7264(N12351,N12355,in0);
and and7265(N12352,in1,N12356);
and and7266(N12353,R1,N12357);
and and7267(N12354,N12358,R5);
and and7272(N12364,N12368,N12369);
and and7273(N12365,in1,R0);
and and7274(N12366,R1,N12370);
and and7275(N12367,N12371,R5);
and and7280(N12377,N12381,in0);
and and7281(N12378,N12382,in2);
and and7282(N12379,N12383,R3);
and and7283(N12380,N12384,N12385);
and and7288(N12390,N12394,in0);
and and7289(N12391,N12395,in2);
and and7290(N12392,N12396,N12397);
and and7291(N12393,R2,N12398);
and and7296(N12403,N12407,N12408);
and and7297(N12404,N12409,N12410);
and and7298(N12405,N12411,R3);
and and7299(N12406,R4,R5);
and and7304(N12416,N12420,in0);
and and7305(N12417,N12421,R0);
and and7306(N12418,N12422,R2);
and and7307(N12419,N12423,N12424);
and and7312(N12429,N12433,in0);
and and7313(N12430,N12434,N12435);
and and7314(N12431,R0,N12436);
and and7315(N12432,R3,N12437);
and and7320(N12442,N12446,N12447);
and and7321(N12443,in2,N12448);
and and7322(N12444,R1,R3);
and and7323(N12445,N12449,N12450);
and and7328(N12455,N12459,in0);
and and7329(N12456,N12460,N12461);
and and7330(N12457,R1,R3);
and and7331(N12458,N12462,N12463);
and and7336(N12468,N12472,in0);
and and7337(N12469,N12473,N12474);
and and7338(N12470,N12475,N12476);
and and7339(N12471,R2,R4);
and and7344(N12481,N12485,in0);
and and7345(N12482,N12486,in2);
and and7346(N12483,R1,R2);
and and7347(N12484,N12487,N12488);
and and7352(N12494,N12498,N12499);
and and7353(N12495,in1,N12500);
and and7354(N12496,R1,R2);
and and7355(N12497,N12501,N12502);
and and7360(N12507,N12511,in1);
and and7361(N12508,in2,R0);
and and7362(N12509,N12512,N12513);
and and7363(N12510,N12514,N12515);
and and7368(N12520,N12524,in0);
and and7369(N12521,in2,N12525);
and and7370(N12522,N12526,N12527);
and and7371(N12523,N12528,R5);
and and7376(N12533,N12537,in0);
and and7377(N12534,N12538,N12539);
and and7378(N12535,R0,R2);
and and7379(N12536,N12540,R5);
and and7384(N12546,N12550,N12551);
and and7385(N12547,in1,N12552);
and and7386(N12548,N12553,R1);
and and7387(N12549,R2,N12554);
and and7392(N12559,N12563,in0);
and and7393(N12560,N12564,R0);
and and7394(N12561,N12565,R3);
and and7395(N12562,R4,N12566);
and and7400(N12572,N12576,in0);
and and7401(N12573,N12577,R0);
and and7402(N12574,N12578,R3);
and and7403(N12575,R4,N12579);
and and7408(N12585,N12589,in0);
and and7409(N12586,N12590,N12591);
and and7410(N12587,N12592,R3);
and and7411(N12588,R4,N12593);
and and7416(N12598,N12602,in0);
and and7417(N12599,in1,N12603);
and and7418(N12600,N12604,N12605);
and and7419(N12601,R3,N12606);
and and7424(N12611,N12615,in0);
and and7425(N12612,in1,N12616);
and and7426(N12613,R2,N12617);
and and7427(N12614,R4,N12618);
and and7432(N12624,N12628,in0);
and and7433(N12625,N12629,R0);
and and7434(N12626,N12630,R2);
and and7435(N12627,N12631,N12632);
and and7440(N12637,N12641,in0);
and and7441(N12638,N12642,N12643);
and and7442(N12639,R0,N12644);
and and7443(N12640,R3,N12645);
and and7448(N12650,N12654,N12655);
and and7449(N12651,N12656,in2);
and and7450(N12652,R0,N12657);
and and7451(N12653,R3,N12658);
and and7456(N12663,N12667,in0);
and and7457(N12664,N12668,R0);
and and7458(N12665,N12669,R3);
and and7459(N12666,N12670,N12671);
and and7464(N12676,N12680,in0);
and and7465(N12677,in1,in2);
and and7466(N12678,R1,R3);
and and7467(N12679,N12681,N12682);
and and7472(N12688,N12692,in0);
and and7473(N12689,in1,in2);
and and7474(N12690,R0,R1);
and and7475(N12691,N12693,N12694);
and and7480(N12700,N12704,N12705);
and and7481(N12701,in2,R0);
and and7482(N12702,R1,R2);
and and7483(N12703,N12706,N12707);
and and7488(N12712,N12716,in0);
and and7489(N12713,in1,in2);
and and7490(N12714,R0,N12717);
and and7491(N12715,N12718,N12719);
and and7496(N12724,N12728,in0);
and and7497(N12725,N12729,R1);
and and7498(N12726,R2,N12730);
and and7499(N12727,N12731,R5);
and and7504(N12736,N12740,N12741);
and and7505(N12737,in1,in2);
and and7506(N12738,R0,N12742);
and and7507(N12739,R2,N12743);
and and7512(N12748,N12752,in0);
and and7513(N12749,in1,in2);
and and7514(N12750,N12753,R2);
and and7515(N12751,N12754,R5);
and and7520(N12760,N12764,in0);
and and7521(N12761,N12765,in2);
and and7522(N12762,R1,N12766);
and and7523(N12763,R3,R4);
and and7528(N12772,N12776,in0);
and and7529(N12773,N12777,N12778);
and and7530(N12774,N12779,R1);
and and7531(N12775,R2,R4);
and and7536(N12784,N12788,N12789);
and and7537(N12785,N12790,in2);
and and7538(N12786,N12791,R1);
and and7539(N12787,R2,R4);
and and7544(N12796,N12800,N12801);
and and7545(N12797,N12802,in2);
and and7546(N12798,R0,N12803);
and and7547(N12799,R3,R4);
and and7552(N12808,N12812,N12813);
and and7553(N12809,N12814,N12815);
and and7554(N12810,R1,R2);
and and7555(N12811,N12816,R4);
and and7560(N12820,N12824,in0);
and and7561(N12821,N12825,in2);
and and7562(N12822,N12826,R2);
and and7563(N12823,N12827,N12828);
and and7568(N12832,N12836,N12837);
and and7569(N12833,N12838,N12839);
and and7570(N12834,R1,N12840);
and and7571(N12835,R3,R5);
and and7576(N12844,N12848,in1);
and and7577(N12845,N12849,R1);
and and7578(N12846,N12850,R3);
and and7579(N12847,N12851,R5);
and and7584(N12856,N12860,N12861);
and and7585(N12857,N12862,N12863);
and and7586(N12858,R1,R2);
and and7587(N12859,R3,R4);
and and7592(N12868,N12872,in0);
and and7593(N12869,in2,R0);
and and7594(N12870,N12873,R2);
and and7595(N12871,N12874,R5);
and and7600(N12880,N12884,in1);
and and7601(N12881,in2,R0);
and and7602(N12882,N12885,R2);
and and7603(N12883,N12886,R5);
and and7608(N12892,N12896,N12897);
and and7609(N12893,N12898,R0);
and and7610(N12894,N12899,R2);
and and7611(N12895,R4,R5);
and and7616(N12904,N12908,N12909);
and and7617(N12905,N12910,R0);
and and7618(N12906,R1,R2);
and and7619(N12907,N12911,N12912);
and and7624(N12916,N12920,N12921);
and and7625(N12917,in2,R1);
and and7626(N12918,N12922,R3);
and and7627(N12919,R4,R5);
and and7632(N12928,N12932,in0);
and and7633(N12929,N12933,N12934);
and and7634(N12930,R1,R3);
and and7635(N12931,R4,R5);
and and7640(N12940,N12944,in0);
and and7641(N12941,N12945,R0);
and and7642(N12942,N12946,N12947);
and and7643(N12943,R4,R5);
and and7648(N12952,N12956,in0);
and and7649(N12953,N12957,N12958);
and and7650(N12954,R0,R1);
and and7651(N12955,R2,N12959);
and and7656(N12964,N12968,in0);
and and7657(N12965,N12969,in2);
and and7658(N12966,R1,R2);
and and7659(N12967,R4,N12970);
and and7664(N12976,N12980,in0);
and and7665(N12977,N12981,N12982);
and and7666(N12978,R1,R2);
and and7667(N12979,R3,N12983);
and and7672(N12988,N12992,in0);
and and7673(N12989,in1,N12993);
and and7674(N12990,R0,R2);
and and7675(N12991,N12994,R4);
and and7680(N13000,N13004,in0);
and and7681(N13001,in2,R0);
and and7682(N13002,N13005,N13006);
and and7683(N13003,N13007,N13008);
and and7688(N13012,N13016,in0);
and and7689(N13013,N13017,N13018);
and and7690(N13014,N13019,R2);
and and7691(N13015,R4,N13020);
and and7696(N13024,N13028,in0);
and and7697(N13025,N13029,R0);
and and7698(N13026,R1,N13030);
and and7699(N13027,N13031,R4);
and and7704(N13036,N13040,in0);
and and7705(N13037,in1,R1);
and and7706(N13038,N13041,R3);
and and7707(N13039,N13042,N13043);
and and7712(N13048,N13052,in0);
and and7713(N13049,N13053,N13054);
and and7714(N13050,N13055,N13056);
and and7715(N13051,R3,R4);
and and7720(N13060,N13064,in1);
and and7721(N13061,N13065,N13066);
and and7722(N13062,N13067,N13068);
and and7723(N13063,R3,R4);
and and7728(N13072,N13076,in1);
and and7729(N13073,N13077,N13078);
and and7730(N13074,N13079,R2);
and and7731(N13075,R3,R4);
and and7736(N13084,N13088,in0);
and and7737(N13085,N13089,in2);
and and7738(N13086,R0,N13090);
and and7739(N13087,N13091,R4);
and and7744(N13096,N13100,in0);
and and7745(N13097,in1,N13101);
and and7746(N13098,R0,N13102);
and and7747(N13099,N13103,R4);
and and7752(N13108,N13112,in0);
and and7753(N13109,in2,R0);
and and7754(N13110,R1,N13113);
and and7755(N13111,N13114,R5);
and and7760(N13120,N13124,in1);
and and7761(N13121,in2,N13125);
and and7762(N13122,N13126,R2);
and and7763(N13123,N13127,R4);
and and7768(N13132,N13136,N13137);
and and7769(N13133,N13138,N13139);
and and7770(N13134,R2,R3);
and and7771(N13135,R4,R5);
and and7776(N13144,N13148,in0);
and and7777(N13145,N13149,N13150);
and and7778(N13146,N13151,R3);
and and7779(N13147,R4,R5);
and and7784(N13156,N13160,in1);
and and7785(N13157,N13161,N13162);
and and7786(N13158,N13163,R3);
and and7787(N13159,R4,R5);
and and7792(N13168,N13172,N13173);
and and7793(N13169,N13174,R0);
and and7794(N13170,R1,R2);
and and7795(N13171,R4,N13175);
and and7800(N13180,N13184,N13185);
and and7801(N13181,in2,R0);
and and7802(N13182,N13186,R3);
and and7803(N13183,N13187,R5);
and and7808(N13192,N13196,N13197);
and and7809(N13193,N13198,in2);
and and7810(N13194,R0,N13199);
and and7811(N13195,R2,R4);
and and7816(N13204,N13208,in0);
and and7817(N13205,N13209,N13210);
and and7818(N13206,R0,N13211);
and and7819(N13207,R2,N13212);
and and7824(N13216,N13220,N13221);
and and7825(N13217,in1,N13222);
and and7826(N13218,R0,N13223);
and and7827(N13219,R3,R5);
and and7832(N13228,N13232,in1);
and and7833(N13229,in2,R0);
and and7834(N13230,N13233,R3);
and and7835(N13231,N13234,N13235);
and and7840(N13240,N13244,in1);
and and7841(N13241,in2,R0);
and and7842(N13242,R1,R3);
and and7843(N13243,N13245,N13246);
and and7848(N13252,N13256,in0);
and and7849(N13253,N13257,N13258);
and and7850(N13254,R2,R3);
and and7851(N13255,N13259,N13260);
and and7856(N13264,N13268,in0);
and and7857(N13265,N13269,N13270);
and and7858(N13266,N13271,R2);
and and7859(N13267,R3,N13272);
and and7864(N13276,N13280,in0);
and and7865(N13277,N13281,R0);
and and7866(N13278,R1,N13282);
and and7867(N13279,R3,N13283);
and and7872(N13288,N13292,in0);
and and7873(N13289,in1,R0);
and and7874(N13290,R1,N13293);
and and7875(N13291,R4,N13294);
and and7880(N13300,N13304,N13305);
and and7881(N13301,N13306,N13307);
and and7882(N13302,R1,R2);
and and7883(N13303,R3,R4);
and and7888(N13312,N13316,in0);
and and7889(N13313,in1,in2);
and and7890(N13314,R0,N13317);
and and7891(N13315,N13318,R3);
and and7896(N13324,N13328,in0);
and and7897(N13325,N13329,R0);
and and7898(N13326,R1,N13330);
and and7899(N13327,N13331,R4);
and and7904(N13336,N13340,N13341);
and and7905(N13337,in1,R0);
and and7906(N13338,R1,N13342);
and and7907(N13339,N13343,R5);
and and7912(N13348,N13352,in0);
and and7913(N13349,N13353,N13354);
and and7914(N13350,N13355,R2);
and and7915(N13351,R3,R4);
and and7920(N13360,N13364,in0);
and and7921(N13361,N13365,in2);
and and7922(N13362,R0,N13366);
and and7923(N13363,N13367,N13368);
and and7928(N13372,N13376,in0);
and and7929(N13373,in1,N13377);
and and7930(N13374,N13378,R3);
and and7931(N13375,N13379,R5);
and and7936(N13384,N13388,N13389);
and and7937(N13385,in1,N13390);
and and7938(N13386,R0,R1);
and and7939(N13387,N13391,R5);
and and7944(N13396,N13400,in2);
and and7945(N13397,R0,N13401);
and and7946(N13398,R2,R3);
and and7947(N13399,R4,R5);
and and7952(N13407,N13411,in1);
and and7953(N13408,R0,N13412);
and and7954(N13409,R2,R3);
and and7955(N13410,R4,R5);
and and7960(N13418,N13422,in0);
and and7961(N13419,in2,N13423);
and and7962(N13420,N13424,R2);
and and7963(N13421,R3,R4);
and and7968(N13429,N13433,in0);
and and7969(N13430,N13434,R0);
and and7970(N13431,N13435,R2);
and and7971(N13432,R3,N13436);
and and7976(N13440,N13444,in0);
and and7977(N13441,in1,N13445);
and and7978(N13442,R1,R2);
and and7979(N13443,R4,R5);
and and7984(N13451,N13455,N13456);
and and7985(N13452,in1,in2);
and and7986(N13453,N13457,R1);
and and7987(N13454,R3,N13458);
and and7992(N13462,N13466,in1);
and and7993(N13463,N13467,R0);
and and7994(N13464,N13468,R2);
and and7995(N13465,R3,N13469);
and and8000(N13473,N13477,in0);
and and8001(N13474,in1,N13478);
and and8002(N13475,R1,R2);
and and8003(N13476,N13479,R5);
and and8008(N13484,N13488,in0);
and and8009(N13485,N13489,R0);
and and8010(N13486,R1,R3);
and and8011(N13487,R4,N13490);
and and8016(N13495,N13499,N13500);
and and8017(N13496,N13501,in2);
and and8018(N13497,R0,R1);
and and8019(N13498,R3,R4);
and and8024(N13506,N13510,in1);
and and8025(N13507,N13511,R0);
and and8026(N13508,R1,R3);
and and8027(N13509,R4,N13512);
and and8032(N13517,N13521,N13522);
and and8033(N13518,in2,R0);
and and8034(N13519,N13523,R3);
and and8035(N13520,R4,N13524);
and and8040(N13528,N13532,in0);
and and8041(N13529,N13533,R0);
and and8042(N13530,N13534,R3);
and and8043(N13531,R4,N13535);
and and8048(N13539,N13543,N13544);
and and8049(N13540,in2,N13545);
and and8050(N13541,R2,N13546);
and and8051(N13542,R4,R5);
and and8056(N13550,N13554,in0);
and and8057(N13551,in1,in2);
and and8058(N13552,R1,N13555);
and and8059(N13553,N13556,R5);
and and8064(N13561,N13565,in0);
and and8065(N13562,N13566,R0);
and and8066(N13563,N13567,R2);
and and8067(N13564,R3,R4);
and and8072(N13572,N13576,N13577);
and and8073(N13573,in1,N13578);
and and8074(N13574,R1,R3);
and and8075(N13575,N13579,R5);
and and8080(N13583,N13587,N13588);
and and8081(N13584,in2,N13589);
and and8082(N13585,R1,R3);
and and8083(N13586,N13590,R5);
and and8088(N13594,N13598,N13599);
and and8089(N13595,N13600,R0);
and and8090(N13596,R1,R3);
and and8091(N13597,R4,R5);
and and8096(N13605,N13609,N13610);
and and8097(N13606,in1,in2);
and and8098(N13607,N13611,R1);
and and8099(N13608,R3,N13612);
and and8104(N13616,N13620,in0);
and and8105(N13617,in2,R1);
and and8106(N13618,N13621,R3);
and and8107(N13619,N13622,R5);
and and8112(N13627,N13631,in0);
and and8113(N13628,in1,in2);
and and8114(N13629,N13632,R3);
and and8115(N13630,N13633,N13634);
and and8120(N13638,N13642,in0);
and and8121(N13639,N13643,R0);
and and8122(N13640,R1,R2);
and and8123(N13641,R3,R4);
and and8128(N13649,N13653,in0);
and and8129(N13650,in1,in2);
and and8130(N13651,R0,N13654);
and and8131(N13652,N13655,R4);
and and8136(N13660,N13664,in0);
and and8137(N13661,N13665,in2);
and and8138(N13662,R0,N13666);
and and8139(N13663,R2,R3);
and and8144(N13671,N13675,in0);
and and8145(N13672,in1,R1);
and and8146(N13673,R2,R3);
and and8147(N13674,N13676,R5);
and and8152(N13682,N13686,N13687);
and and8153(N13683,in1,in2);
and and8154(N13684,R1,R2);
and and8155(N13685,R3,R5);
and and8160(N13693,N13697,in0);
and and8161(N13694,in1,in2);
and and8162(N13695,R0,N13698);
and and8163(N13696,R2,N13699);
and and8168(N13704,N13708,in0);
and and8169(N13705,N13709,in2);
and and8170(N13706,R0,N13710);
and and8171(N13707,R3,N13711);
and and8176(N13715,N13719,in0);
and and8177(N13716,in1,N13720);
and and8178(N13717,R0,N13721);
and and8179(N13718,R3,N13722);
and and8184(N13726,N13730,in1);
and and8185(N13727,in2,N13731);
and and8186(N13728,N13732,R2);
and and8187(N13729,R4,N13733);
and and8192(N13737,N13741,in0);
and and8193(N13738,N13742,N13743);
and and8194(N13739,R1,R2);
and and8195(N13740,R4,R5);
and and8200(N13748,N13752,in1);
and and8201(N13749,in2,N13753);
and and8202(N13750,R2,R3);
and and8203(N13751,R4,N13754);
and and8208(N13759,N13763,in0);
and and8209(N13760,in1,N13764);
and and8210(N13761,N13765,R2);
and and8211(N13762,N13766,R5);
and and8216(N13770,N13774,in0);
and and8217(N13771,N13775,R0);
and and8218(N13772,R1,R2);
and and8219(N13773,N13776,R4);
and and8224(N13781,N13785,in0);
and and8225(N13782,N13786,in2);
and and8226(N13783,R0,R2);
and and8227(N13784,N13787,R4);
and and8232(N13792,N13796,in0);
and and8233(N13793,in1,N13797);
and and8234(N13794,R0,N13798);
and and8235(N13795,R2,R4);
and and8240(N13803,N13807,in0);
and and8241(N13804,in1,N13808);
and and8242(N13805,R1,R3);
and and8243(N13806,R4,N13809);
and and8248(N13814,N13818,in0);
and and8249(N13815,in1,in2);
and and8250(N13816,N13819,R1);
and and8251(N13817,R3,N13820);
and and8256(N13825,N13829,in0);
and and8257(N13826,in1,in2);
and and8258(N13827,N13830,N13831);
and and8259(N13828,R2,R4);
and and8264(N13836,N13840,in0);
and and8265(N13837,in1,in2);
and and8266(N13838,R0,R2);
and and8267(N13839,N13841,N13842);
and and8272(N13847,N13851,in0);
and and8273(N13848,in1,in2);
and and8274(N13849,R0,N13852);
and and8275(N13850,R2,N13853);
and and8280(N13858,N13862,in0);
and and8281(N13859,in1,in2);
and and8282(N13860,R0,N13863);
and and8283(N13861,N13864,R4);
and and8288(N13869,N13873,in0);
and and8289(N13870,in1,N13874);
and and8290(N13871,R0,N13875);
and and8291(N13872,N13876,R4);
and and8296(N13880,N13884,N13885);
and and8297(N13881,in1,N13886);
and and8298(N13882,R0,R1);
and and8299(N13883,R2,R4);
and and8304(N13891,N13895,in0);
and and8305(N13892,in1,in2);
and and8306(N13893,R0,R1);
and and8307(N13894,N13896,R5);
and and8312(N13902,N13906,in0);
and and8313(N13903,in1,N13907);
and and8314(N13904,N13908,N13909);
and and8315(N13905,R3,R4);
and and8320(N13913,N13917,in0);
and and8321(N13914,in1,N13918);
and and8322(N13915,R0,N13919);
and and8323(N13916,R3,R4);
and and8328(N13924,N13928,in0);
and and8329(N13925,in1,N13929);
and and8330(N13926,N13930,R3);
and and8331(N13927,R4,R5);
and and8336(N13935,N13939,in0);
and and8337(N13936,in2,N13940);
and and8338(N13937,N13941,R2);
and and8339(N13938,R3,N13942);
and and8344(N13946,N13950,in0);
and and8345(N13947,in1,in2);
and and8346(N13948,R0,R1);
and and8347(N13949,N13951,R5);
and and8352(N13957,N13961,in0);
and and8353(N13958,in1,R0);
and and8354(N13959,R1,R2);
and and8355(N13960,N13962,R5);
and and8360(N13967,N13971,in0);
and and8361(N13968,in1,in2);
and and8362(N13969,R1,R2);
and and8363(N13970,R3,R4);
and and8368(N13977,N13981,in0);
and and8369(N13978,N13982,R0);
and and8370(N13979,R1,R2);
and and8371(N13980,R3,N13983);
and and8376(N13987,N13991,in0);
and and8377(N13988,N13992,N13993);
and and8378(N13989,R2,R3);
and and8379(N13990,R4,R5);
and and8384(N13997,N14001,in0);
and and8385(N13998,N14002,R1);
and and8386(N13999,R2,R3);
and and8387(N14000,N14003,R5);
and and8392(N14007,N14011,in0);
and and8393(N14008,in1,N14012);
and and8394(N14009,N14013,R1);
and and8395(N14010,R2,R4);
and and8400(N14017,N14021,in0);
and and8401(N14018,in2,N14022);
and and8402(N14019,R1,N14023);
and and8403(N14020,R3,R5);
and and8408(N14027,N14031,in0);
and and8409(N14028,in1,N14032);
and and8410(N14029,R1,N14033);
and and8411(N14030,R3,R5);
and and8416(N14037,N14041,in1);
and and8417(N14038,in2,R0);
and and8418(N14039,R1,R2);
and and8419(N14040,R3,R4);
and and8424(N14047,N14051,in0);
and and8425(N14048,in2,R0);
and and8426(N14049,R1,R2);
and and8427(N14050,N14052,N14053);
and and8432(N14057,N14061,N14062);
and and8433(N14058,R0,R1);
and and8434(N14059,R2,R3);
and and8435(N14060,R4,R5);
and and8440(N14067,N14071,in0);
and and8441(N14068,R0,R1);
and and8442(N14069,R2,N14072);
and and8443(N14070,N14073,R5);
and and8448(N14077,N14081,N14082);
and and8449(N14078,N14083,R0);
and and8450(N14079,R2,R3);
and and8451(N14080,R4,R5);
and and8456(N14087,N14091,in1);
and and8457(N14088,in2,R0);
and and8458(N14089,N14092,R2);
and and8459(N14090,R3,R4);
and and8464(N14097,N14101,in0);
and and8465(N14098,in1,in2);
and and8466(N14099,R0,N14102);
and and8467(N14100,R3,R4);
and and8472(N14107,N14111,in1);
and and8473(N14108,in2,R1);
and and8474(N14109,R2,R3);
and and8475(N14110,R4,R5);
and and8480(N14117,N14121,in1);
and and8481(N14118,in2,R1);
and and8482(N14119,R2,R3);
and and8483(N14120,R4,N14122);
and and8488(N14126,N14130,in1);
and and8489(N14127,in2,R0);
and and8490(N14128,R2,R3);
and and8491(N14129,R4,N14131);
and and8496(N14135,N14139,in0);
and and8497(N14136,in1,N14140);
and and8498(N14137,R0,R2);
and and8499(N14138,R3,R4);
and and8504(N14144,N14148,in0);
and and8505(N14145,in1,in2);
and and8506(N14146,R0,R1);
and and8507(N14147,R3,R4);
and and8512(N14153,N14157,N14158);
and and8513(N14154,in1,R0);
and and8514(N14155,R1,R2);
and and8515(N14156,R3,R4);
and and8520(N14162,N14166,in0);
and and8521(N14163,in2,R0);
and and8522(N14164,R1,R3);
and and8523(N14165,R4,R5);
and and8528(N14171,N14175,in0);
and and8529(N14172,in1,R0);
and and8530(N14173,R1,R3);
and and8531(N14174,R4,R5);
and and8536(N14180,N14184,in0);
and and8537(N14181,in1,R0);
and and8538(N14182,R1,R2);
and and8539(N14183,R3,N14185);
and and8544(N14189,N14193,in2);
and and8545(N14190,R0,R1);
and and8546(N14191,R2,R3);
and and8547(N14192,R4,R5);
and and8552(N14198,N14202,in0);
and and8553(N14199,in1,N14203);
and and8554(N14200,R0,R1);
and and8555(N14201,R2,R3);
and and8560(N14207,R0,N14211);
and and8561(N14208,N14212,N14213);
and and8562(N14209,N14214,N14215);
and and8563(N14210,N14216,N14217);
and and8567(N14221,in1,N14225);
and and8568(N14222,N14226,N14227);
and and8569(N14223,N14228,N14229);
and and8570(N14224,N14230,N14231);
and and8574(N14235,N14239,R0);
and and8575(N14236,N14240,N14241);
and and8576(N14237,N14242,N14243);
and and8577(N14238,N14244,N14245);
and and8581(N14249,in1,N14253);
and and8582(N14250,N14254,N14255);
and and8583(N14251,N14256,N14257);
and and8584(N14252,N14258,N14259);
and and8588(N14263,in0,N14267);
and and8589(N14264,N14268,N14269);
and and8590(N14265,N14270,N14271);
and and8591(N14266,R5,N14272);
and and8595(N14276,N14280,R0);
and and8596(N14277,N14281,N14282);
and and8597(N14278,N14283,N14284);
and and8598(N14279,R5,N14285);
and and8602(N14289,N14293,N14294);
and and8603(N14290,N14295,R2);
and and8604(N14291,N14296,N14297);
and and8605(N14292,R6,N14298);
and and8609(N14302,N14306,N14307);
and and8610(N14303,R1,N14308);
and and8611(N14304,N14309,R5);
and and8612(N14305,N14310,N14311);
and and8616(N14315,N14319,N14320);
and and8617(N14316,N14321,N14322);
and and8618(N14317,R3,N14323);
and and8619(N14318,R6,N14324);
and and8623(N14328,in1,R0);
and and8624(N14329,N14332,N14333);
and and8625(N14330,N14334,N14335);
and and8626(N14331,N14336,N14337);
and and8630(N14341,in1,N14345);
and and8631(N14342,N14346,R3);
and and8632(N14343,N14347,N14348);
and and8633(N14344,N14349,N14350);
and and8637(N14354,in0,N14358);
and and8638(N14355,R1,R2);
and and8639(N14356,N14359,N14360);
and and8640(N14357,N14361,N14362);
and and8644(N14366,in0,R0);
and and8645(N14367,N14370,R2);
and and8646(N14368,N14371,N14372);
and and8647(N14369,N14373,N14374);
and and8651(N14378,N14382,N14383);
and and8652(N14379,R1,R2);
and and8653(N14380,N14384,R5);
and and8654(N14381,N14385,N14386);
and and8658(N14390,N14394,N14395);
and and8659(N14391,R0,R1);
and and8660(N14392,N14396,N14397);
and and8661(N14393,N14398,R7);
and and8665(N14402,in0,R0);
and and8666(N14403,N14406,N14407);
and and8667(N14404,R3,N14408);
and and8668(N14405,N14409,N14410);
and and8672(N14414,N14418,R0);
and and8673(N14415,N14419,N14420);
and and8674(N14416,N14421,N14422);
and and8675(N14417,R6,R7);
and and8679(N14426,in0,N14430);
and and8680(N14427,N14431,N14432);
and and8681(N14428,R3,N14433);
and and8682(N14429,N14434,R7);
and and8686(N14438,N14442,in2);
and and8687(N14439,R2,N14443);
and and8688(N14440,R4,N14444);
and and8689(N14441,N14445,N14446);
and and8693(N14450,N14454,in1);
and and8694(N14451,R2,N14455);
and and8695(N14452,R4,N14456);
and and8696(N14453,N14457,N14458);
and and8700(N14462,N14466,N14467);
and and8701(N14463,R0,R1);
and and8702(N14464,R3,N14468);
and and8703(N14465,N14469,N14470);
and and8707(N14474,in0,N14478);
and and8708(N14475,N14479,R3);
and and8709(N14476,N14480,R5);
and and8710(N14477,N14481,N14482);
and and8714(N14486,in2,N14490);
and and8715(N14487,R1,N14491);
and and8716(N14488,N14492,R5);
and and8717(N14489,N14493,N14494);
and and8721(N14498,in0,N14502);
and and8722(N14499,N14503,N14504);
and and8723(N14500,R3,N14505);
and and8724(N14501,N14506,R7);
and and8728(N14510,in0,R0);
and and8729(N14511,N14514,R2);
and and8730(N14512,N14515,N14516);
and and8731(N14513,N14517,R7);
and and8735(N14521,in0,R0);
and and8736(N14522,N14525,N14526);
and and8737(N14523,N14527,N14528);
and and8738(N14524,R5,R6);
and and8742(N14532,in0,R0);
and and8743(N14533,N14536,R3);
and and8744(N14534,N14537,N14538);
and and8745(N14535,N14539,R7);
and and8749(N14543,N14547,N14548);
and and8750(N14544,R2,N14549);
and and8751(N14545,N14550,R5);
and and8752(N14546,R6,R7);
and and8756(N14554,in0,N14558);
and and8757(N14555,N14559,R2);
and and8758(N14556,N14560,R4);
and and8759(N14557,R6,N14561);
and and8763(N14565,in0,N14569);
and and8764(N14566,N14570,R3);
and and8765(N14567,R4,N14571);
and and8766(N14568,N14572,R7);
and and8770(N14576,N14580,R0);
and and8771(N14577,R1,N14581);
and and8772(N14578,N14582,R5);
and and8773(N14579,N14583,R7);
and and8777(N14587,in0,N14591);
and and8778(N14588,R0,R1);
and and8779(N14589,R3,N14592);
and and8780(N14590,N14593,N14594);
and and8784(N14598,in0,N14602);
and and8785(N14599,R0,R1);
and and8786(N14600,R3,N14603);
and and8787(N14601,N14604,N14605);
and and8791(N14609,in1,R1);
and and8792(N14610,N14613,R3);
and and8793(N14611,R4,R5);
and and8794(N14612,N14614,N14615);
and and8798(N14619,N14623,R0);
and and8799(N14620,R1,N14624);
and and8800(N14621,R3,N14625);
and and8801(N14622,R6,R7);
and and8805(N14629,in2,N14633);
and and8806(N14630,N14634,R2);
and and8807(N14631,R3,R4);
and and8808(N14632,N14635,R7);
and and8812(N14639,in0,N14643);
and and8813(N14640,R2,R3);
and and8814(N14641,R4,N14644);
and and8815(N14642,R6,N14645);
and and8819(N14649,in0,R0);
and and8820(N14650,N14653,R3);
and and8821(N14651,R4,N14654);
and and8822(N14652,N14655,R7);
and and8826(N14659,N14663,R0);
and and8827(N14660,R1,N14664);
and and8828(N14661,R3,R5);
and and8829(N14662,R6,R7);
and and8833(N14668,in0,R0);
and and8834(N14669,N14672,R2);
and and8835(N14670,R3,R4);
and and8836(N14671,R6,N14673);
and and8840(N14677,R0,R1);
and and8841(N14678,R2,R3);
and and8842(N14679,N14681,R5);
and and8843(N14680,R6,N14682);
and and8847(N14686,in1,N14690);
and and8848(N14687,R1,R2);
and and8849(N14688,R4,R5);
and and8850(N14689,N14691,R7);
and and8854(N14695,in0,in2);
and and8855(N14696,N14699,R2);
and and8856(N14697,R3,R4);
and and8857(N14698,N14700,R7);
and and8861(N14704,in1,in2);
and and8862(N14705,R0,R1);
and and8863(N14706,R3,R5);
and and8864(N14707,R6,R7);
and and8868(N14711,N14714,N14715);
and and8869(N14712,N14716,R4);
and and8870(N14713,N14717,R7);
and and8874(N14721,R1,R2);
and and8875(N14722,R3,N14724);
and and8876(N14723,R6,N14725);
and and5061(N8892,N8900,R5);
and and5062(N8893,N8901,N8902);
and and5070(N8910,N8916,N8917);
and and5071(N8911,N8918,N8919);
and and5079(N8927,R3,N8934);
and and5080(N8928,N8935,N8936);
and and5088(N8944,N8951,N8952);
and and5089(N8945,N8953,R7);
and and5097(N8961,R4,R5);
and and5098(N8962,N8969,N8970);
and and5106(N8978,R4,N8985);
and and5107(N8979,N8986,N8987);
and and5115(N8995,N9000,N9001);
and and5116(N8996,N9002,N9003);
and and5124(N9011,N9016,N9017);
and and5125(N9012,N9018,N9019);
and and5133(N9027,N9034,R5);
and and5134(N9028,N9035,R7);
and and5142(N9043,R4,N9049);
and and5143(N9044,N9050,N9051);
and and5151(N9059,N9065,N9066);
and and5152(N9060,N9067,R7);
and and5160(N9075,N9080,N9081);
and and5161(N9076,N9082,N9083);
and and5169(N9091,N9097,R5);
and and5170(N9092,N9098,N9099);
and and5178(N9107,N9112,N9113);
and and5179(N9108,N9114,N9115);
and and5187(N9123,N9128,N9129);
and and5188(N9124,N9130,N9131);
and and5196(N9139,N9145,N9146);
and and5197(N9140,R5,N9147);
and and5205(N9155,N9161,N9162);
and and5206(N9156,R6,N9163);
and and5214(N9171,R4,N9178);
and and5215(N9172,R6,N9179);
and and5223(N9187,R3,R4);
and and5224(N9188,N9194,N9195);
and and5232(N9203,N9209,R5);
and and5233(N9204,N9210,N9211);
and and5241(N9219,N9226,R4);
and and5242(N9220,N9227,R7);
and and5250(N9235,R3,R5);
and and5251(N9236,N9241,N9242);
and and5259(N9250,R3,N9256);
and and5260(N9251,N9257,R7);
and and5268(N9265,N9270,R5);
and and5269(N9266,N9271,N9272);
and and5277(N9280,N9287,R5);
and and5278(N9281,R6,R7);
and and5286(N9295,N9301,R5);
and and5287(N9296,R6,N9302);
and and5295(N9310,N9316,R5);
and and5296(N9311,R6,N9317);
and and5304(N9325,R4,N9330);
and and5305(N9326,N9331,N9332);
and and5313(N9340,N9345,R5);
and and5314(N9341,N9346,N9347);
and and5322(N9355,N9360,R5);
and and5323(N9356,N9361,N9362);
and and5331(N9370,N9374,N9375);
and and5332(N9371,N9376,N9377);
and and5340(N9385,N9391,R5);
and and5341(N9386,N9392,R7);
and and5349(N9400,R4,R5);
and and5350(N9401,N9406,N9407);
and and5358(N9415,R3,R4);
and and5359(N9416,N9422,R7);
and and5367(N9430,N9436,R5);
and and5368(N9431,R6,N9437);
and and5376(N9445,N9451,N9452);
and and5377(N9446,R6,R7);
and and5385(N9460,N9466,N9467);
and and5386(N9461,R6,R7);
and and5394(N9475,N9480,R5);
and and5395(N9476,N9481,N9482);
and and5403(N9490,R4,N9496);
and and5404(N9491,N9497,R7);
and and5412(N9505,R3,N9511);
and and5413(N9506,N9512,R6);
and and5421(N9520,N9525,R4);
and and5422(N9521,N9526,N9527);
and and5430(N9535,R4,N9540);
and and5431(N9536,N9541,N9542);
and and5439(N9550,R3,R4);
and and5440(N9551,N9556,N9557);
and and5448(N9565,R4,N9570);
and and5449(N9566,N9571,N9572);
and and5457(N9580,N9586,N9587);
and and5458(N9581,R6,R7);
and and5466(N9595,R3,N9602);
and and5467(N9596,R6,R7);
and and5475(N9610,R4,N9616);
and and5476(N9611,R6,N9617);
and and5484(N9625,R4,R5);
and and5485(N9626,N9631,N9632);
and and5493(N9640,R3,N9646);
and and5494(N9641,N9647,R7);
and and5502(N9655,N9661,R4);
and and5503(N9656,N9662,R6);
and and5511(N9670,N9675,N9676);
and and5512(N9671,R6,N9677);
and and5520(N9685,R3,R5);
and and5521(N9686,R6,N9692);
and and5529(N9700,N9706,R5);
and and5530(N9701,N9707,R7);
and and5538(N9715,N9720,N9721);
and and5539(N9716,N9722,R7);
and and5547(N9730,N9735,R5);
and and5548(N9731,N9736,N9737);
and and5556(N9745,R4,R5);
and and5557(N9746,N9751,R7);
and and5565(N9759,R4,R5);
and and5566(N9760,N9765,R7);
and and5574(N9773,R4,N9779);
and and5575(N9774,R6,R7);
and and5583(N9787,R4,N9793);
and and5584(N9788,R6,R7);
and and5592(N9801,R3,N9805);
and and5593(N9802,N9806,N9807);
and and5601(N9815,N9819,N9820);
and and5602(N9816,N9821,R7);
and and5610(N9829,N9833,N9834);
and and5611(N9830,N9835,R7);
and and5619(N9843,R3,R4);
and and5620(N9844,N9848,N9849);
and and5628(N9857,N9862,R5);
and and5629(N9858,R6,N9863);
and and5637(N9871,N9876,R5);
and and5638(N9872,R6,N9877);
and and5646(N9885,N9889,N9890);
and and5647(N9886,N9891,R7);
and and5655(N9899,N9903,N9904);
and and5656(N9900,N9905,R7);
and and5664(N9913,R3,N9917);
and and5665(N9914,N9918,N9919);
and and5673(N9927,R4,R5);
and and5674(N9928,R6,R7);
and and5682(N9941,R4,N9945);
and and5683(N9942,N9946,N9947);
and and5691(N9955,R4,N9960);
and and5692(N9956,N9961,R7);
and and5700(N9969,N9974,N9975);
and and5701(N9970,R6,R7);
and and5709(N9983,N9988,R5);
and and5710(N9984,R6,N9989);
and and5718(N9997,R4,N10002);
and and5719(N9998,R6,N10003);
and and5727(N10011,R4,N10016);
and and5728(N10012,N10017,R7);
and and5736(N10025,R4,N10030);
and and5737(N10026,N10031,R7);
and and5745(N10039,R4,R5);
and and5746(N10040,R6,R7);
and and5754(N10053,R3,N10058);
and and5755(N10054,R6,N10059);
and and5763(N10067,N10071,N10072);
and and5764(N10068,R6,N10073);
and and5772(N10081,R4,R5);
and and5773(N10082,N10086,N10087);
and and5781(N10095,R4,N10099);
and and5782(N10096,N10100,N10101);
and and5790(N10109,R3,N10113);
and and5791(N10110,N10114,N10115);
and and5799(N10123,R3,N10127);
and and5800(N10124,N10128,N10129);
and and5808(N10137,R4,R5);
and and5809(N10138,N10142,N10143);
and and5817(N10151,N10157,R5);
and and5818(N10152,R6,R7);
and and5826(N10165,N10170,R5);
and and5827(N10166,N10171,R7);
and and5835(N10179,R3,N10184);
and and5836(N10180,N10185,R7);
and and5844(N10193,R3,N10199);
and and5845(N10194,R5,R6);
and and5853(N10207,R3,N10212);
and and5854(N10208,N10213,R7);
and and5862(N10221,R3,R4);
and and5863(N10222,N10227,R7);
and and5871(N10235,R3,N10240);
and and5872(N10236,N10241,R7);
and and5880(N10249,R4,N10254);
and and5881(N10250,N10255,R7);
and and5889(N10263,N10268,R4);
and and5890(N10264,N10269,R7);
and and5898(N10277,N10282,R5);
and and5899(N10278,R6,N10283);
and and5907(N10291,N10295,R5);
and and5908(N10292,N10296,N10297);
and and5916(N10305,R4,R5);
and and5917(N10306,N10309,N10310);
and and5925(N10318,R3,N10322);
and and5926(N10319,R5,N10323);
and and5934(N10331,R3,N10336);
and and5935(N10332,R6,R7);
and and5943(N10344,R3,N10349);
and and5944(N10345,R6,R7);
and and5952(N10357,N10360,N10361);
and and5953(N10358,R6,N10362);
and and5961(N10370,R4,N10375);
and and5962(N10371,R6,R7);
and and5970(N10383,R4,N10388);
and and5971(N10384,R6,R7);
and and5979(N10396,R3,N10400);
and and5980(N10397,N10401,R7);
and and5988(N10409,N10414,R5);
and and5989(N10410,R6,R7);
and and5997(N10422,N10427,R5);
and and5998(N10423,R6,R7);
and and6006(N10435,R4,R5);
and and6007(N10436,R6,N10440);
and and6015(N10448,N10453,R5);
and and6016(N10449,R6,R7);
and and6024(N10461,R3,R4);
and and6025(N10462,R6,R7);
and and6033(N10474,R3,R5);
and and6034(N10475,R6,R7);
and and6042(N10487,R3,R5);
and and6043(N10488,R6,R7);
and and6051(N10500,R4,R5);
and and6052(N10501,N10505,R7);
and and6060(N10513,R4,R5);
and and6061(N10514,N10517,N10518);
and and6069(N10526,R4,R5);
and and6070(N10527,N10530,N10531);
and and6078(N10539,R3,R4);
and and6079(N10540,N10544,R7);
and and6087(N10552,N10556,R4);
and and6088(N10553,R6,N10557);
and and6096(N10565,R3,R4);
and and6097(N10566,N10569,N10570);
and and6105(N10578,R4,R5);
and and6106(N10579,R6,R7);
and and6114(N10591,R4,R5);
and and6115(N10592,R6,R7);
and and6123(N10604,N10607,N10608);
and and6124(N10605,R6,N10609);
and and6132(N10617,R4,N10620);
and and6133(N10618,N10621,N10622);
and and6141(N10630,R4,R5);
and and6142(N10631,R6,N10635);
and and6150(N10643,R4,R5);
and and6151(N10644,N10648,R7);
and and6159(N10656,R3,R5);
and and6160(N10657,R6,R7);
and and6168(N10669,R3,N10673);
and and6169(N10670,N10674,R7);
and and6177(N10682,R3,N10686);
and and6178(N10683,N10687,R7);
and and6186(N10695,R3,R4);
and and6187(N10696,R5,R7);
and and6195(N10708,N10711,N10712);
and and6196(N10709,R6,N10713);
and and6204(N10721,N10725,R5);
and and6205(N10722,R6,N10726);
and and6213(N10734,N10738,R5);
and and6214(N10735,N10739,R7);
and and6222(N10747,R3,N10752);
and and6223(N10748,R5,R7);
and and6231(N10760,R3,N10765);
and and6232(N10761,R6,R7);
and and6240(N10773,R3,N10778);
and and6241(N10774,R6,R7);
and and6249(N10786,R4,R5);
and and6250(N10787,R6,N10791);
and and6258(N10799,R4,R5);
and and6259(N10800,R6,N10804);
and and6267(N10812,R3,R5);
and and6268(N10813,R6,N10817);
and and6276(N10825,N10828,R5);
and and6277(N10826,N10829,R7);
and and6285(N10837,N10840,N10841);
and and6286(N10838,R6,R7);
and and6294(N10849,N10853,R5);
and and6295(N10850,R6,R7);
and and6303(N10861,R3,R4);
and and6304(N10862,N10865,R7);
and and6312(N10873,R3,N10877);
and and6313(N10874,R5,R7);
and and6321(N10885,R3,R5);
and and6322(N10886,N10888,N10889);
and and6330(N10897,N10900,R5);
and and6331(N10898,N10901,R7);
and and6339(N10909,N10912,R5);
and and6340(N10910,R6,N10913);
and and6348(N10921,N10923,N10924);
and and6349(N10922,N10925,R7);
and and6357(N10933,R4,R5);
and and6358(N10934,R6,R7);
and and6366(N10945,N10948,R4);
and and6367(N10946,N10949,R7);
and and6375(N10957,R4,R5);
and and6376(N10958,R6,R7);
and and6384(N10969,R4,N10972);
and and6385(N10970,N10973,R7);
and and6393(N10981,N10985,R4);
and and6394(N10982,R6,R7);
and and6402(N10993,R4,N10996);
and and6403(N10994,R6,N10997);
and and6411(N11005,R3,R4);
and and6412(N11006,R5,N11009);
and and6420(N11017,R4,R5);
and and6421(N11018,N11021,R7);
and and6429(N11029,N11032,N11033);
and and6430(N11030,R6,R7);
and and6438(N11041,R4,R5);
and and6439(N11042,N11045,R7);
and and6447(N11053,N11055,R4);
and and6448(N11054,N11056,N11057);
and and6456(N11065,R4,N11069);
and and6457(N11066,R6,R7);
and and6465(N11077,R4,R5);
and and6466(N11078,N11081,R7);
and and6474(N11089,N11093,R5);
and and6475(N11090,R6,R7);
and and6483(N11101,R4,N11104);
and and6484(N11102,N11105,R7);
and and6492(N11113,N11116,R4);
and and6493(N11114,N11117,R7);
and and6501(N11125,R3,N11128);
and and6502(N11126,N11129,R7);
and and6510(N11137,R3,R5);
and and6511(N11138,N11141,R7);
and and6519(N11149,R4,R5);
and and6520(N11150,R6,N11152);
and and6528(N11160,R4,R5);
and and6529(N11161,R6,R7);
and and6537(N11171,R4,R5);
and and6538(N11172,R6,R7);
and and6546(N11182,R4,R5);
and and6547(N11183,R6,R7);
and and6555(N11193,R4,R5);
and and6556(N11194,R6,N11196);
and and6564(N11204,N11207,R4);
and and6565(N11205,R5,R6);
and and6573(N11215,N11218,R4);
and and6574(N11216,R5,R6);
and and6582(N11226,N11229,R5);
and and6583(N11227,R6,R7);
and and6591(N11237,R4,R5);
and and6592(N11238,N11240,R7);
and and6600(N11248,N11251,R5);
and and6601(N11249,R6,R7);
and and6609(N11259,N11261,R4);
and and6610(N11260,N11262,R6);
and and6618(N11270,R4,R5);
and and6619(N11271,R6,R7);
and and6627(N11281,R4,N11284);
and and6628(N11282,R6,R7);
and and6636(N11292,R4,R5);
and and6637(N11293,N11295,R7);
and and6645(N11303,N11306,R4);
and and6646(N11304,R5,R6);
and and6654(N11314,R3,N11317);
and and6655(N11315,R6,R7);
and and6663(N11325,R4,R5);
and and6664(N11326,R6,R7);
and and6672(N11335,R4,R5);
and and6673(N11336,R6,R7);
and and6681(N11345,N11347,R4);
and and6682(N11346,R5,R7);
and and6690(N11355,R4,R5);
and and6691(N11356,R6,R7);
and and6699(N11365,R4,R5);
and and6700(N11366,R6,R7);
and and6708(N11375,N11382,N11383);
and and6716(N11391,R6,N11399);
and and6724(N11407,N11414,N11415);
and and6732(N11423,N11430,N11431);
and and6740(N11439,N11446,N11447);
and and6748(N11455,N11462,N11463);
and and6756(N11471,N11479,R7);
and and6764(N11487,N11493,N11494);
and and6772(N11502,N11508,N11509);
and and6780(N11517,N11523,N11524);
and and6788(N11532,N11539,R7);
and and6796(N11547,R5,N11554);
and and6804(N11562,R5,N11569);
and and6812(N11577,N11583,N11584);
and and6820(N11592,N11598,R7);
and and6828(N11606,R6,N11612);
and and6836(N11620,R6,N11626);
and and6844(N11634,N11639,N11640);
and and6852(N11648,N11653,N11654);
and and6860(N11662,R5,N11668);
and and6868(N11676,N11682,R7);
and and6876(N11690,N11696,R7);
and and6884(N11704,N11709,N11710);
and and6892(N11718,N11723,N11724);
and and6900(N11732,N11737,N11738);
and and6908(N11746,N11751,N11752);
and and6916(N11760,N11765,N11766);
and and6924(N11774,R5,N11780);
and and6932(N11788,N11793,N11794);
and and6940(N11802,N11808,R7);
and and6948(N11816,N11822,R7);
and and6956(N11830,N11836,R7);
and and6964(N11844,R6,N11850);
and and6972(N11858,N11863,N11864);
and and6980(N11872,R5,N11878);
and and6988(N11886,N11891,N11892);
and and6996(N11900,R6,N11906);
and and7004(N11914,R6,N11920);
and and7012(N11928,N11933,N11934);
and and7020(N11942,R6,N11948);
and and7028(N11956,N11962,R7);
and and7036(N11970,R6,N11976);
and and7044(N11984,N11989,N11990);
and and7052(N11998,N12003,N12004);
and and7060(N12012,N12018,R6);
and and7068(N12026,N12032,R7);
and and7076(N12040,R5,N12046);
and and7084(N12054,N12059,N12060);
and and7092(N12068,R6,N12074);
and and7100(N12082,N12086,N12087);
and and7108(N12095,N12100,R7);
and and7116(N12108,N12113,R7);
and and7124(N12121,N12126,R7);
and and7132(N12134,R6,N12139);
and and7140(N12147,N12152,R7);
and and7148(N12160,R6,N12165);
and and7156(N12173,N12177,N12178);
and and7164(N12186,N12191,R7);
and and7172(N12199,N12203,N12204);
and and7180(N12212,N12217,R7);
and and7188(N12225,R6,R7);
and and7196(N12238,N12242,N12243);
and and7204(N12251,R6,N12256);
and and7212(N12264,R6,N12269);
and and7220(N12277,R6,N12282);
and and7228(N12290,N12294,N12295);
and and7236(N12303,N12307,N12308);
and and7244(N12316,R4,N12321);
and and7252(N12329,N12333,N12334);
and and7260(N12342,R6,N12347);
and and7268(N12355,N12359,N12360);
and and7276(N12368,N12372,N12373);
and and7284(N12381,R6,N12386);
and and7292(N12394,R4,N12399);
and and7300(N12407,N12412,R7);
and and7308(N12420,R6,N12425);
and and7316(N12433,N12438,R6);
and and7324(N12446,N12451,R7);
and and7332(N12459,N12464,R7);
and and7340(N12472,N12477,R7);
and and7348(N12485,N12489,N12490);
and and7356(N12498,R5,N12503);
and and7364(N12511,N12516,R7);
and and7372(N12524,N12529,R7);
and and7380(N12537,N12541,N12542);
and and7388(N12550,R5,N12555);
and and7396(N12563,N12567,N12568);
and and7404(N12576,N12580,N12581);
and and7412(N12589,R6,N12594);
and and7420(N12602,R6,N12607);
and and7428(N12615,N12619,N12620);
and and7436(N12628,R6,N12633);
and and7444(N12641,R6,N12646);
and and7452(N12654,R5,N12659);
and and7460(N12667,R6,N12672);
and and7468(N12680,N12683,N12684);
and and7476(N12692,N12695,N12696);
and and7484(N12704,R6,N12708);
and and7492(N12716,N12720,R5);
and and7500(N12728,R6,N12732);
and and7508(N12740,N12744,R7);
and and7516(N12752,N12755,N12756);
and and7524(N12764,N12767,N12768);
and and7532(N12776,N12780,R7);
and and7540(N12788,N12792,R7);
and and7548(N12800,N12804,R7);
and and7556(N12812,R6,R7);
and and7564(N12824,R6,R7);
and and7572(N12836,R6,R7);
and and7580(N12848,R6,N12852);
and and7588(N12860,R6,N12864);
and and7596(N12872,N12875,N12876);
and and7604(N12884,N12887,N12888);
and and7612(N12896,N12900,R7);
and and7620(N12908,R6,R7);
and and7628(N12920,N12923,N12924);
and and7636(N12932,N12935,N12936);
and and7644(N12944,R6,N12948);
and and7652(N12956,R4,N12960);
and and7660(N12968,N12971,N12972);
and and7668(N12980,R5,N12984);
and and7676(N12992,N12995,N12996);
and and7684(N13004,R6,R7);
and and7692(N13016,R6,R7);
and and7700(N13028,R5,N13032);
and and7708(N13040,R6,N13044);
and and7716(N13052,R5,R6);
and and7724(N13064,R5,R6);
and and7732(N13076,N13080,R7);
and and7740(N13088,R5,N13092);
and and7748(N13100,R5,N13104);
and and7756(N13112,N13115,N13116);
and and7764(N13124,R6,N13128);
and and7772(N13136,R6,N13140);
and and7780(N13148,N13152,R7);
and and7788(N13160,N13164,R7);
and and7796(N13172,N13176,R7);
and and7804(N13184,R6,N13188);
and and7812(N13196,N13200,R7);
and and7820(N13208,R4,R7);
and and7828(N13220,N13224,R7);
and and7836(N13232,R6,N13236);
and and7844(N13244,N13247,N13248);
and and7852(N13256,R6,R7);
and and7860(N13268,R5,R6);
and and7868(N13280,R5,N13284);
and and7876(N13292,N13295,N13296);
and and7884(N13304,R6,N13308);
and and7892(N13316,N13319,N13320);
and and7900(N13328,R5,N13332);
and and7908(N13340,N13344,R7);
and and7916(N13352,R6,N13356);
and and7924(N13364,R5,R6);
and and7932(N13376,N13380,R7);
and and7940(N13388,N13392,R7);
and and7948(N13400,N13402,N13403);
and and7956(N13411,N13413,N13414);
and and7964(N13422,R5,N13425);
and and7972(N13433,R5,R7);
and and7980(N13444,N13446,N13447);
and and7988(N13455,R5,R7);
and and7996(N13466,R6,R7);
and and8004(N13477,N13480,R7);
and and8012(N13488,R6,N13491);
and and8020(N13499,R6,N13502);
and and8028(N13510,R6,N13513);
and and8036(N13521,R6,R7);
and and8044(N13532,R6,R7);
and and8052(N13543,R6,R7);
and and8060(N13554,N13557,R7);
and and8068(N13565,N13568,R7);
and and8076(N13576,R6,R7);
and and8084(N13587,R6,R7);
and and8092(N13598,R6,N13601);
and and8100(N13609,R5,R6);
and and8108(N13620,R6,N13623);
and and8116(N13631,R6,R7);
and and8124(N13642,N13644,N13645);
and and8132(N13653,R6,N13656);
and and8140(N13664,R6,N13667);
and and8148(N13675,N13677,N13678);
and and8156(N13686,N13688,N13689);
and and8164(N13697,R4,N13700);
and and8172(N13708,R6,R7);
and and8180(N13719,R6,R7);
and and8188(N13730,R6,R7);
and and8196(N13741,N13744,R7);
and and8204(N13752,R6,N13755);
and and8212(N13763,R6,R7);
and and8220(N13774,N13777,R7);
and and8228(N13785,N13788,R7);
and and8236(N13796,N13799,R7);
and and8244(N13807,N13810,R7);
and and8252(N13818,N13821,R7);
and and8260(N13829,N13832,R7);
and and8268(N13840,N13843,R7);
and and8276(N13851,R5,N13854);
and and8284(N13862,N13865,R7);
and and8292(N13873,R5,R6);
and and8300(N13884,N13887,R7);
and and8308(N13895,N13897,N13898);
and and8316(N13906,R5,R6);
and and8324(N13917,N13920,R7);
and and8332(N13928,N13931,R7);
and and8340(N13939,R5,R6);
and and8348(N13950,N13952,N13953);
and and8356(N13961,R6,N13963);
and and8364(N13971,N13972,N13973);
and and8372(N13981,R5,R7);
and and8380(N13991,R6,R7);
and and8388(N14001,R6,R7);
and and8396(N14011,R6,R7);
and and8404(N14021,R6,R7);
and and8412(N14031,R6,R7);
and and8420(N14041,N14042,N14043);
and and8428(N14051,R6,R7);
and and8436(N14061,N14063,R7);
and and8444(N14071,R6,R7);
and and8452(N14081,R6,R7);
and and8460(N14091,R5,N14093);
and and8468(N14101,N14103,R7);
and and8476(N14111,N14112,N14113);
and and8484(N14121,R6,R7);
and and8492(N14130,R6,R7);
and and8500(N14139,R6,R7);
and and8508(N14148,R6,N14149);
and and8516(N14157,R5,R6);
and and8524(N14166,R6,N14167);
and and8532(N14175,R6,N14176);
and and8540(N14184,R5,R7);
and and8548(N14193,N14194,R7);
and and8556(N14202,R5,R7);
and and8877(N15146,N15147,N15148);
and and8886(N15164,N15165,N15166);
and and8895(N15181,N15182,N15183);
and and8904(N15198,N15199,N15200);
and and8913(N15214,N15215,N15216);
and and8922(N15230,N15231,N15232);
and and8931(N15246,N15247,N15248);
and and8940(N15262,N15263,N15264);
and and8949(N15278,N15279,N15280);
and and8958(N15294,N15295,N15296);
and and8967(N15310,N15311,N15312);
and and8976(N15326,N15327,N15328);
and and8985(N15342,N15343,N15344);
and and8994(N15357,N15358,N15359);
and and9003(N15372,N15373,N15374);
and and9012(N15387,N15388,N15389);
and and9021(N15402,N15403,N15404);
and and9030(N15417,N15418,N15419);
and and9039(N15432,N15433,N15434);
and and9048(N15447,N15448,N15449);
and and9057(N15462,N15463,N15464);
and and9066(N15477,N15478,N15479);
and and9075(N15492,N15493,N15494);
and and9084(N15507,N15508,N15509);
and and9093(N15522,N15523,N15524);
and and9102(N15537,N15538,N15539);
and and9111(N15552,N15553,N15554);
and and9120(N15566,N15567,N15568);
and and9129(N15580,N15581,N15582);
and and9138(N15594,N15595,N15596);
and and9147(N15608,N15609,N15610);
and and9156(N15622,N15623,N15624);
and and9165(N15636,N15637,N15638);
and and9174(N15650,N15651,N15652);
and and9183(N15664,N15665,N15666);
and and9192(N15678,N15679,N15680);
and and9201(N15692,N15693,N15694);
and and9210(N15706,N15707,N15708);
and and9219(N15720,N15721,N15722);
and and9228(N15734,N15735,N15736);
and and9237(N15748,N15749,N15750);
and and9246(N15762,N15763,N15764);
and and9255(N15776,N15777,N15778);
and and9264(N15790,N15791,N15792);
and and9273(N15804,N15805,N15806);
and and9282(N15818,N15819,N15820);
and and9291(N15832,N15833,N15834);
and and9300(N15846,N15847,N15848);
and and9309(N15860,N15861,N15862);
and and9318(N15874,N15875,N15876);
and and9327(N15888,N15889,N15890);
and and9336(N15902,N15903,N15904);
and and9345(N15916,N15917,N15918);
and and9354(N15930,N15931,N15932);
and and9363(N15944,N15945,N15946);
and and9372(N15958,N15959,N15960);
and and9381(N15972,N15973,N15974);
and and9390(N15986,N15987,N15988);
and and9399(N16000,N16001,N16002);
and and9408(N16014,N16015,N16016);
and and9417(N16028,N16029,N16030);
and and9426(N16042,N16043,N16044);
and and9435(N16056,N16057,N16058);
and and9444(N16070,N16071,N16072);
and and9453(N16084,N16085,N16086);
and and9462(N16098,N16099,N16100);
and and9471(N16111,N16112,N16113);
and and9480(N16124,N16125,N16126);
and and9489(N16137,N16138,N16139);
and and9498(N16150,N16151,N16152);
and and9507(N16163,N16164,N16165);
and and9516(N16176,N16177,N16178);
and and9525(N16189,N16190,N16191);
and and9534(N16202,N16203,N16204);
and and9543(N16215,N16216,N16217);
and and9552(N16228,N16229,N16230);
and and9561(N16241,N16242,N16243);
and and9570(N16254,N16255,N16256);
and and9579(N16267,N16268,N16269);
and and9588(N16280,N16281,N16282);
and and9597(N16293,N16294,N16295);
and and9606(N16306,N16307,N16308);
and and9615(N16319,N16320,N16321);
and and9624(N16332,N16333,N16334);
and and9633(N16345,N16346,N16347);
and and9642(N16358,N16359,N16360);
and and9651(N16371,N16372,N16373);
and and9660(N16384,N16385,N16386);
and and9669(N16397,N16398,N16399);
and and9678(N16410,N16411,N16412);
and and9687(N16422,N16423,N16424);
and and9696(N16434,N16435,N16436);
and and9705(N16446,N16447,N16448);
and and9714(N16458,N16459,N16460);
and and9723(N16470,N16471,N16472);
and and9732(N16482,N16483,N16484);
and and9741(N16494,N16495,N16496);
and and9750(N16506,N16507,N16508);
and and9759(N16518,N16519,N16520);
and and9768(N16530,N16531,N16532);
and and9777(N16542,N16543,N16544);
and and9786(N16554,N16555,N16556);
and and9795(N16566,N16567,N16568);
and and9804(N16578,N16579,N16580);
and and9813(N16590,N16591,N16592);
and and9822(N16602,N16603,N16604);
and and9831(N16614,N16615,N16616);
and and9840(N16626,N16627,N16628);
and and9849(N16638,N16639,N16640);
and and9858(N16650,N16651,N16652);
and and9867(N16662,N16663,N16664);
and and9876(N16674,N16675,N16676);
and and9885(N16686,N16687,N16688);
and and9894(N16698,N16699,N16700);
and and9903(N16710,N16711,N16712);
and and9912(N16722,N16723,N16724);
and and9921(N16734,N16735,N16736);
and and9930(N16746,N16747,N16748);
and and9939(N16758,N16759,N16760);
and and9948(N16770,N16771,N16772);
and and9957(N16782,N16783,N16784);
and and9966(N16794,N16795,N16796);
and and9975(N16806,N16807,N16808);
and and9984(N16818,N16819,N16820);
and and9993(N16830,N16831,N16832);
and and10002(N16842,N16843,N16844);
and and10011(N16854,N16855,N16856);
and and10020(N16866,N16867,N16868);
and and10029(N16878,N16879,N16880);
and and10038(N16890,N16891,N16892);
and and10047(N16901,N16902,N16903);
and and10056(N16912,N16913,N16914);
and and10065(N16923,N16924,N16925);
and and10074(N16934,N16935,N16936);
and and10083(N16945,N16946,N16947);
and and10092(N16955,N16956,N16957);
and and10101(N16965,N16966,N16967);
and and10110(N16975,N16976,N16977);
and and10119(N16985,N16986,N16987);
and and10128(N16995,N16996,N16997);
and and10137(N17005,N17006,N17007);
and and10146(N17015,N17016,N17017);
and and10155(N17025,N17026,N17027);
and and10163(N17041,N17042,N17043);
and and10171(N17057,N17058,N17059);
and and10179(N17072,N17073,N17074);
and and10187(N17087,N17088,N17089);
and and10195(N17102,N17103,N17104);
and and10203(N17117,N17118,N17119);
and and10211(N17132,N17133,N17134);
and and10219(N17147,N17148,N17149);
and and10227(N17162,N17163,N17164);
and and10235(N17177,N17178,N17179);
and and10243(N17192,N17193,N17194);
and and10251(N17207,N17208,N17209);
and and10259(N17222,N17223,N17224);
and and10267(N17237,N17238,N17239);
and and10275(N17252,N17253,N17254);
and and10283(N17267,N17268,N17269);
and and10291(N17282,N17283,N17284);
and and10299(N17297,N17298,N17299);
and and10307(N17311,N17312,N17313);
and and10315(N17325,N17326,N17327);
and and10323(N17339,N17340,N17341);
and and10331(N17353,N17354,N17355);
and and10339(N17367,N17368,N17369);
and and10347(N17381,N17382,N17383);
and and10355(N17395,N17396,N17397);
and and10363(N17409,N17410,N17411);
and and10371(N17423,N17424,N17425);
and and10379(N17437,N17438,N17439);
and and10387(N17451,N17452,N17453);
and and10395(N17465,N17466,N17467);
and and10403(N17479,N17480,N17481);
and and10411(N17493,N17494,N17495);
and and10419(N17507,N17508,N17509);
and and10427(N17521,N17522,N17523);
and and10435(N17535,N17536,N17537);
and and10443(N17549,N17550,N17551);
and and10451(N17563,N17564,N17565);
and and10459(N17577,N17578,N17579);
and and10467(N17591,N17592,N17593);
and and10475(N17605,N17606,N17607);
and and10483(N17619,N17620,N17621);
and and10491(N17633,N17634,N17635);
and and10499(N17647,N17648,N17649);
and and10507(N17661,N17662,N17663);
and and10515(N17675,N17676,N17677);
and and10523(N17689,N17690,N17691);
and and10531(N17703,N17704,N17705);
and and10539(N17717,N17718,N17719);
and and10547(N17731,N17732,N17733);
and and10555(N17745,N17746,N17747);
and and10563(N17759,N17760,N17761);
and and10571(N17772,N17773,N17774);
and and10579(N17785,N17786,N17787);
and and10587(N17798,N17799,N17800);
and and10595(N17811,N17812,N17813);
and and10603(N17824,N17825,N17826);
and and10611(N17837,N17838,N17839);
and and10619(N17850,N17851,N17852);
and and10627(N17863,N17864,N17865);
and and10635(N17876,N17877,N17878);
and and10643(N17889,N17890,N17891);
and and10651(N17902,N17903,N17904);
and and10659(N17915,N17916,N17917);
and and10667(N17928,N17929,N17930);
and and10675(N17941,N17942,N17943);
and and10683(N17954,N17955,N17956);
and and10691(N17967,N17968,N17969);
and and10699(N17980,N17981,N17982);
and and10707(N17993,N17994,N17995);
and and10715(N18006,N18007,N18008);
and and10723(N18019,N18020,N18021);
and and10731(N18032,N18033,N18034);
and and10739(N18045,N18046,N18047);
and and10747(N18058,N18059,N18060);
and and10755(N18071,N18072,N18073);
and and10763(N18084,N18085,N18086);
and and10771(N18097,N18098,N18099);
and and10779(N18110,N18111,N18112);
and and10787(N18123,N18124,N18125);
and and10795(N18136,N18137,N18138);
and and10803(N18149,N18150,N18151);
and and10811(N18162,N18163,N18164);
and and10819(N18175,N18176,N18177);
and and10827(N18188,N18189,N18190);
and and10835(N18201,N18202,N18203);
and and10843(N18214,N18215,N18216);
and and10851(N18227,N18228,N18229);
and and10859(N18240,N18241,N18242);
and and10867(N18253,N18254,N18255);
and and10875(N18266,N18267,N18268);
and and10883(N18279,N18280,N18281);
and and10891(N18292,N18293,N18294);
and and10899(N18305,N18306,N18307);
and and10907(N18318,N18319,N18320);
and and10915(N18331,N18332,N18333);
and and10923(N18344,N18345,N18346);
and and10931(N18357,N18358,N18359);
and and10939(N18370,N18371,N18372);
and and10947(N18383,N18384,N18385);
and and10955(N18396,N18397,N18398);
and and10963(N18409,N18410,N18411);
and and10971(N18422,N18423,N18424);
and and10979(N18435,N18436,N18437);
and and10987(N18448,N18449,N18450);
and and10995(N18461,N18462,N18463);
and and11003(N18474,N18475,N18476);
and and11011(N18487,N18488,N18489);
and and11019(N18500,N18501,N18502);
and and11027(N18513,N18514,N18515);
and and11035(N18526,N18527,N18528);
and and11043(N18539,N18540,N18541);
and and11051(N18552,N18553,N18554);
and and11059(N18565,N18566,N18567);
and and11067(N18578,N18579,N18580);
and and11075(N18591,N18592,N18593);
and and11083(N18603,N18604,N18605);
and and11091(N18615,N18616,N18617);
and and11099(N18627,N18628,N18629);
and and11107(N18639,N18640,N18641);
and and11115(N18651,N18652,N18653);
and and11123(N18663,N18664,N18665);
and and11131(N18675,N18676,N18677);
and and11139(N18687,N18688,N18689);
and and11147(N18699,N18700,N18701);
and and11155(N18711,N18712,N18713);
and and11163(N18723,N18724,N18725);
and and11171(N18735,N18736,N18737);
and and11179(N18747,N18748,N18749);
and and11187(N18759,N18760,N18761);
and and11195(N18771,N18772,N18773);
and and11203(N18783,N18784,N18785);
and and11211(N18795,N18796,N18797);
and and11219(N18807,N18808,N18809);
and and11227(N18819,N18820,N18821);
and and11235(N18831,N18832,N18833);
and and11243(N18843,N18844,N18845);
and and11251(N18855,N18856,N18857);
and and11259(N18867,N18868,N18869);
and and11267(N18879,N18880,N18881);
and and11275(N18891,N18892,N18893);
and and11283(N18903,N18904,N18905);
and and11291(N18915,N18916,N18917);
and and11299(N18927,N18928,N18929);
and and11307(N18939,N18940,N18941);
and and11315(N18951,N18952,N18953);
and and11323(N18963,N18964,N18965);
and and11331(N18975,N18976,N18977);
and and11339(N18987,N18988,N18989);
and and11347(N18999,N19000,N19001);
and and11355(N19011,N19012,N19013);
and and11363(N19023,N19024,N19025);
and and11371(N19035,N19036,N19037);
and and11379(N19047,N19048,N19049);
and and11387(N19059,N19060,N19061);
and and11395(N19071,N19072,N19073);
and and11403(N19083,N19084,N19085);
and and11411(N19095,N19096,N19097);
and and11419(N19107,N19108,N19109);
and and11427(N19119,N19120,N19121);
and and11435(N19131,N19132,N19133);
and and11443(N19143,N19144,N19145);
and and11451(N19155,N19156,N19157);
and and11459(N19166,N19167,N19168);
and and11467(N19177,N19178,N19179);
and and11475(N19188,N19189,N19190);
and and11483(N19199,N19200,N19201);
and and11491(N19210,N19211,N19212);
and and11499(N19221,N19222,N19223);
and and11507(N19232,N19233,N19234);
and and11515(N19243,N19244,N19245);
and and11523(N19254,N19255,N19256);
and and11531(N19265,N19266,N19267);
and and11539(N19276,N19277,N19278);
and and11547(N19287,N19288,N19289);
and and11555(N19298,N19299,N19300);
and and11563(N19309,N19310,N19311);
and and11571(N19320,N19321,N19322);
and and11579(N19331,N19332,N19333);
and and11587(N19342,N19343,N19344);
and and11595(N19353,N19354,N19355);
and and11603(N19364,N19365,N19366);
and and11611(N19375,N19376,N19377);
and and11619(N19386,N19387,N19388);
and and11627(N19397,N19398,N19399);
and and11635(N19408,N19409,N19410);
and and11643(N19419,N19420,N19421);
and and11651(N19430,N19431,N19432);
and and11659(N19441,N19442,N19443);
and and11667(N19452,N19453,N19454);
and and11675(N19463,N19464,N19465);
and and11683(N19474,N19475,N19476);
and and11691(N19485,N19486,N19487);
and and11699(N19496,N19497,N19498);
and and11707(N19507,N19508,N19509);
and and11715(N19518,N19519,N19520);
and and11723(N19529,N19530,N19531);
and and11731(N19540,N19541,N19542);
and and11739(N19551,N19552,N19553);
and and11747(N19562,N19563,N19564);
and and11755(N19573,N19574,N19575);
and and11763(N19583,N19584,N19585);
and and11771(N19593,N19594,N19595);
and and11779(N19603,N19604,N19605);
and and11787(N19613,N19614,N19615);
and and11795(N19623,N19624,N19625);
and and11803(N19633,N19634,N19635);
and and11811(N19643,N19644,N19645);
and and11819(N19653,N19654,N19655);
and and11827(N19663,N19664,N19665);
and and11835(N19673,N19674,N19675);
and and11843(N19683,N19684,N19685);
and and11851(N19693,N19694,N19695);
and and11859(N19703,N19704,N19705);
and and11867(N19713,N19714,N19715);
and and11875(N19723,N19724,N19725);
and and11883(N19733,N19734,N19735);
and and11891(N19743,N19744,N19745);
and and11899(N19753,N19754,N19755);
and and11907(N19763,N19764,N19765);
and and11915(N19772,N19773,N19774);
and and11923(N19781,N19782,N19783);
and and11931(N19790,N19791,N19792);
and and11939(N19799,N19800,N19801);
and and11947(N19808,N19809,N19810);
and and11955(N19817,N19818,N19819);
and and11963(N19826,N19827,N19828);
and and11971(N19835,N19836,N19837);
and and11979(N19844,N19845,N19846);
and and11987(N19852,N19853,N19854);
and and11994(N19866,N19867,N19868);
and and12001(N19880,N19881,N19882);
and and12008(N19894,N19895,N19896);
and and12015(N19908,N19909,N19910);
and and12022(N19922,N19923,N19924);
and and12029(N19935,N19936,N19937);
and and12036(N19948,N19949,N19950);
and and12043(N19961,N19962,N19963);
and and12050(N19973,N19974,N19975);
and and12057(N19985,N19986,N19987);
and and12064(N19997,N19998,N19999);
and and12071(N20009,N20010,N20011);
and and12078(N20021,N20022,N20023);
and and12085(N20033,N20034,N20035);
and and12092(N20045,N20046,N20047);
and and12099(N20057,N20058,N20059);
and and12106(N20069,N20070,N20071);
and and12113(N20081,N20082,N20083);
and and12120(N20092,N20093,N20094);
and and12127(N20103,N20104,N20105);
and and12134(N20114,N20115,N20116);
and and12141(N20125,N20126,N20127);
and and12148(N20136,N20137,N20138);
and and12155(N20147,N20148,N20149);
and and12162(N20158,N20159,N20160);
and and12169(N20169,N20170,N20171);
and and12176(N20180,N20181,N20182);
and and12183(N20191,N20192,N20193);
and and12190(N20202,N20203,N20204);
and and12197(N20213,N20214,N20215);
and and12204(N20224,N20225,N20226);
and and12211(N20234,N20235,N20236);
and and12218(N20244,N20245,N20246);
and and12225(N20254,N20255,N20256);
and and12232(N20264,N20265,N20266);
and and12239(N20274,N20275,N20276);
and and12246(N20284,N20285,N20286);
and and12253(N20294,N20295,N20296);
and and12260(N20304,N20305,N20306);
and and12267(N20314,N20315,N20316);
and and12274(N20324,N20325,N20326);
and and12281(N20334,N20335,N20336);
and and12288(N20343,N20344,N20345);
and and12295(N20352,N20353,N20354);
and and12302(N20361,N20362,N20363);
and and12309(N20370,N20371,N20372);
and and12316(N20378,N20379,N20380);
and and12323(N20386,N20387,N20388);
and and12330(N20394,N20395,N20396);
and and8878(N15147,N15149,N15150);
and and8879(N15148,N15151,N15152);
and and8887(N15165,N15167,N15168);
and and8888(N15166,N15169,N15170);
and and8896(N15182,N15184,N15185);
and and8897(N15183,N15186,N15187);
and and8905(N15199,N15201,N15202);
and and8906(N15200,N15203,N15204);
and and8914(N15215,N15217,N15218);
and and8915(N15216,N15219,N15220);
and and8923(N15231,N15233,N15234);
and and8924(N15232,N15235,N15236);
and and8932(N15247,N15249,N15250);
and and8933(N15248,N15251,N15252);
and and8941(N15263,N15265,N15266);
and and8942(N15264,N15267,N15268);
and and8950(N15279,N15281,N15282);
and and8951(N15280,N15283,N15284);
and and8959(N15295,N15297,N15298);
and and8960(N15296,N15299,N15300);
and and8968(N15311,N15313,N15314);
and and8969(N15312,N15315,N15316);
and and8977(N15327,N15329,N15330);
and and8978(N15328,N15331,N15332);
and and8986(N15343,N15345,N15346);
and and8987(N15344,N15347,N15348);
and and8995(N15358,N15360,N15361);
and and8996(N15359,N15362,N15363);
and and9004(N15373,N15375,N15376);
and and9005(N15374,N15377,N15378);
and and9013(N15388,N15390,N15391);
and and9014(N15389,N15392,N15393);
and and9022(N15403,N15405,N15406);
and and9023(N15404,N15407,N15408);
and and9031(N15418,N15420,N15421);
and and9032(N15419,N15422,N15423);
and and9040(N15433,N15435,N15436);
and and9041(N15434,N15437,N15438);
and and9049(N15448,N15450,N15451);
and and9050(N15449,N15452,N15453);
and and9058(N15463,N15465,N15466);
and and9059(N15464,N15467,N15468);
and and9067(N15478,N15480,N15481);
and and9068(N15479,N15482,N15483);
and and9076(N15493,N15495,N15496);
and and9077(N15494,N15497,N15498);
and and9085(N15508,N15510,N15511);
and and9086(N15509,N15512,N15513);
and and9094(N15523,N15525,N15526);
and and9095(N15524,N15527,N15528);
and and9103(N15538,N15540,N15541);
and and9104(N15539,N15542,N15543);
and and9112(N15553,N15555,N15556);
and and9113(N15554,N15557,N15558);
and and9121(N15567,N15569,N15570);
and and9122(N15568,N15571,N15572);
and and9130(N15581,N15583,N15584);
and and9131(N15582,N15585,N15586);
and and9139(N15595,N15597,N15598);
and and9140(N15596,N15599,N15600);
and and9148(N15609,N15611,N15612);
and and9149(N15610,N15613,N15614);
and and9157(N15623,N15625,N15626);
and and9158(N15624,N15627,N15628);
and and9166(N15637,N15639,N15640);
and and9167(N15638,N15641,N15642);
and and9175(N15651,N15653,N15654);
and and9176(N15652,N15655,N15656);
and and9184(N15665,N15667,N15668);
and and9185(N15666,N15669,N15670);
and and9193(N15679,N15681,N15682);
and and9194(N15680,N15683,N15684);
and and9202(N15693,N15695,N15696);
and and9203(N15694,N15697,N15698);
and and9211(N15707,N15709,N15710);
and and9212(N15708,N15711,N15712);
and and9220(N15721,N15723,N15724);
and and9221(N15722,N15725,N15726);
and and9229(N15735,N15737,N15738);
and and9230(N15736,N15739,N15740);
and and9238(N15749,N15751,N15752);
and and9239(N15750,N15753,N15754);
and and9247(N15763,N15765,N15766);
and and9248(N15764,N15767,N15768);
and and9256(N15777,N15779,N15780);
and and9257(N15778,N15781,N15782);
and and9265(N15791,N15793,N15794);
and and9266(N15792,N15795,N15796);
and and9274(N15805,N15807,N15808);
and and9275(N15806,N15809,N15810);
and and9283(N15819,N15821,N15822);
and and9284(N15820,N15823,N15824);
and and9292(N15833,N15835,N15836);
and and9293(N15834,N15837,N15838);
and and9301(N15847,N15849,N15850);
and and9302(N15848,N15851,N15852);
and and9310(N15861,N15863,N15864);
and and9311(N15862,N15865,N15866);
and and9319(N15875,N15877,N15878);
and and9320(N15876,N15879,N15880);
and and9328(N15889,N15891,N15892);
and and9329(N15890,N15893,N15894);
and and9337(N15903,N15905,N15906);
and and9338(N15904,N15907,N15908);
and and9346(N15917,N15919,N15920);
and and9347(N15918,N15921,N15922);
and and9355(N15931,N15933,N15934);
and and9356(N15932,N15935,N15936);
and and9364(N15945,N15947,N15948);
and and9365(N15946,N15949,N15950);
and and9373(N15959,N15961,N15962);
and and9374(N15960,N15963,N15964);
and and9382(N15973,N15975,N15976);
and and9383(N15974,N15977,N15978);
and and9391(N15987,N15989,N15990);
and and9392(N15988,N15991,N15992);
and and9400(N16001,N16003,N16004);
and and9401(N16002,N16005,N16006);
and and9409(N16015,N16017,N16018);
and and9410(N16016,N16019,N16020);
and and9418(N16029,N16031,N16032);
and and9419(N16030,N16033,N16034);
and and9427(N16043,N16045,N16046);
and and9428(N16044,N16047,N16048);
and and9436(N16057,N16059,N16060);
and and9437(N16058,N16061,N16062);
and and9445(N16071,N16073,N16074);
and and9446(N16072,N16075,N16076);
and and9454(N16085,N16087,N16088);
and and9455(N16086,N16089,N16090);
and and9463(N16099,N16101,N16102);
and and9464(N16100,N16103,N16104);
and and9472(N16112,N16114,N16115);
and and9473(N16113,N16116,N16117);
and and9481(N16125,N16127,N16128);
and and9482(N16126,N16129,N16130);
and and9490(N16138,N16140,N16141);
and and9491(N16139,N16142,N16143);
and and9499(N16151,N16153,N16154);
and and9500(N16152,N16155,N16156);
and and9508(N16164,N16166,N16167);
and and9509(N16165,N16168,N16169);
and and9517(N16177,N16179,N16180);
and and9518(N16178,N16181,N16182);
and and9526(N16190,N16192,N16193);
and and9527(N16191,N16194,N16195);
and and9535(N16203,N16205,N16206);
and and9536(N16204,N16207,N16208);
and and9544(N16216,N16218,N16219);
and and9545(N16217,N16220,N16221);
and and9553(N16229,N16231,N16232);
and and9554(N16230,N16233,N16234);
and and9562(N16242,N16244,N16245);
and and9563(N16243,N16246,N16247);
and and9571(N16255,N16257,N16258);
and and9572(N16256,N16259,N16260);
and and9580(N16268,N16270,N16271);
and and9581(N16269,N16272,N16273);
and and9589(N16281,N16283,N16284);
and and9590(N16282,N16285,N16286);
and and9598(N16294,N16296,N16297);
and and9599(N16295,N16298,N16299);
and and9607(N16307,N16309,N16310);
and and9608(N16308,N16311,N16312);
and and9616(N16320,N16322,N16323);
and and9617(N16321,N16324,N16325);
and and9625(N16333,N16335,N16336);
and and9626(N16334,N16337,N16338);
and and9634(N16346,N16348,N16349);
and and9635(N16347,N16350,N16351);
and and9643(N16359,N16361,N16362);
and and9644(N16360,N16363,N16364);
and and9652(N16372,N16374,N16375);
and and9653(N16373,N16376,N16377);
and and9661(N16385,N16387,N16388);
and and9662(N16386,N16389,N16390);
and and9670(N16398,N16400,N16401);
and and9671(N16399,N16402,N16403);
and and9679(N16411,N16413,N16414);
and and9680(N16412,N16415,N16416);
and and9688(N16423,N16425,N16426);
and and9689(N16424,N16427,N16428);
and and9697(N16435,N16437,N16438);
and and9698(N16436,N16439,N16440);
and and9706(N16447,N16449,N16450);
and and9707(N16448,N16451,N16452);
and and9715(N16459,N16461,N16462);
and and9716(N16460,N16463,N16464);
and and9724(N16471,N16473,N16474);
and and9725(N16472,N16475,N16476);
and and9733(N16483,N16485,N16486);
and and9734(N16484,N16487,N16488);
and and9742(N16495,N16497,N16498);
and and9743(N16496,N16499,N16500);
and and9751(N16507,N16509,N16510);
and and9752(N16508,N16511,N16512);
and and9760(N16519,N16521,N16522);
and and9761(N16520,N16523,N16524);
and and9769(N16531,N16533,N16534);
and and9770(N16532,N16535,N16536);
and and9778(N16543,N16545,N16546);
and and9779(N16544,N16547,N16548);
and and9787(N16555,N16557,N16558);
and and9788(N16556,N16559,N16560);
and and9796(N16567,N16569,N16570);
and and9797(N16568,N16571,N16572);
and and9805(N16579,N16581,N16582);
and and9806(N16580,N16583,N16584);
and and9814(N16591,N16593,N16594);
and and9815(N16592,N16595,N16596);
and and9823(N16603,N16605,N16606);
and and9824(N16604,N16607,N16608);
and and9832(N16615,N16617,N16618);
and and9833(N16616,N16619,N16620);
and and9841(N16627,N16629,N16630);
and and9842(N16628,N16631,N16632);
and and9850(N16639,N16641,N16642);
and and9851(N16640,N16643,N16644);
and and9859(N16651,N16653,N16654);
and and9860(N16652,N16655,N16656);
and and9868(N16663,N16665,N16666);
and and9869(N16664,N16667,N16668);
and and9877(N16675,N16677,N16678);
and and9878(N16676,N16679,N16680);
and and9886(N16687,N16689,N16690);
and and9887(N16688,N16691,N16692);
and and9895(N16699,N16701,N16702);
and and9896(N16700,N16703,N16704);
and and9904(N16711,N16713,N16714);
and and9905(N16712,N16715,N16716);
and and9913(N16723,N16725,N16726);
and and9914(N16724,N16727,N16728);
and and9922(N16735,N16737,N16738);
and and9923(N16736,N16739,N16740);
and and9931(N16747,N16749,N16750);
and and9932(N16748,N16751,N16752);
and and9940(N16759,N16761,N16762);
and and9941(N16760,N16763,N16764);
and and9949(N16771,N16773,N16774);
and and9950(N16772,N16775,N16776);
and and9958(N16783,N16785,N16786);
and and9959(N16784,N16787,N16788);
and and9967(N16795,N16797,N16798);
and and9968(N16796,N16799,N16800);
and and9976(N16807,N16809,N16810);
and and9977(N16808,N16811,N16812);
and and9985(N16819,N16821,N16822);
and and9986(N16820,N16823,N16824);
and and9994(N16831,N16833,N16834);
and and9995(N16832,N16835,N16836);
and and10003(N16843,N16845,N16846);
and and10004(N16844,N16847,N16848);
and and10012(N16855,N16857,N16858);
and and10013(N16856,N16859,N16860);
and and10021(N16867,N16869,N16870);
and and10022(N16868,N16871,N16872);
and and10030(N16879,N16881,N16882);
and and10031(N16880,N16883,N16884);
and and10039(N16891,N16893,N16894);
and and10040(N16892,N16895,N16896);
and and10048(N16902,N16904,N16905);
and and10049(N16903,N16906,N16907);
and and10057(N16913,N16915,N16916);
and and10058(N16914,N16917,N16918);
and and10066(N16924,N16926,N16927);
and and10067(N16925,N16928,N16929);
and and10075(N16935,N16937,N16938);
and and10076(N16936,N16939,N16940);
and and10084(N16946,N16948,N16949);
and and10085(N16947,N16950,N16951);
and and10093(N16956,N16958,N16959);
and and10094(N16957,N16960,N16961);
and and10102(N16966,N16968,N16969);
and and10103(N16967,N16970,N16971);
and and10111(N16976,N16978,N16979);
and and10112(N16977,N16980,N16981);
and and10120(N16986,N16988,N16989);
and and10121(N16987,N16990,N16991);
and and10129(N16996,N16998,N16999);
and and10130(N16997,N17000,N17001);
and and10138(N17006,N17008,N17009);
and and10139(N17007,N17010,N17011);
and and10147(N17016,N17018,N17019);
and and10148(N17017,N17020,N17021);
and and10156(N17026,N17028,N17029);
and and10157(N17027,N17030,N17031);
and and10164(N17042,N17044,N17045);
and and10165(N17043,N17046,N17047);
and and10172(N17058,N17060,N17061);
and and10173(N17059,N17062,N17063);
and and10180(N17073,N17075,N17076);
and and10181(N17074,N17077,N17078);
and and10188(N17088,N17090,N17091);
and and10189(N17089,N17092,N17093);
and and10196(N17103,N17105,N17106);
and and10197(N17104,N17107,N17108);
and and10204(N17118,N17120,N17121);
and and10205(N17119,N17122,N17123);
and and10212(N17133,N17135,N17136);
and and10213(N17134,N17137,N17138);
and and10220(N17148,N17150,N17151);
and and10221(N17149,N17152,N17153);
and and10228(N17163,N17165,N17166);
and and10229(N17164,N17167,N17168);
and and10236(N17178,N17180,N17181);
and and10237(N17179,N17182,N17183);
and and10244(N17193,N17195,N17196);
and and10245(N17194,N17197,N17198);
and and10252(N17208,N17210,N17211);
and and10253(N17209,N17212,N17213);
and and10260(N17223,N17225,N17226);
and and10261(N17224,N17227,N17228);
and and10268(N17238,N17240,N17241);
and and10269(N17239,N17242,N17243);
and and10276(N17253,N17255,N17256);
and and10277(N17254,N17257,N17258);
and and10284(N17268,N17270,N17271);
and and10285(N17269,N17272,N17273);
and and10292(N17283,N17285,N17286);
and and10293(N17284,N17287,N17288);
and and10300(N17298,N17300,N17301);
and and10301(N17299,N17302,N17303);
and and10308(N17312,N17314,N17315);
and and10309(N17313,N17316,N17317);
and and10316(N17326,N17328,N17329);
and and10317(N17327,N17330,N17331);
and and10324(N17340,N17342,N17343);
and and10325(N17341,N17344,N17345);
and and10332(N17354,N17356,N17357);
and and10333(N17355,N17358,N17359);
and and10340(N17368,N17370,N17371);
and and10341(N17369,N17372,N17373);
and and10348(N17382,N17384,N17385);
and and10349(N17383,N17386,N17387);
and and10356(N17396,N17398,N17399);
and and10357(N17397,N17400,N17401);
and and10364(N17410,N17412,N17413);
and and10365(N17411,N17414,N17415);
and and10372(N17424,N17426,N17427);
and and10373(N17425,N17428,N17429);
and and10380(N17438,N17440,N17441);
and and10381(N17439,N17442,N17443);
and and10388(N17452,N17454,N17455);
and and10389(N17453,N17456,N17457);
and and10396(N17466,N17468,N17469);
and and10397(N17467,N17470,N17471);
and and10404(N17480,N17482,N17483);
and and10405(N17481,N17484,N17485);
and and10412(N17494,N17496,N17497);
and and10413(N17495,N17498,N17499);
and and10420(N17508,N17510,N17511);
and and10421(N17509,N17512,N17513);
and and10428(N17522,N17524,N17525);
and and10429(N17523,N17526,N17527);
and and10436(N17536,N17538,N17539);
and and10437(N17537,N17540,N17541);
and and10444(N17550,N17552,N17553);
and and10445(N17551,N17554,N17555);
and and10452(N17564,N17566,N17567);
and and10453(N17565,N17568,N17569);
and and10460(N17578,N17580,N17581);
and and10461(N17579,N17582,N17583);
and and10468(N17592,N17594,N17595);
and and10469(N17593,N17596,N17597);
and and10476(N17606,N17608,N17609);
and and10477(N17607,N17610,N17611);
and and10484(N17620,N17622,N17623);
and and10485(N17621,N17624,N17625);
and and10492(N17634,N17636,N17637);
and and10493(N17635,N17638,N17639);
and and10500(N17648,N17650,N17651);
and and10501(N17649,N17652,N17653);
and and10508(N17662,N17664,N17665);
and and10509(N17663,N17666,N17667);
and and10516(N17676,N17678,N17679);
and and10517(N17677,N17680,N17681);
and and10524(N17690,N17692,N17693);
and and10525(N17691,N17694,N17695);
and and10532(N17704,N17706,N17707);
and and10533(N17705,N17708,N17709);
and and10540(N17718,N17720,N17721);
and and10541(N17719,N17722,N17723);
and and10548(N17732,N17734,N17735);
and and10549(N17733,N17736,N17737);
and and10556(N17746,N17748,N17749);
and and10557(N17747,N17750,N17751);
and and10564(N17760,N17762,N17763);
and and10565(N17761,N17764,N17765);
and and10572(N17773,N17775,N17776);
and and10573(N17774,N17777,N17778);
and and10580(N17786,N17788,N17789);
and and10581(N17787,N17790,N17791);
and and10588(N17799,N17801,N17802);
and and10589(N17800,N17803,N17804);
and and10596(N17812,N17814,N17815);
and and10597(N17813,N17816,N17817);
and and10604(N17825,N17827,N17828);
and and10605(N17826,N17829,N17830);
and and10612(N17838,N17840,N17841);
and and10613(N17839,N17842,N17843);
and and10620(N17851,N17853,N17854);
and and10621(N17852,N17855,N17856);
and and10628(N17864,N17866,N17867);
and and10629(N17865,N17868,N17869);
and and10636(N17877,N17879,N17880);
and and10637(N17878,N17881,N17882);
and and10644(N17890,N17892,N17893);
and and10645(N17891,N17894,N17895);
and and10652(N17903,N17905,N17906);
and and10653(N17904,N17907,N17908);
and and10660(N17916,N17918,N17919);
and and10661(N17917,N17920,N17921);
and and10668(N17929,N17931,N17932);
and and10669(N17930,N17933,N17934);
and and10676(N17942,N17944,N17945);
and and10677(N17943,N17946,N17947);
and and10684(N17955,N17957,N17958);
and and10685(N17956,N17959,N17960);
and and10692(N17968,N17970,N17971);
and and10693(N17969,N17972,N17973);
and and10700(N17981,N17983,N17984);
and and10701(N17982,N17985,N17986);
and and10708(N17994,N17996,N17997);
and and10709(N17995,N17998,N17999);
and and10716(N18007,N18009,N18010);
and and10717(N18008,N18011,N18012);
and and10724(N18020,N18022,N18023);
and and10725(N18021,N18024,N18025);
and and10732(N18033,N18035,N18036);
and and10733(N18034,N18037,N18038);
and and10740(N18046,N18048,N18049);
and and10741(N18047,N18050,N18051);
and and10748(N18059,N18061,N18062);
and and10749(N18060,N18063,N18064);
and and10756(N18072,N18074,N18075);
and and10757(N18073,N18076,N18077);
and and10764(N18085,N18087,N18088);
and and10765(N18086,N18089,N18090);
and and10772(N18098,N18100,N18101);
and and10773(N18099,N18102,N18103);
and and10780(N18111,N18113,N18114);
and and10781(N18112,N18115,N18116);
and and10788(N18124,N18126,N18127);
and and10789(N18125,N18128,N18129);
and and10796(N18137,N18139,N18140);
and and10797(N18138,N18141,N18142);
and and10804(N18150,N18152,N18153);
and and10805(N18151,N18154,N18155);
and and10812(N18163,N18165,N18166);
and and10813(N18164,N18167,N18168);
and and10820(N18176,N18178,N18179);
and and10821(N18177,N18180,N18181);
and and10828(N18189,N18191,N18192);
and and10829(N18190,N18193,N18194);
and and10836(N18202,N18204,N18205);
and and10837(N18203,N18206,N18207);
and and10844(N18215,N18217,N18218);
and and10845(N18216,N18219,N18220);
and and10852(N18228,N18230,N18231);
and and10853(N18229,N18232,N18233);
and and10860(N18241,N18243,N18244);
and and10861(N18242,N18245,N18246);
and and10868(N18254,N18256,N18257);
and and10869(N18255,N18258,N18259);
and and10876(N18267,N18269,N18270);
and and10877(N18268,N18271,N18272);
and and10884(N18280,N18282,N18283);
and and10885(N18281,N18284,N18285);
and and10892(N18293,N18295,N18296);
and and10893(N18294,N18297,N18298);
and and10900(N18306,N18308,N18309);
and and10901(N18307,N18310,N18311);
and and10908(N18319,N18321,N18322);
and and10909(N18320,N18323,N18324);
and and10916(N18332,N18334,N18335);
and and10917(N18333,N18336,N18337);
and and10924(N18345,N18347,N18348);
and and10925(N18346,N18349,N18350);
and and10932(N18358,N18360,N18361);
and and10933(N18359,N18362,N18363);
and and10940(N18371,N18373,N18374);
and and10941(N18372,N18375,N18376);
and and10948(N18384,N18386,N18387);
and and10949(N18385,N18388,N18389);
and and10956(N18397,N18399,N18400);
and and10957(N18398,N18401,N18402);
and and10964(N18410,N18412,N18413);
and and10965(N18411,N18414,N18415);
and and10972(N18423,N18425,N18426);
and and10973(N18424,N18427,N18428);
and and10980(N18436,N18438,N18439);
and and10981(N18437,N18440,N18441);
and and10988(N18449,N18451,N18452);
and and10989(N18450,N18453,N18454);
and and10996(N18462,N18464,N18465);
and and10997(N18463,N18466,N18467);
and and11004(N18475,N18477,N18478);
and and11005(N18476,N18479,N18480);
and and11012(N18488,N18490,N18491);
and and11013(N18489,N18492,N18493);
and and11020(N18501,N18503,N18504);
and and11021(N18502,N18505,N18506);
and and11028(N18514,N18516,N18517);
and and11029(N18515,N18518,N18519);
and and11036(N18527,N18529,N18530);
and and11037(N18528,N18531,N18532);
and and11044(N18540,N18542,N18543);
and and11045(N18541,N18544,N18545);
and and11052(N18553,N18555,N18556);
and and11053(N18554,N18557,N18558);
and and11060(N18566,N18568,N18569);
and and11061(N18567,N18570,N18571);
and and11068(N18579,N18581,N18582);
and and11069(N18580,N18583,N18584);
and and11076(N18592,N18594,N18595);
and and11077(N18593,N18596,N18597);
and and11084(N18604,N18606,N18607);
and and11085(N18605,N18608,N18609);
and and11092(N18616,N18618,N18619);
and and11093(N18617,N18620,N18621);
and and11100(N18628,N18630,N18631);
and and11101(N18629,N18632,N18633);
and and11108(N18640,N18642,N18643);
and and11109(N18641,N18644,N18645);
and and11116(N18652,N18654,N18655);
and and11117(N18653,N18656,N18657);
and and11124(N18664,N18666,N18667);
and and11125(N18665,N18668,N18669);
and and11132(N18676,N18678,N18679);
and and11133(N18677,N18680,N18681);
and and11140(N18688,N18690,N18691);
and and11141(N18689,N18692,N18693);
and and11148(N18700,N18702,N18703);
and and11149(N18701,N18704,N18705);
and and11156(N18712,N18714,N18715);
and and11157(N18713,N18716,N18717);
and and11164(N18724,N18726,N18727);
and and11165(N18725,N18728,N18729);
and and11172(N18736,N18738,N18739);
and and11173(N18737,N18740,N18741);
and and11180(N18748,N18750,N18751);
and and11181(N18749,N18752,N18753);
and and11188(N18760,N18762,N18763);
and and11189(N18761,N18764,N18765);
and and11196(N18772,N18774,N18775);
and and11197(N18773,N18776,N18777);
and and11204(N18784,N18786,N18787);
and and11205(N18785,N18788,N18789);
and and11212(N18796,N18798,N18799);
and and11213(N18797,N18800,N18801);
and and11220(N18808,N18810,N18811);
and and11221(N18809,N18812,N18813);
and and11228(N18820,N18822,N18823);
and and11229(N18821,N18824,N18825);
and and11236(N18832,N18834,N18835);
and and11237(N18833,N18836,N18837);
and and11244(N18844,N18846,N18847);
and and11245(N18845,N18848,N18849);
and and11252(N18856,N18858,N18859);
and and11253(N18857,N18860,N18861);
and and11260(N18868,N18870,N18871);
and and11261(N18869,N18872,N18873);
and and11268(N18880,N18882,N18883);
and and11269(N18881,N18884,N18885);
and and11276(N18892,N18894,N18895);
and and11277(N18893,N18896,N18897);
and and11284(N18904,N18906,N18907);
and and11285(N18905,N18908,N18909);
and and11292(N18916,N18918,N18919);
and and11293(N18917,N18920,N18921);
and and11300(N18928,N18930,N18931);
and and11301(N18929,N18932,N18933);
and and11308(N18940,N18942,N18943);
and and11309(N18941,N18944,N18945);
and and11316(N18952,N18954,N18955);
and and11317(N18953,N18956,N18957);
and and11324(N18964,N18966,N18967);
and and11325(N18965,N18968,N18969);
and and11332(N18976,N18978,N18979);
and and11333(N18977,N18980,N18981);
and and11340(N18988,N18990,N18991);
and and11341(N18989,N18992,N18993);
and and11348(N19000,N19002,N19003);
and and11349(N19001,N19004,N19005);
and and11356(N19012,N19014,N19015);
and and11357(N19013,N19016,N19017);
and and11364(N19024,N19026,N19027);
and and11365(N19025,N19028,N19029);
and and11372(N19036,N19038,N19039);
and and11373(N19037,N19040,N19041);
and and11380(N19048,N19050,N19051);
and and11381(N19049,N19052,N19053);
and and11388(N19060,N19062,N19063);
and and11389(N19061,N19064,N19065);
and and11396(N19072,N19074,N19075);
and and11397(N19073,N19076,N19077);
and and11404(N19084,N19086,N19087);
and and11405(N19085,N19088,N19089);
and and11412(N19096,N19098,N19099);
and and11413(N19097,N19100,N19101);
and and11420(N19108,N19110,N19111);
and and11421(N19109,N19112,N19113);
and and11428(N19120,N19122,N19123);
and and11429(N19121,N19124,N19125);
and and11436(N19132,N19134,N19135);
and and11437(N19133,N19136,N19137);
and and11444(N19144,N19146,N19147);
and and11445(N19145,N19148,N19149);
and and11452(N19156,N19158,N19159);
and and11453(N19157,N19160,N19161);
and and11460(N19167,N19169,N19170);
and and11461(N19168,N19171,N19172);
and and11468(N19178,N19180,N19181);
and and11469(N19179,N19182,N19183);
and and11476(N19189,N19191,N19192);
and and11477(N19190,N19193,N19194);
and and11484(N19200,N19202,N19203);
and and11485(N19201,N19204,N19205);
and and11492(N19211,N19213,N19214);
and and11493(N19212,N19215,N19216);
and and11500(N19222,N19224,N19225);
and and11501(N19223,N19226,N19227);
and and11508(N19233,N19235,N19236);
and and11509(N19234,N19237,N19238);
and and11516(N19244,N19246,N19247);
and and11517(N19245,N19248,N19249);
and and11524(N19255,N19257,N19258);
and and11525(N19256,N19259,N19260);
and and11532(N19266,N19268,N19269);
and and11533(N19267,N19270,N19271);
and and11540(N19277,N19279,N19280);
and and11541(N19278,N19281,N19282);
and and11548(N19288,N19290,N19291);
and and11549(N19289,N19292,N19293);
and and11556(N19299,N19301,N19302);
and and11557(N19300,N19303,N19304);
and and11564(N19310,N19312,N19313);
and and11565(N19311,N19314,N19315);
and and11572(N19321,N19323,N19324);
and and11573(N19322,N19325,N19326);
and and11580(N19332,N19334,N19335);
and and11581(N19333,N19336,N19337);
and and11588(N19343,N19345,N19346);
and and11589(N19344,N19347,N19348);
and and11596(N19354,N19356,N19357);
and and11597(N19355,N19358,N19359);
and and11604(N19365,N19367,N19368);
and and11605(N19366,N19369,N19370);
and and11612(N19376,N19378,N19379);
and and11613(N19377,N19380,N19381);
and and11620(N19387,N19389,N19390);
and and11621(N19388,N19391,N19392);
and and11628(N19398,N19400,N19401);
and and11629(N19399,N19402,N19403);
and and11636(N19409,N19411,N19412);
and and11637(N19410,N19413,N19414);
and and11644(N19420,N19422,N19423);
and and11645(N19421,N19424,N19425);
and and11652(N19431,N19433,N19434);
and and11653(N19432,N19435,N19436);
and and11660(N19442,N19444,N19445);
and and11661(N19443,N19446,N19447);
and and11668(N19453,N19455,N19456);
and and11669(N19454,N19457,N19458);
and and11676(N19464,N19466,N19467);
and and11677(N19465,N19468,N19469);
and and11684(N19475,N19477,N19478);
and and11685(N19476,N19479,N19480);
and and11692(N19486,N19488,N19489);
and and11693(N19487,N19490,N19491);
and and11700(N19497,N19499,N19500);
and and11701(N19498,N19501,N19502);
and and11708(N19508,N19510,N19511);
and and11709(N19509,N19512,N19513);
and and11716(N19519,N19521,N19522);
and and11717(N19520,N19523,N19524);
and and11724(N19530,N19532,N19533);
and and11725(N19531,N19534,N19535);
and and11732(N19541,N19543,N19544);
and and11733(N19542,N19545,N19546);
and and11740(N19552,N19554,N19555);
and and11741(N19553,N19556,N19557);
and and11748(N19563,N19565,N19566);
and and11749(N19564,N19567,N19568);
and and11756(N19574,N19576,N19577);
and and11757(N19575,N19578,N19579);
and and11764(N19584,N19586,N19587);
and and11765(N19585,N19588,N19589);
and and11772(N19594,N19596,N19597);
and and11773(N19595,N19598,N19599);
and and11780(N19604,N19606,N19607);
and and11781(N19605,N19608,N19609);
and and11788(N19614,N19616,N19617);
and and11789(N19615,N19618,N19619);
and and11796(N19624,N19626,N19627);
and and11797(N19625,N19628,N19629);
and and11804(N19634,N19636,N19637);
and and11805(N19635,N19638,N19639);
and and11812(N19644,N19646,N19647);
and and11813(N19645,N19648,N19649);
and and11820(N19654,N19656,N19657);
and and11821(N19655,N19658,N19659);
and and11828(N19664,N19666,N19667);
and and11829(N19665,N19668,N19669);
and and11836(N19674,N19676,N19677);
and and11837(N19675,N19678,N19679);
and and11844(N19684,N19686,N19687);
and and11845(N19685,N19688,N19689);
and and11852(N19694,N19696,N19697);
and and11853(N19695,N19698,N19699);
and and11860(N19704,N19706,N19707);
and and11861(N19705,N19708,N19709);
and and11868(N19714,N19716,N19717);
and and11869(N19715,N19718,N19719);
and and11876(N19724,N19726,N19727);
and and11877(N19725,N19728,N19729);
and and11884(N19734,N19736,N19737);
and and11885(N19735,N19738,N19739);
and and11892(N19744,N19746,N19747);
and and11893(N19745,N19748,N19749);
and and11900(N19754,N19756,N19757);
and and11901(N19755,N19758,N19759);
and and11908(N19764,N19766,N19767);
and and11909(N19765,N19768,N19769);
and and11916(N19773,N19775,N19776);
and and11917(N19774,N19777,N19778);
and and11924(N19782,N19784,N19785);
and and11925(N19783,N19786,N19787);
and and11932(N19791,N19793,N19794);
and and11933(N19792,N19795,N19796);
and and11940(N19800,N19802,N19803);
and and11941(N19801,N19804,N19805);
and and11948(N19809,N19811,N19812);
and and11949(N19810,N19813,N19814);
and and11956(N19818,N19820,N19821);
and and11957(N19819,N19822,N19823);
and and11964(N19827,N19829,N19830);
and and11965(N19828,N19831,N19832);
and and11972(N19836,N19838,N19839);
and and11973(N19837,N19840,N19841);
and and11980(N19845,N19847,N19848);
and and11981(N19846,N19849,N19850);
and and11988(N19853,N19855,N19856);
and and11989(N19854,N19857,N19858);
and and11995(N19867,N19869,N19870);
and and11996(N19868,N19871,N19872);
and and12002(N19881,N19883,N19884);
and and12003(N19882,N19885,N19886);
and and12009(N19895,N19897,N19898);
and and12010(N19896,N19899,N19900);
and and12016(N19909,N19911,N19912);
and and12017(N19910,N19913,N19914);
and and12023(N19923,N19925,N19926);
and and12024(N19924,N19927,N19928);
and and12030(N19936,N19938,N19939);
and and12031(N19937,N19940,N19941);
and and12037(N19949,N19951,N19952);
and and12038(N19950,N19953,N19954);
and and12044(N19962,N19964,N19965);
and and12045(N19963,N19966,N19967);
and and12051(N19974,N19976,N19977);
and and12052(N19975,N19978,N19979);
and and12058(N19986,N19988,N19989);
and and12059(N19987,N19990,N19991);
and and12065(N19998,N20000,N20001);
and and12066(N19999,N20002,N20003);
and and12072(N20010,N20012,N20013);
and and12073(N20011,N20014,N20015);
and and12079(N20022,N20024,N20025);
and and12080(N20023,N20026,N20027);
and and12086(N20034,N20036,N20037);
and and12087(N20035,N20038,N20039);
and and12093(N20046,N20048,N20049);
and and12094(N20047,N20050,N20051);
and and12100(N20058,N20060,N20061);
and and12101(N20059,N20062,N20063);
and and12107(N20070,N20072,N20073);
and and12108(N20071,N20074,N20075);
and and12114(N20082,N20084,N20085);
and and12115(N20083,N20086,N20087);
and and12121(N20093,N20095,N20096);
and and12122(N20094,N20097,N20098);
and and12128(N20104,N20106,N20107);
and and12129(N20105,N20108,N20109);
and and12135(N20115,N20117,N20118);
and and12136(N20116,N20119,N20120);
and and12142(N20126,N20128,N20129);
and and12143(N20127,N20130,N20131);
and and12149(N20137,N20139,N20140);
and and12150(N20138,N20141,N20142);
and and12156(N20148,N20150,N20151);
and and12157(N20149,N20152,N20153);
and and12163(N20159,N20161,N20162);
and and12164(N20160,N20163,N20164);
and and12170(N20170,N20172,N20173);
and and12171(N20171,N20174,N20175);
and and12177(N20181,N20183,N20184);
and and12178(N20182,N20185,N20186);
and and12184(N20192,N20194,N20195);
and and12185(N20193,N20196,N20197);
and and12191(N20203,N20205,N20206);
and and12192(N20204,N20207,N20208);
and and12198(N20214,N20216,N20217);
and and12199(N20215,N20218,N20219);
and and12205(N20225,N20227,N20228);
and and12206(N20226,N20229,N20230);
and and12212(N20235,N20237,N20238);
and and12213(N20236,N20239,N20240);
and and12219(N20245,N20247,N20248);
and and12220(N20246,N20249,N20250);
and and12226(N20255,N20257,N20258);
and and12227(N20256,N20259,N20260);
and and12233(N20265,N20267,N20268);
and and12234(N20266,N20269,N20270);
and and12240(N20275,N20277,N20278);
and and12241(N20276,N20279,N20280);
and and12247(N20285,N20287,N20288);
and and12248(N20286,N20289,N20290);
and and12254(N20295,N20297,N20298);
and and12255(N20296,N20299,N20300);
and and12261(N20305,N20307,N20308);
and and12262(N20306,N20309,N20310);
and and12268(N20315,N20317,N20318);
and and12269(N20316,N20319,N20320);
and and12275(N20325,N20327,N20328);
and and12276(N20326,N20329,N20330);
and and12282(N20335,N20337,N20338);
and and12283(N20336,N20339,N20340);
and and12289(N20344,N20346,N20347);
and and12290(N20345,N20348,N20349);
and and12296(N20353,N20355,N20356);
and and12297(N20354,N20357,N20358);
and and12303(N20362,N20364,N20365);
and and12304(N20363,N20366,N20367);
and and12310(N20371,N20373,N20374);
and and12311(N20372,N20375,N20376);
and and12317(N20379,N20381,N20382);
and and12318(N20380,N20383,N20384);
and and12324(N20387,N20389,N20390);
and and12325(N20388,N20391,N20392);
and and12331(N20395,N20397,N20398);
and and12332(N20396,N20399,in0);
and and8880(N15149,N15153,N15154);
and and8881(N15150,N15155,in1);
and and8882(N15151,N15156,N15157);
and and8883(N15152,N15158,N15159);
and and8889(N15167,N15171,N15172);
and and8890(N15168,in1,N15173);
and and8891(N15169,N15174,N15175);
and and8892(N15170,N15176,N15177);
and and8898(N15184,N15188,N15189);
and and8899(N15185,in1,N15190);
and and8900(N15186,N15191,N15192);
and and8901(N15187,N15193,N15194);
and and8907(N15201,N15205,N15206);
and and8908(N15202,N15207,N15208);
and and8909(N15203,R0,N15209);
and and8910(N15204,R2,R3);
and and8916(N15217,N15221,N15222);
and and8917(N15218,in0,in1);
and and8918(N15219,N15223,N15224);
and and8919(N15220,N15225,R3);
and and8925(N15233,N15237,N15238);
and and8926(N15234,N15239,in2);
and and8927(N15235,R0,N15240);
and and8928(N15236,R2,N15241);
and and8934(N15249,N15253,N15254);
and and8935(N15250,N15255,N15256);
and and8936(N15251,in2,N15257);
and and8937(N15252,N15258,R2);
and and8943(N15265,N15269,N15270);
and and8944(N15266,N15271,in1);
and and8945(N15267,N15272,N15273);
and and8946(N15268,N15274,R2);
and and8952(N15281,N15285,N15286);
and and8953(N15282,N15287,in1);
and and8954(N15283,N15288,N15289);
and and8955(N15284,N15290,N15291);
and and8961(N15297,N15301,N15302);
and and8962(N15298,N15303,N15304);
and and8963(N15299,N15305,R0);
and and8964(N15300,N15306,N15307);
and and8970(N15313,N15317,N15318);
and and8971(N15314,N15319,N15320);
and and8972(N15315,N15321,N15322);
and and8973(N15316,R1,N15323);
and and8979(N15329,N15333,N15334);
and and8980(N15330,N15335,N15336);
and and8981(N15331,in2,N15337);
and and8982(N15332,N15338,N15339);
and and8988(N15345,N15349,N15350);
and and8989(N15346,N15351,N15352);
and and8990(N15347,R0,N15353);
and and8991(N15348,N15354,N15355);
and and8997(N15360,N15364,N15365);
and and8998(N15361,in0,in2);
and and8999(N15362,N15366,R1);
and and9000(N15363,N15367,R3);
and and9006(N15375,N15379,N15380);
and and9007(N15376,N15381,in1);
and and9008(N15377,N15382,N15383);
and and9009(N15378,R2,N15384);
and and9015(N15390,N15394,N15395);
and and9016(N15391,N15396,N15397);
and and9017(N15392,N15398,N15399);
and and9018(N15393,R2,N15400);
and and9024(N15405,N15409,N15410);
and and9025(N15406,in0,in1);
and and9026(N15407,in2,N15411);
and and9027(N15408,N15412,N15413);
and and9033(N15420,N15424,N15425);
and and9034(N15421,N15426,in1);
and and9035(N15422,N15427,R0);
and and9036(N15423,N15428,N15429);
and and9042(N15435,N15439,N15440);
and and9043(N15436,N15441,in1);
and and9044(N15437,in2,N15442);
and and9045(N15438,N15443,R2);
and and9051(N15450,N15454,N15455);
and and9052(N15451,N15456,N15457);
and and9053(N15452,in2,R0);
and and9054(N15453,N15458,N15459);
and and9060(N15465,N15469,N15470);
and and9061(N15466,N15471,N15472);
and and9062(N15467,N15473,N15474);
and and9063(N15468,R1,R3);
and and9069(N15480,N15484,N15485);
and and9070(N15481,N15486,in1);
and and9071(N15482,N15487,R1);
and and9072(N15483,R2,N15488);
and and9078(N15495,N15499,N15500);
and and9079(N15496,N15501,N15502);
and and9080(N15497,in2,R0);
and and9081(N15498,N15503,R3);
and and9087(N15510,N15514,N15515);
and and9088(N15511,N15516,in1);
and and9089(N15512,N15517,N15518);
and and9090(N15513,R1,R3);
and and9096(N15525,N15529,N15530);
and and9097(N15526,N15531,in2);
and and9098(N15527,N15532,R1);
and and9099(N15528,N15533,R3);
and and9105(N15540,N15544,N15545);
and and9106(N15541,N15546,in1);
and and9107(N15542,N15547,N15548);
and and9108(N15543,N15549,R2);
and and9114(N15555,N15559,N15560);
and and9115(N15556,in1,in2);
and and9116(N15557,R0,N15561);
and and9117(N15558,R2,R3);
and and9123(N15569,N15573,N15574);
and and9124(N15570,N15575,in2);
and and9125(N15571,N15576,N15577);
and and9126(N15572,R2,R3);
and and9132(N15583,N15587,N15588);
and and9133(N15584,N15589,N15590);
and and9134(N15585,R0,R1);
and and9135(N15586,R2,N15591);
and and9141(N15597,N15601,N15602);
and and9142(N15598,N15603,in1);
and and9143(N15599,N15604,R0);
and and9144(N15600,R1,R2);
and and9150(N15611,N15615,N15616);
and and9151(N15612,N15617,N15618);
and and9152(N15613,N15619,R0);
and and9153(N15614,N15620,R2);
and and9159(N15625,N15629,N15630);
and and9160(N15626,N15631,in1);
and and9161(N15627,N15632,R0);
and and9162(N15628,N15633,R2);
and and9168(N15639,N15643,N15644);
and and9169(N15640,N15645,in1);
and and9170(N15641,in2,N15646);
and and9171(N15642,R2,R3);
and and9177(N15653,N15657,N15658);
and and9178(N15654,in0,in1);
and and9179(N15655,N15659,N15660);
and and9180(N15656,N15661,R3);
and and9186(N15667,N15671,N15672);
and and9187(N15668,N15673,N15674);
and and9188(N15669,R0,R1);
and and9189(N15670,N15675,R3);
and and9195(N15681,N15685,N15686);
and and9196(N15682,N15687,N15688);
and and9197(N15683,in2,R1);
and and9198(N15684,R2,N15689);
and and9204(N15695,N15699,N15700);
and and9205(N15696,N15701,in1);
and and9206(N15697,N15702,N15703);
and and9207(N15698,R1,R2);
and and9213(N15709,N15713,N15714);
and and9214(N15710,N15715,N15716);
and and9215(N15711,N15717,R0);
and and9216(N15712,N15718,N15719);
and and9222(N15723,N15727,N15728);
and and9223(N15724,in0,N15729);
and and9224(N15725,in2,R0);
and and9225(N15726,R1,N15730);
and and9231(N15737,N15741,N15742);
and and9232(N15738,N15743,N15744);
and and9233(N15739,N15745,N15746);
and and9234(N15740,R2,N15747);
and and9240(N15751,N15755,N15756);
and and9241(N15752,in0,in1);
and and9242(N15753,in2,N15757);
and and9243(N15754,N15758,R2);
and and9249(N15765,N15769,N15770);
and and9250(N15766,N15771,N15772);
and and9251(N15767,N15773,R0);
and and9252(N15768,R1,R2);
and and9258(N15779,N15783,N15784);
and and9259(N15780,in0,N15785);
and and9260(N15781,in2,N15786);
and and9261(N15782,R1,R3);
and and9267(N15793,N15797,N15798);
and and9268(N15794,in1,in2);
and and9269(N15795,N15799,N15800);
and and9270(N15796,N15801,R3);
and and9276(N15807,N15811,N15812);
and and9277(N15808,in1,in2);
and and9278(N15809,N15813,N15814);
and and9279(N15810,R2,N15815);
and and9285(N15821,N15825,N15826);
and and9286(N15822,in0,N15827);
and and9287(N15823,N15828,N15829);
and and9288(N15824,R1,N15830);
and and9294(N15835,N15839,N15840);
and and9295(N15836,N15841,N15842);
and and9296(N15837,in2,R0);
and and9297(N15838,N15843,R2);
and and9303(N15849,N15853,N15854);
and and9304(N15850,N15855,N15856);
and and9305(N15851,N15857,R0);
and and9306(N15852,R1,R2);
and and9312(N15863,N15867,N15868);
and and9313(N15864,N15869,N15870);
and and9314(N15865,R0,N15871);
and and9315(N15866,N15872,N15873);
and and9321(N15877,N15881,N15882);
and and9322(N15878,in1,in2);
and and9323(N15879,N15883,R1);
and and9324(N15880,R2,N15884);
and and9330(N15891,N15895,N15896);
and and9331(N15892,N15897,in2);
and and9332(N15893,N15898,N15899);
and and9333(N15894,R2,N15900);
and and9339(N15905,N15909,N15910);
and and9340(N15906,in1,in2);
and and9341(N15907,R0,N15911);
and and9342(N15908,N15912,R3);
and and9348(N15919,N15923,N15924);
and and9349(N15920,N15925,in1);
and and9350(N15921,in2,R0);
and and9351(N15922,N15926,N15927);
and and9357(N15933,N15937,N15938);
and and9358(N15934,in1,in2);
and and9359(N15935,N15939,R1);
and and9360(N15936,N15940,R3);
and and9366(N15947,N15951,N15952);
and and9367(N15948,N15953,in2);
and and9368(N15949,N15954,N15955);
and and9369(N15950,N15956,R3);
and and9375(N15961,N15965,N15966);
and and9376(N15962,in0,N15967);
and and9377(N15963,in2,R0);
and and9378(N15964,N15968,N15969);
and and9384(N15975,N15979,N15980);
and and9385(N15976,N15981,in1);
and and9386(N15977,in2,R0);
and and9387(N15978,N15982,N15983);
and and9393(N15989,N15993,N15994);
and and9394(N15990,N15995,in1);
and and9395(N15991,N15996,N15997);
and and9396(N15992,N15998,R2);
and and9402(N16003,N16007,N16008);
and and9403(N16004,in1,N16009);
and and9404(N16005,N16010,N16011);
and and9405(N16006,R2,N16012);
and and9411(N16017,N16021,N16022);
and and9412(N16018,in0,N16023);
and and9413(N16019,in2,N16024);
and and9414(N16020,R2,N16025);
and and9420(N16031,N16035,N16036);
and and9421(N16032,N16037,N16038);
and and9422(N16033,in2,R0);
and and9423(N16034,N16039,N16040);
and and9429(N16045,N16049,N16050);
and and9430(N16046,N16051,in1);
and and9431(N16047,N16052,R0);
and and9432(N16048,N16053,N16054);
and and9438(N16059,N16063,N16064);
and and9439(N16060,in1,N16065);
and and9440(N16061,N16066,N16067);
and and9441(N16062,R2,R3);
and and9447(N16073,N16077,N16078);
and and9448(N16074,in0,in1);
and and9449(N16075,in2,N16079);
and and9450(N16076,N16080,N16081);
and and9456(N16087,N16091,N16092);
and and9457(N16088,N16093,N16094);
and and9458(N16089,R0,R1);
and and9459(N16090,N16095,R3);
and and9465(N16101,N16105,N16106);
and and9466(N16102,in1,N16107);
and and9467(N16103,R0,N16108);
and and9468(N16104,R2,R3);
and and9474(N16114,N16118,N16119);
and and9475(N16115,in1,N16120);
and and9476(N16116,R0,R1);
and and9477(N16117,R2,N16121);
and and9483(N16127,N16131,N16132);
and and9484(N16128,N16133,N16134);
and and9485(N16129,in2,N16135);
and and9486(N16130,R1,R2);
and and9492(N16140,N16144,N16145);
and and9493(N16141,N16146,N16147);
and and9494(N16142,N16148,R1);
and and9495(N16143,R2,R3);
and and9501(N16153,N16157,N16158);
and and9502(N16154,in0,in1);
and and9503(N16155,N16159,R1);
and and9504(N16156,R2,N16160);
and and9510(N16166,N16170,N16171);
and and9511(N16167,N16172,N16173);
and and9512(N16168,N16174,R0);
and and9513(N16169,R2,R3);
and and9519(N16179,N16183,N16184);
and and9520(N16180,N16185,in2);
and and9521(N16181,R0,R1);
and and9522(N16182,N16186,R3);
and and9528(N16192,N16196,N16197);
and and9529(N16193,N16198,N16199);
and and9530(N16194,N16200,R1);
and and9531(N16195,R2,R3);
and and9537(N16205,N16209,N16210);
and and9538(N16206,in1,in2);
and and9539(N16207,N16211,R1);
and and9540(N16208,R2,N16212);
and and9546(N16218,N16222,N16223);
and and9547(N16219,in0,in1);
and and9548(N16220,N16224,R1);
and and9549(N16221,R2,N16225);
and and9555(N16231,N16235,N16236);
and and9556(N16232,in0,in1);
and and9557(N16233,in2,N16237);
and and9558(N16234,N16238,R2);
and and9564(N16244,N16248,N16249);
and and9565(N16245,N16250,N16251);
and and9566(N16246,R0,R1);
and and9567(N16247,N16252,R3);
and and9573(N16257,N16261,N16262);
and and9574(N16258,N16263,in1);
and and9575(N16259,N16264,R0);
and and9576(N16260,R1,R2);
and and9582(N16270,N16274,N16275);
and and9583(N16271,N16276,in1);
and and9584(N16272,N16277,N16278);
and and9585(N16273,R1,R2);
and and9591(N16283,N16287,N16288);
and and9592(N16284,in1,N16289);
and and9593(N16285,R0,R1);
and and9594(N16286,R2,R3);
and and9600(N16296,N16300,N16301);
and and9601(N16297,N16302,in1);
and and9602(N16298,in2,N16303);
and and9603(N16299,N16304,R2);
and and9609(N16309,N16313,N16314);
and and9610(N16310,in0,in1);
and and9611(N16311,N16315,R0);
and and9612(N16312,R1,N16316);
and and9618(N16322,N16326,N16327);
and and9619(N16323,in0,N16328);
and and9620(N16324,N16329,R0);
and and9621(N16325,N16330,N16331);
and and9627(N16335,N16339,N16340);
and and9628(N16336,in0,N16341);
and and9629(N16337,N16342,N16343);
and and9630(N16338,N16344,R2);
and and9636(N16348,N16352,N16353);
and and9637(N16349,N16354,N16355);
and and9638(N16350,in2,N16356);
and and9639(N16351,N16357,R2);
and and9645(N16361,N16365,N16366);
and and9646(N16362,in0,in1);
and and9647(N16363,in2,R0);
and and9648(N16364,N16367,R3);
and and9654(N16374,N16378,N16379);
and and9655(N16375,in0,N16380);
and and9656(N16376,in2,N16381);
and and9657(N16377,R1,N16382);
and and9663(N16387,N16391,N16392);
and and9664(N16388,N16393,in2);
and and9665(N16389,R0,N16394);
and and9666(N16390,R2,N16395);
and and9672(N16400,N16404,N16405);
and and9673(N16401,in0,N16406);
and and9674(N16402,in2,N16407);
and and9675(N16403,N16408,R2);
and and9681(N16413,N16417,N16418);
and and9682(N16414,in0,in2);
and and9683(N16415,R0,N16419);
and and9684(N16416,R2,R3);
and and9690(N16425,N16429,N16430);
and and9691(N16426,N16431,in1);
and and9692(N16427,in2,R0);
and and9693(N16428,N16432,R2);
and and9699(N16437,N16441,N16442);
and and9700(N16438,in0,in1);
and and9701(N16439,in2,N16443);
and and9702(N16440,R2,R3);
and and9708(N16449,N16453,N16454);
and and9709(N16450,N16455,in1);
and and9710(N16451,in2,R0);
and and9711(N16452,R2,R3);
and and9717(N16461,N16465,N16466);
and and9718(N16462,in1,in2);
and and9719(N16463,N16467,N16468);
and and9720(N16464,R2,R3);
and and9726(N16473,N16477,N16478);
and and9727(N16474,in0,in2);
and and9728(N16475,R0,R1);
and and9729(N16476,R2,N16479);
and and9735(N16485,N16489,N16490);
and and9736(N16486,in0,in1);
and and9737(N16487,in2,N16491);
and and9738(N16488,R1,R2);
and and9744(N16497,N16501,N16502);
and and9745(N16498,N16503,in1);
and and9746(N16499,in2,N16504);
and and9747(N16500,R1,R2);
and and9753(N16509,N16513,N16514);
and and9754(N16510,in0,in1);
and and9755(N16511,N16515,R0);
and and9756(N16512,N16516,R2);
and and9762(N16521,N16525,N16526);
and and9763(N16522,in1,in2);
and and9764(N16523,R0,N16527);
and and9765(N16524,R2,N16528);
and and9771(N16533,N16537,N16538);
and and9772(N16534,N16539,in2);
and and9773(N16535,R0,N16540);
and and9774(N16536,N16541,R3);
and and9780(N16545,N16549,N16550);
and and9781(N16546,in0,in1);
and and9782(N16547,in2,N16551);
and and9783(N16548,N16552,R3);
and and9789(N16557,N16561,N16562);
and and9790(N16558,in0,N16563);
and and9791(N16559,R0,N16564);
and and9792(N16560,R2,R3);
and and9798(N16569,N16573,N16574);
and and9799(N16570,N16575,N16576);
and and9800(N16571,in2,R1);
and and9801(N16572,R2,R3);
and and9807(N16581,N16585,N16586);
and and9808(N16582,in0,N16587);
and and9809(N16583,in2,R0);
and and9810(N16584,N16588,N16589);
and and9816(N16593,N16597,N16598);
and and9817(N16594,in0,in1);
and and9818(N16595,N16599,R0);
and and9819(N16596,N16600,N16601);
and and9825(N16605,N16609,N16610);
and and9826(N16606,N16611,in1);
and and9827(N16607,in2,R0);
and and9828(N16608,N16612,N16613);
and and9834(N16617,N16621,N16622);
and and9835(N16618,N16623,N16624);
and and9836(N16619,in2,R0);
and and9837(N16620,R1,R3);
and and9843(N16629,N16633,N16634);
and and9844(N16630,N16635,N16636);
and and9845(N16631,N16637,R1);
and and9846(N16632,R2,R3);
and and9852(N16641,N16645,N16646);
and and9853(N16642,in0,in1);
and and9854(N16643,in2,N16647);
and and9855(N16644,R1,R2);
and and9861(N16653,N16657,N16658);
and and9862(N16654,N16659,in1);
and and9863(N16655,N16660,R1);
and and9864(N16656,R2,N16661);
and and9870(N16665,N16669,N16670);
and and9871(N16666,in0,in1);
and and9872(N16667,N16671,N16672);
and and9873(N16668,R1,R2);
and and9879(N16677,N16681,N16682);
and and9880(N16678,in0,N16683);
and and9881(N16679,in2,N16684);
and and9882(N16680,R1,R3);
and and9888(N16689,N16693,N16694);
and and9889(N16690,in0,N16695);
and and9890(N16691,in2,R0);
and and9891(N16692,R1,R2);
and and9897(N16701,N16705,N16706);
and and9898(N16702,in0,in2);
and and9899(N16703,R0,N16707);
and and9900(N16704,R2,R3);
and and9906(N16713,N16717,N16718);
and and9907(N16714,in0,in2);
and and9908(N16715,R0,N16719);
and and9909(N16716,N16720,N16721);
and and9915(N16725,N16729,N16730);
and and9916(N16726,in0,in1);
and and9917(N16727,N16731,R0);
and and9918(N16728,N16732,N16733);
and and9924(N16737,N16741,N16742);
and and9925(N16738,N16743,in1);
and and9926(N16739,in2,R0);
and and9927(N16740,R1,N16744);
and and9933(N16749,N16753,N16754);
and and9934(N16750,in0,in1);
and and9935(N16751,in2,R0);
and and9936(N16752,N16755,N16756);
and and9942(N16761,N16765,N16766);
and and9943(N16762,in0,in2);
and and9944(N16763,R0,N16767);
and and9945(N16764,N16768,R3);
and and9951(N16773,N16777,N16778);
and and9952(N16774,N16779,in1);
and and9953(N16775,in2,R0);
and and9954(N16776,N16780,R3);
and and9960(N16785,N16789,N16790);
and and9961(N16786,in0,in1);
and and9962(N16787,N16791,N16792);
and and9963(N16788,R2,R3);
and and9969(N16797,N16801,N16802);
and and9970(N16798,in0,in1);
and and9971(N16799,in2,N16803);
and and9972(N16800,N16804,R2);
and and9978(N16809,N16813,N16814);
and and9979(N16810,in0,in1);
and and9980(N16811,in2,R0);
and and9981(N16812,R1,N16815);
and and9987(N16821,N16825,N16826);
and and9988(N16822,in0,in1);
and and9989(N16823,N16827,R0);
and and9990(N16824,R1,R2);
and and9996(N16833,N16837,N16838);
and and9997(N16834,in0,in1);
and and9998(N16835,in2,R0);
and and9999(N16836,N16839,R3);
and and10005(N16845,N16849,N16850);
and and10006(N16846,in0,in1);
and and10007(N16847,in2,N16851);
and and10008(N16848,N16852,R2);
and and10014(N16857,N16861,N16862);
and and10015(N16858,in0,N16863);
and and10016(N16859,in2,R0);
and and10017(N16860,R2,N16864);
and and10023(N16869,N16873,N16874);
and and10024(N16870,in0,in1);
and and10025(N16871,N16875,R0);
and and10026(N16872,R2,N16876);
and and10032(N16881,N16885,N16886);
and and10033(N16882,N16887,in1);
and and10034(N16883,N16888,R0);
and and10035(N16884,R1,R2);
and and10041(N16893,N16897,N16898);
and and10042(N16894,in0,in2);
and and10043(N16895,N16899,N16900);
and and10044(N16896,R2,R3);
and and10050(N16904,N16908,N16909);
and and10051(N16905,in0,in1);
and and10052(N16906,N16910,R1);
and and10053(N16907,R2,R3);
and and10059(N16915,N16919,N16920);
and and10060(N16916,N16921,in1);
and and10061(N16917,in2,R0);
and and10062(N16918,R1,R2);
and and10068(N16926,N16930,N16931);
and and10069(N16927,in0,in1);
and and10070(N16928,in2,R0);
and and10071(N16929,N16932,R2);
and and10077(N16937,N16941,N16942);
and and10078(N16938,in1,N16943);
and and10079(N16939,R0,N16944);
and and10080(N16940,R2,R3);
and and10086(N16948,N16952,N16953);
and and10087(N16949,in0,in1);
and and10088(N16950,in2,R0);
and and10089(N16951,R2,R3);
and and10095(N16958,N16962,N16963);
and and10096(N16959,in0,in1);
and and10097(N16960,in2,N16964);
and and10098(N16961,R1,R2);
and and10104(N16968,N16972,N16973);
and and10105(N16969,in0,in1);
and and10106(N16970,in2,R0);
and and10107(N16971,R2,R3);
and and10113(N16978,N16982,N16983);
and and10114(N16979,in0,in1);
and and10115(N16980,in2,R0);
and and10116(N16981,N16984,R3);
and and10122(N16988,N16992,N16993);
and and10123(N16989,in0,in1);
and and10124(N16990,in2,R0);
and and10125(N16991,R1,R3);
and and10131(N16998,N17002,N17003);
and and10132(N16999,in0,in1);
and and10133(N17000,N17004,R1);
and and10134(N17001,R2,R3);
and and10140(N17008,N17012,N17013);
and and10141(N17009,N17014,in1);
and and10142(N17010,in2,R0);
and and10143(N17011,R1,R2);
and and10149(N17018,N17022,N17023);
and and10150(N17019,in0,in1);
and and10151(N17020,R0,R1);
and and10152(N17021,R2,R3);
and and10158(N17028,N17032,N17033);
and and10159(N17029,in2,N17034);
and and10160(N17030,N17035,N17036);
and and10161(N17031,N17037,N17038);
and and10166(N17044,N17048,N17049);
and and10167(N17045,N17050,N17051);
and and10168(N17046,N17052,R3);
and and10169(N17047,N17053,N17054);
and and10174(N17060,N17064,N17065);
and and10175(N17061,N17066,N17067);
and and10176(N17062,R1,N17068);
and and10177(N17063,N17069,N17070);
and and10182(N17075,N17079,in1);
and and10183(N17076,N17080,N17081);
and and10184(N17077,N17082,N17083);
and and10185(N17078,N17084,N17085);
and and10190(N17090,N17094,N17095);
and and10191(N17091,in2,N17096);
and and10192(N17092,N17097,N17098);
and and10193(N17093,N17099,R4);
and and10198(N17105,N17109,in0);
and and10199(N17106,N17110,N17111);
and and10200(N17107,R2,N17112);
and and10201(N17108,N17113,N17114);
and and10206(N17120,N17124,N17125);
and and10207(N17121,N17126,R0);
and and10208(N17122,N17127,N17128);
and and10209(N17123,N17129,N17130);
and and10214(N17135,N17139,N17140);
and and10215(N17136,in2,N17141);
and and10216(N17137,N17142,R3);
and and10217(N17138,N17143,N17144);
and and10222(N17150,N17154,N17155);
and and10223(N17151,N17156,N17157);
and and10224(N17152,N17158,R2);
and and10225(N17153,N17159,N17160);
and and10230(N17165,N17169,N17170);
and and10231(N17166,N17171,in2);
and and10232(N17167,N17172,N17173);
and and10233(N17168,N17174,N17175);
and and10238(N17180,N17184,N17185);
and and10239(N17181,N17186,N17187);
and and10240(N17182,N17188,N17189);
and and10241(N17183,N17190,R5);
and and10246(N17195,N17199,N17200);
and and10247(N17196,N17201,N17202);
and and10248(N17197,N17203,N17204);
and and10249(N17198,R3,N17205);
and and10254(N17210,N17214,N17215);
and and10255(N17211,N17216,N17217);
and and10256(N17212,R2,N17218);
and and10257(N17213,R4,N17219);
and and10262(N17225,N17229,N17230);
and and10263(N17226,in1,in2);
and and10264(N17227,N17231,N17232);
and and10265(N17228,N17233,N17234);
and and10270(N17240,N17244,N17245);
and and10271(N17241,N17246,R1);
and and10272(N17242,N17247,N17248);
and and10273(N17243,N17249,N17250);
and and10278(N17255,N17259,N17260);
and and10279(N17256,N17261,N17262);
and and10280(N17257,N17263,R2);
and and10281(N17258,N17264,N17265);
and and10286(N17270,N17274,N17275);
and and10287(N17271,N17276,N17277);
and and10288(N17272,R0,N17278);
and and10289(N17273,N17279,N17280);
and and10294(N17285,N17289,N17290);
and and10295(N17286,N17291,R0);
and and10296(N17287,N17292,N17293);
and and10297(N17288,N17294,N17295);
and and10302(N17300,N17304,in1);
and and10303(N17301,N17305,N17306);
and and10304(N17302,R1,N17307);
and and10305(N17303,R3,N17308);
and and10310(N17314,N17318,in0);
and and10311(N17315,R0,N17319);
and and10312(N17316,N17320,N17321);
and and10313(N17317,N17322,N17323);
and and10318(N17328,N17332,N17333);
and and10319(N17329,in2,R0);
and and10320(N17330,N17334,N17335);
and and10321(N17331,R4,N17336);
and and10326(N17342,N17346,in2);
and and10327(N17343,R0,N17347);
and and10328(N17344,N17348,N17349);
and and10329(N17345,N17350,R5);
and and10334(N17356,N17360,N17361);
and and10335(N17357,N17362,R1);
and and10336(N17358,R2,R3);
and and10337(N17359,N17363,N17364);
and and10342(N17370,N17374,in0);
and and10343(N17371,N17375,R0);
and and10344(N17372,N17376,R2);
and and10345(N17373,N17377,N17378);
and and10350(N17384,N17388,in0);
and and10351(N17385,N17389,N17390);
and and10352(N17386,N17391,R2);
and and10353(N17387,N17392,N17393);
and and10358(N17398,N17402,in1);
and and10359(N17399,N17403,N17404);
and and10360(N17400,N17405,R2);
and and10361(N17401,N17406,N17407);
and and10366(N17412,N17416,N17417);
and and10367(N17413,N17418,N17419);
and and10368(N17414,N17420,N17421);
and and10369(N17415,N17422,R3);
and and10374(N17426,N17430,in0);
and and10375(N17427,N17431,R0);
and and10376(N17428,N17432,N17433);
and and10377(N17429,R3,N17434);
and and10382(N17440,N17444,in0);
and and10383(N17441,N17445,N17446);
and and10384(N17442,N17447,R2);
and and10385(N17443,R3,N17448);
and and10390(N17454,N17458,in0);
and and10391(N17455,N17459,N17460);
and and10392(N17456,N17461,N17462);
and and10393(N17457,N17463,R5);
and and10398(N17468,N17472,N17473);
and and10399(N17469,N17474,N17475);
and and10400(N17470,R2,N17476);
and and10401(N17471,N17477,N17478);
and and10406(N17482,N17486,N17487);
and and10407(N17483,N17488,N17489);
and and10408(N17484,N17490,R3);
and and10409(N17485,N17491,N17492);
and and10414(N17496,N17500,N17501);
and and10415(N17497,in2,N17502);
and and10416(N17498,N17503,N17504);
and and10417(N17499,R3,R4);
and and10422(N17510,N17514,N17515);
and and10423(N17511,N17516,N17517);
and and10424(N17512,R2,R3);
and and10425(N17513,R4,N17518);
and and10430(N17524,N17528,N17529);
and and10431(N17525,N17530,N17531);
and and10432(N17526,R1,N17532);
and and10433(N17527,R3,N17533);
and and10438(N17538,N17542,N17543);
and and10439(N17539,N17544,N17545);
and and10440(N17540,N17546,R3);
and and10441(N17541,R4,N17547);
and and10446(N17552,N17556,N17557);
and and10447(N17553,N17558,in2);
and and10448(N17554,R1,N17559);
and and10449(N17555,N17560,R5);
and and10454(N17566,N17570,in0);
and and10455(N17567,N17571,N17572);
and and10456(N17568,N17573,N17574);
and and10457(N17569,R3,N17575);
and and10462(N17580,N17584,N17585);
and and10463(N17581,in2,N17586);
and and10464(N17582,N17587,N17588);
and and10465(N17583,R3,N17589);
and and10470(N17594,N17598,N17599);
and and10471(N17595,in1,N17600);
and and10472(N17596,N17601,N17602);
and and10473(N17597,N17603,R3);
and and10478(N17608,N17612,in0);
and and10479(N17609,N17613,N17614);
and and10480(N17610,R2,N17615);
and and10481(N17611,R4,N17616);
and and10486(N17622,N17626,N17627);
and and10487(N17623,N17628,R0);
and and10488(N17624,R2,N17629);
and and10489(N17625,N17630,N17631);
and and10494(N17636,N17640,in0);
and and10495(N17637,N17641,N17642);
and and10496(N17638,N17643,R3);
and and10497(N17639,N17644,R5);
and and10502(N17650,N17654,N17655);
and and10503(N17651,in1,N17656);
and and10504(N17652,N17657,R3);
and and10505(N17653,N17658,R5);
and and10510(N17664,N17668,N17669);
and and10511(N17665,in1,N17670);
and and10512(N17666,N17671,R2);
and and10513(N17667,N17672,N17673);
and and10518(N17678,N17682,N17683);
and and10519(N17679,N17684,N17685);
and and10520(N17680,R1,R2);
and and10521(N17681,N17686,N17687);
and and10526(N17692,N17696,in2);
and and10527(N17693,R0,N17697);
and and10528(N17694,N17698,N17699);
and and10529(N17695,N17700,N17701);
and and10534(N17706,N17710,in0);
and and10535(N17707,in1,N17711);
and and10536(N17708,N17712,N17713);
and and10537(N17709,N17714,R5);
and and10542(N17720,N17724,N17725);
and and10543(N17721,N17726,N17727);
and and10544(N17722,N17728,R2);
and and10545(N17723,R3,R4);
and and10550(N17734,N17738,in0);
and and10551(N17735,N17739,N17740);
and and10552(N17736,N17741,N17742);
and and10553(N17737,R3,N17743);
and and10558(N17748,N17752,in0);
and and10559(N17749,N17753,N17754);
and and10560(N17750,R2,N17755);
and and10561(N17751,R4,N17756);
and and10566(N17762,N17766,N17767);
and and10567(N17763,N17768,N17769);
and and10568(N17764,R2,R3);
and and10569(N17765,N17770,R5);
and and10574(N17775,N17779,in0);
and and10575(N17776,in1,R1);
and and10576(N17777,N17780,N17781);
and and10577(N17778,N17782,N17783);
and and10582(N17788,N17792,in0);
and and10583(N17789,in1,in2);
and and10584(N17790,N17793,N17794);
and and10585(N17791,N17795,N17796);
and and10590(N17801,N17805,in0);
and and10591(N17802,N17806,R0);
and and10592(N17803,R1,R2);
and and10593(N17804,N17807,N17808);
and and10598(N17814,N17818,in0);
and and10599(N17815,in1,N17819);
and and10600(N17816,N17820,R2);
and and10601(N17817,N17821,N17822);
and and10606(N17827,N17831,in0);
and and10607(N17828,in1,N17832);
and and10608(N17829,R0,N17833);
and and10609(N17830,N17834,N17835);
and and10614(N17840,N17844,in1);
and and10615(N17841,in2,N17845);
and and10616(N17842,R1,R2);
and and10617(N17843,N17846,N17847);
and and10622(N17853,N17857,in0);
and and10623(N17854,N17858,N17859);
and and10624(N17855,R2,N17860);
and and10625(N17856,N17861,R5);
and and10630(N17866,N17870,in0);
and and10631(N17867,in1,N17871);
and and10632(N17868,R0,N17872);
and and10633(N17869,R2,N17873);
and and10638(N17879,N17883,N17884);
and and10639(N17880,in2,R0);
and and10640(N17881,N17885,R2);
and and10641(N17882,N17886,N17887);
and and10646(N17892,N17896,in0);
and and10647(N17893,in1,N17897);
and and10648(N17894,R2,R3);
and and10649(N17895,N17898,N17899);
and and10654(N17905,N17909,N17910);
and and10655(N17906,N17911,in2);
and and10656(N17907,N17912,R1);
and and10657(N17908,N17913,R5);
and and10662(N17918,N17922,in2);
and and10663(N17919,R0,N17923);
and and10664(N17920,N17924,N17925);
and and10665(N17921,R4,N17926);
and and10670(N17931,N17935,in0);
and and10671(N17932,N17936,R0);
and and10672(N17933,N17937,N17938);
and and10673(N17934,N17939,R4);
and and10678(N17944,N17948,N17949);
and and10679(N17945,N17950,R1);
and and10680(N17946,R2,N17951);
and and10681(N17947,R4,N17952);
and and10686(N17957,N17961,in0);
and and10687(N17958,in1,in2);
and and10688(N17959,N17962,N17963);
and and10689(N17960,N17964,N17965);
and and10694(N17970,N17974,N17975);
and and10695(N17971,N17976,R0);
and and10696(N17972,N17977,N17978);
and and10697(N17973,R3,R4);
and and10702(N17983,N17987,in0);
and and10703(N17984,N17988,N17989);
and and10704(N17985,N17990,N17991);
and and10705(N17986,R3,N17992);
and and10710(N17996,N18000,in1);
and and10711(N17997,N18001,N18002);
and and10712(N17998,R2,N18003);
and and10713(N17999,N18004,N18005);
and and10718(N18009,N18013,N18014);
and and10719(N18010,N18015,R0);
and and10720(N18011,N18016,R2);
and and10721(N18012,N18017,R5);
and and10726(N18022,N18026,in0);
and and10727(N18023,N18027,N18028);
and and10728(N18024,R0,N18029);
and and10729(N18025,R2,R5);
and and10734(N18035,N18039,N18040);
and and10735(N18036,in2,R0);
and and10736(N18037,N18041,R2);
and and10737(N18038,N18042,R5);
and and10742(N18048,N18052,N18053);
and and10743(N18049,in1,R0);
and and10744(N18050,N18054,R2);
and and10745(N18051,N18055,R5);
and and10750(N18061,N18065,in0);
and and10751(N18062,N18066,R0);
and and10752(N18063,N18067,N18068);
and and10753(N18064,N18069,N18070);
and and10758(N18074,N18078,N18079);
and and10759(N18075,N18080,R0);
and and10760(N18076,N18081,N18082);
and and10761(N18077,R4,R5);
and and10766(N18087,N18091,N18092);
and and10767(N18088,N18093,in2);
and and10768(N18089,R0,N18094);
and and10769(N18090,R3,N18095);
and and10774(N18100,N18104,in0);
and and10775(N18101,N18105,N18106);
and and10776(N18102,N18107,R2);
and and10777(N18103,R3,R4);
and and10782(N18113,N18117,in0);
and and10783(N18114,N18118,R0);
and and10784(N18115,N18119,R3);
and and10785(N18116,R4,N18120);
and and10790(N18126,N18130,in0);
and and10791(N18127,N18131,R0);
and and10792(N18128,N18132,R2);
and and10793(N18129,N18133,R4);
and and10798(N18139,N18143,N18144);
and and10799(N18140,in1,R0);
and and10800(N18141,N18145,R2);
and and10801(N18142,N18146,R4);
and and10806(N18152,N18156,N18157);
and and10807(N18153,in1,N18158);
and and10808(N18154,R0,N18159);
and and10809(N18155,N18160,N18161);
and and10814(N18165,N18169,N18170);
and and10815(N18166,R0,R1);
and and10816(N18167,N18171,N18172);
and and10817(N18168,R4,R5);
and and10822(N18178,N18182,in0);
and and10823(N18179,N18183,R1);
and and10824(N18180,N18184,R3);
and and10825(N18181,N18185,N18186);
and and10830(N18191,N18195,in1);
and and10831(N18192,N18196,N18197);
and and10832(N18193,N18198,R3);
and and10833(N18194,R4,N18199);
and and10838(N18204,N18208,in0);
and and10839(N18205,N18209,N18210);
and and10840(N18206,N18211,R3);
and and10841(N18207,R4,N18212);
and and10846(N18217,N18221,in1);
and and10847(N18218,in2,N18222);
and and10848(N18219,R1,N18223);
and and10849(N18220,N18224,R5);
and and10854(N18230,N18234,N18235);
and and10855(N18231,N18236,N18237);
and and10856(N18232,R1,R2);
and and10857(N18233,R3,N18238);
and and10862(N18243,N18247,in0);
and and10863(N18244,in1,N18248);
and and10864(N18245,N18249,N18250);
and and10865(N18246,N18251,R3);
and and10870(N18256,N18260,in0);
and and10871(N18257,in1,N18261);
and and10872(N18258,N18262,N18263);
and and10873(N18259,R3,N18264);
and and10878(N18269,N18273,N18274);
and and10879(N18270,N18275,N18276);
and and10880(N18271,N18277,R3);
and and10881(N18272,R4,R5);
and and10886(N18282,N18286,in0);
and and10887(N18283,N18287,N18288);
and and10888(N18284,R0,N18289);
and and10889(N18285,R2,N18290);
and and10894(N18295,N18299,N18300);
and and10895(N18296,N18301,R0);
and and10896(N18297,N18302,R3);
and and10897(N18298,N18303,R5);
and and10902(N18308,N18312,in1);
and and10903(N18309,N18313,R0);
and and10904(N18310,N18314,R3);
and and10905(N18311,N18315,N18316);
and and10910(N18321,N18325,N18326);
and and10911(N18322,in2,R0);
and and10912(N18323,N18327,R3);
and and10913(N18324,N18328,N18329);
and and10918(N18334,N18338,N18339);
and and10919(N18335,in1,R0);
and and10920(N18336,R1,N18340);
and and10921(N18337,R3,N18341);
and and10926(N18347,N18351,N18352);
and and10927(N18348,in2,R0);
and and10928(N18349,R1,R3);
and and10929(N18350,N18353,N18354);
and and10934(N18360,N18364,in0);
and and10935(N18361,N18365,R0);
and and10936(N18362,R1,N18366);
and and10937(N18363,R3,N18367);
and and10942(N18373,N18377,N18378);
and and10943(N18374,N18379,N18380);
and and10944(N18375,N18381,R2);
and and10945(N18376,R3,N18382);
and and10950(N18386,N18390,in0);
and and10951(N18387,N18391,in2);
and and10952(N18388,N18392,R3);
and and10953(N18389,N18393,R5);
and and10958(N18399,N18403,N18404);
and and10959(N18400,N18405,in2);
and and10960(N18401,N18406,R2);
and and10961(N18402,N18407,R4);
and and10966(N18412,N18416,N18417);
and and10967(N18413,N18418,N18419);
and and10968(N18414,R2,R3);
and and10969(N18415,N18420,R5);
and and10974(N18425,N18429,N18430);
and and10975(N18426,N18431,R0);
and and10976(N18427,R1,R3);
and and10977(N18428,N18432,R5);
and and10982(N18438,N18442,in0);
and and10983(N18439,N18443,N18444);
and and10984(N18440,R2,N18445);
and and10985(N18441,N18446,R5);
and and10990(N18451,N18455,in0);
and and10991(N18452,in1,R0);
and and10992(N18453,N18456,N18457);
and and10993(N18454,R3,N18458);
and and10998(N18464,N18468,N18469);
and and10999(N18465,in1,N18470);
and and11000(N18466,R2,R3);
and and11001(N18467,N18471,R5);
and and11006(N18477,N18481,in1);
and and11007(N18478,N18482,R1);
and and11008(N18479,N18483,R3);
and and11009(N18480,R4,N18484);
and and11014(N18490,N18494,in2);
and and11015(N18491,N18495,N18496);
and and11016(N18492,N18497,R3);
and and11017(N18493,N18498,N18499);
and and11022(N18503,N18507,N18508);
and and11023(N18504,N18509,R0);
and and11024(N18505,N18510,N18511);
and and11025(N18506,R4,R5);
and and11030(N18516,N18520,in0);
and and11031(N18517,N18521,in2);
and and11032(N18518,N18522,N18523);
and and11033(N18519,R3,R4);
and and11038(N18529,N18533,N18534);
and and11039(N18530,N18535,N18536);
and and11040(N18531,N18537,R3);
and and11041(N18532,R4,R5);
and and11046(N18542,N18546,in0);
and and11047(N18543,N18547,R0);
and and11048(N18544,N18548,R2);
and and11049(N18545,N18549,N18550);
and and11054(N18555,N18559,in0);
and and11055(N18556,N18560,R0);
and and11056(N18557,N18561,R2);
and and11057(N18558,N18562,N18563);
and and11062(N18568,N18572,in0);
and and11063(N18569,N18573,N18574);
and and11064(N18570,R0,N18575);
and and11065(N18571,N18576,N18577);
and and11070(N18581,N18585,N18586);
and and11071(N18582,N18587,N18588);
and and11072(N18583,R0,N18589);
and and11073(N18584,R2,R5);
and and11078(N18594,N18598,in0);
and and11079(N18595,in1,N18599);
and and11080(N18596,R0,R1);
and and11081(N18597,R2,N18600);
and and11086(N18606,N18610,in1);
and and11087(N18607,N18611,R0);
and and11088(N18608,R1,R2);
and and11089(N18609,N18612,N18613);
and and11094(N18618,N18622,in0);
and and11095(N18619,N18623,N18624);
and and11096(N18620,R1,R2);
and and11097(N18621,R3,R4);
and and11102(N18630,N18634,in0);
and and11103(N18631,in1,in2);
and and11104(N18632,R0,R2);
and and11105(N18633,N18635,N18636);
and and11110(N18642,N18646,in0);
and and11111(N18643,N18647,N18648);
and and11112(N18644,R1,R2);
and and11113(N18645,N18649,R5);
and and11118(N18654,N18658,N18659);
and and11119(N18655,N18660,R0);
and and11120(N18656,R1,R3);
and and11121(N18657,R4,N18661);
and and11126(N18666,N18670,in1);
and and11127(N18667,in2,N18671);
and and11128(N18668,R1,R2);
and and11129(N18669,N18672,R5);
and and11134(N18678,N18682,in1);
and and11135(N18679,in2,R0);
and and11136(N18680,R1,N18683);
and and11137(N18681,N18684,R4);
and and11142(N18690,N18694,N18695);
and and11143(N18691,in1,in2);
and and11144(N18692,R1,N18696);
and and11145(N18693,N18697,R5);
and and11150(N18702,N18706,N18707);
and and11151(N18703,N18708,N18709);
and and11152(N18704,R1,N18710);
and and11153(N18705,R3,R5);
and and11158(N18714,N18718,N18719);
and and11159(N18715,R0,R1);
and and11160(N18716,R2,N18720);
and and11161(N18717,R4,N18721);
and and11166(N18726,N18730,in1);
and and11167(N18727,N18731,R1);
and and11168(N18728,N18732,R3);
and and11169(N18729,N18733,R5);
and and11174(N18738,N18742,N18743);
and and11175(N18739,R0,R1);
and and11176(N18740,R2,R3);
and and11177(N18741,N18744,N18745);
and and11182(N18750,N18754,N18755);
and and11183(N18751,R0,N18756);
and and11184(N18752,R2,N18757);
and and11185(N18753,R4,R5);
and and11190(N18762,N18766,N18767);
and and11191(N18763,in1,R1);
and and11192(N18764,N18768,R3);
and and11193(N18765,R4,R5);
and and11198(N18774,N18778,in1);
and and11199(N18775,R0,R1);
and and11200(N18776,N18779,N18780);
and and11201(N18777,R4,N18781);
and and11206(N18786,N18790,in0);
and and11207(N18787,N18791,R0);
and and11208(N18788,R1,R2);
and and11209(N18789,N18792,R4);
and and11214(N18798,N18802,in0);
and and11215(N18799,in2,N18803);
and and11216(N18800,R2,R3);
and and11217(N18801,R4,N18804);
and and11222(N18810,N18814,in1);
and and11223(N18811,in2,N18815);
and and11224(N18812,R2,R3);
and and11225(N18813,R4,N18816);
and and11230(N18822,N18826,in0);
and and11231(N18823,N18827,N18828);
and and11232(N18824,R0,R1);
and and11233(N18825,R2,R3);
and and11238(N18834,N18838,in0);
and and11239(N18835,in1,N18839);
and and11240(N18836,R1,N18840);
and and11241(N18837,R3,N18841);
and and11246(N18846,N18850,in0);
and and11247(N18847,N18851,N18852);
and and11248(N18848,N18853,N18854);
and and11249(N18849,R3,R4);
and and11254(N18858,N18862,N18863);
and and11255(N18859,in2,N18864);
and and11256(N18860,R2,R3);
and and11257(N18861,R4,N18865);
and and11262(N18870,N18874,in0);
and and11263(N18871,N18875,N18876);
and and11264(N18872,R2,R3);
and and11265(N18873,R4,N18877);
and and11270(N18882,N18886,in0);
and and11271(N18883,N18887,N18888);
and and11272(N18884,R2,N18889);
and and11273(N18885,N18890,R5);
and and11278(N18894,N18898,in0);
and and11279(N18895,in1,in2);
and and11280(N18896,N18899,N18900);
and and11281(N18897,R2,N18901);
and and11286(N18906,N18910,in0);
and and11287(N18907,N18911,N18912);
and and11288(N18908,N18913,R3);
and and11289(N18909,R4,R5);
and and11294(N18918,N18922,in1);
and and11295(N18919,in2,R0);
and and11296(N18920,R2,N18923);
and and11297(N18921,N18924,N18925);
and and11302(N18930,N18934,in0);
and and11303(N18931,N18935,N18936);
and and11304(N18932,R0,R2);
and and11305(N18933,N18937,R4);
and and11310(N18942,N18946,in1);
and and11311(N18943,in2,N18947);
and and11312(N18944,N18948,R2);
and and11313(N18945,N18949,R4);
and and11318(N18954,N18958,in0);
and and11319(N18955,N18959,R0);
and and11320(N18956,R1,N18960);
and and11321(N18957,R3,N18961);
and and11326(N18966,N18970,N18971);
and and11327(N18967,N18972,in2);
and and11328(N18968,R1,R2);
and and11329(N18969,N18973,R5);
and and11334(N18978,N18982,in0);
and and11335(N18979,in2,N18983);
and and11336(N18980,R1,N18984);
and and11337(N18981,N18985,R5);
and and11342(N18990,N18994,N18995);
and and11343(N18991,N18996,N18997);
and and11344(N18992,R1,R2);
and and11345(N18993,R4,N18998);
and and11350(N19002,N19006,in0);
and and11351(N19003,in2,R0);
and and11352(N19004,N19007,N19008);
and and11353(N19005,N19009,N19010);
and and11358(N19014,N19018,in0);
and and11359(N19015,in1,N19019);
and and11360(N19016,R0,R1);
and and11361(N19017,R2,N19020);
and and11366(N19026,N19030,N19031);
and and11367(N19027,in2,N19032);
and and11368(N19028,R2,N19033);
and and11369(N19029,R4,N19034);
and and11374(N19038,N19042,in1);
and and11375(N19039,in2,R0);
and and11376(N19040,R1,N19043);
and and11377(N19041,N19044,R4);
and and11382(N19050,N19054,in0);
and and11383(N19051,in1,N19055);
and and11384(N19052,R0,R1);
and and11385(N19053,N19056,N19057);
and and11390(N19062,N19066,in0);
and and11391(N19063,N19067,in2);
and and11392(N19064,N19068,N19069);
and and11393(N19065,N19070,R3);
and and11398(N19074,N19078,N19079);
and and11399(N19075,N19080,in2);
and and11400(N19076,R0,R1);
and and11401(N19077,N19081,R4);
and and11406(N19086,N19090,in0);
and and11407(N19087,N19091,in2);
and and11408(N19088,R0,N19092);
and and11409(N19089,R3,N19093);
and and11414(N19098,N19102,in0);
and and11415(N19099,in1,N19103);
and and11416(N19100,N19104,R3);
and and11417(N19101,N19105,R5);
and and11422(N19110,N19114,in0);
and and11423(N19111,in1,R0);
and and11424(N19112,R1,N19115);
and and11425(N19113,R3,N19116);
and and11430(N19122,N19126,in1);
and and11431(N19123,N19127,N19128);
and and11432(N19124,R2,R3);
and and11433(N19125,N19129,R5);
and and11438(N19134,N19138,in0);
and and11439(N19135,N19139,R0);
and and11440(N19136,R1,N19140);
and and11441(N19137,R3,N19141);
and and11446(N19146,N19150,N19151);
and and11447(N19147,in1,in2);
and and11448(N19148,R0,R1);
and and11449(N19149,N19152,R3);
and and11454(N19158,N19162,in1);
and and11455(N19159,N19163,R1);
and and11456(N19160,R2,R3);
and and11457(N19161,N19164,R5);
and and11462(N19169,N19173,N19174);
and and11463(N19170,in1,N19175);
and and11464(N19171,R0,R1);
and and11465(N19172,R2,R5);
and and11470(N19180,N19184,N19185);
and and11471(N19181,in2,R0);
and and11472(N19182,N19186,R3);
and and11473(N19183,R4,N19187);
and and11478(N19191,N19195,in0);
and and11479(N19192,in1,in2);
and and11480(N19193,R0,R2);
and and11481(N19194,N19196,N19197);
and and11486(N19202,N19206,in0);
and and11487(N19203,in1,R0);
and and11488(N19204,N19207,R2);
and and11489(N19205,N19208,R4);
and and11494(N19213,N19217,N19218);
and and11495(N19214,in2,R0);
and and11496(N19215,R1,R2);
and and11497(N19216,R3,N19219);
and and11502(N19224,N19228,in0);
and and11503(N19225,N19229,R0);
and and11504(N19226,N19230,R2);
and and11505(N19227,R3,R4);
and and11510(N19235,N19239,in0);
and and11511(N19236,N19240,in2);
and and11512(N19237,N19241,R1);
and and11513(N19238,R2,R4);
and and11518(N19246,N19250,N19251);
and and11519(N19247,N19252,R1);
and and11520(N19248,R2,N19253);
and and11521(N19249,R4,R5);
and and11526(N19257,N19261,N19262);
and and11527(N19258,in1,N19263);
and and11528(N19259,R1,R3);
and and11529(N19260,N19264,R5);
and and11534(N19268,N19272,N19273);
and and11535(N19269,N19274,R0);
and and11536(N19270,R1,R3);
and and11537(N19271,R4,R5);
and and11542(N19279,N19283,in0);
and and11543(N19280,in2,R1);
and and11544(N19281,N19284,R3);
and and11545(N19282,N19285,R5);
and and11550(N19290,N19294,in1);
and and11551(N19291,in2,R0);
and and11552(N19292,N19295,R2);
and and11553(N19293,N19296,R5);
and and11558(N19301,N19305,N19306);
and and11559(N19302,in2,R0);
and and11560(N19303,R1,R2);
and and11561(N19304,R3,R4);
and and11566(N19312,N19316,in0);
and and11567(N19313,in1,in2);
and and11568(N19314,R0,N19317);
and and11569(N19315,R2,N19318);
and and11574(N19323,N19327,in0);
and and11575(N19324,N19328,R0);
and and11576(N19325,R1,R2);
and and11577(N19326,N19329,N19330);
and and11582(N19334,N19338,in0);
and and11583(N19335,N19339,R0);
and and11584(N19336,N19340,R2);
and and11585(N19337,R3,R4);
and and11590(N19345,N19349,N19350);
and and11591(N19346,in1,R0);
and and11592(N19347,N19351,N19352);
and and11593(N19348,R4,R5);
and and11598(N19356,N19360,in0);
and and11599(N19357,in1,in2);
and and11600(N19358,R0,N19361);
and and11601(N19359,R2,N19362);
and and11606(N19367,N19371,N19372);
and and11607(N19368,R0,R1);
and and11608(N19369,R2,N19373);
and and11609(N19370,R4,N19374);
and and11614(N19378,N19382,in0);
and and11615(N19379,in2,N19383);
and and11616(N19380,N19384,R2);
and and11617(N19381,R4,N19385);
and and11622(N19389,N19393,N19394);
and and11623(N19390,N19395,R0);
and and11624(N19391,R1,R2);
and and11625(N19392,R4,R5);
and and11630(N19400,N19404,N19405);
and and11631(N19401,R0,R1);
and and11632(N19402,R2,N19406);
and and11633(N19403,N19407,R5);
and and11638(N19411,N19415,in0);
and and11639(N19412,N19416,N19417);
and and11640(N19413,N19418,R1);
and and11641(N19414,R2,R4);
and and11646(N19422,N19426,N19427);
and and11647(N19423,in2,N19428);
and and11648(N19424,R1,R2);
and and11649(N19425,R4,R5);
and and11654(N19433,N19437,in1);
and and11655(N19434,N19438,R0);
and and11656(N19435,N19439,R3);
and and11657(N19436,R4,R5);
and and11662(N19444,N19448,in0);
and and11663(N19445,N19449,in2);
and and11664(N19446,R0,N19450);
and and11665(N19447,R3,R5);
and and11670(N19455,N19459,in0);
and and11671(N19456,in1,R0);
and and11672(N19457,N19460,R3);
and and11673(N19458,N19461,R5);
and and11678(N19466,N19470,N19471);
and and11679(N19467,in1,in2);
and and11680(N19468,R0,N19472);
and and11681(N19469,R3,R5);
and and11686(N19477,N19481,in0);
and and11687(N19478,in2,R0);
and and11688(N19479,N19482,R2);
and and11689(N19480,N19483,R4);
and and11694(N19488,N19492,in0);
and and11695(N19489,in1,R0);
and and11696(N19490,N19493,R2);
and and11697(N19491,N19494,R4);
and and11702(N19499,N19503,N19504);
and and11703(N19500,in1,in2);
and and11704(N19501,N19505,R1);
and and11705(N19502,R3,R4);
and and11710(N19510,N19514,in0);
and and11711(N19511,N19515,N19516);
and and11712(N19512,R0,R2);
and and11713(N19513,N19517,R4);
and and11718(N19521,N19525,in0);
and and11719(N19522,N19526,R0);
and and11720(N19523,N19527,R2);
and and11721(N19524,R3,R4);
and and11726(N19532,N19536,in0);
and and11727(N19533,in1,N19537);
and and11728(N19534,N19538,R3);
and and11729(N19535,R4,R5);
and and11734(N19543,N19547,in1);
and and11735(N19544,in2,R0);
and and11736(N19545,R1,N19548);
and and11737(N19546,R4,N19549);
and and11742(N19554,N19558,in1);
and and11743(N19555,in2,N19559);
and and11744(N19556,R1,R3);
and and11745(N19557,R4,N19560);
and and11750(N19565,N19569,in0);
and and11751(N19566,in1,in2);
and and11752(N19567,R0,R1);
and and11753(N19568,N19570,R5);
and and11758(N19576,N19580,in0);
and and11759(N19577,N19581,R1);
and and11760(N19578,N19582,R3);
and and11761(N19579,R4,R5);
and and11766(N19586,N19590,in0);
and and11767(N19587,in1,N19591);
and and11768(N19588,R1,R2);
and and11769(N19589,R3,N19592);
and and11774(N19596,N19600,in1);
and and11775(N19597,in2,R0);
and and11776(N19598,R1,R3);
and and11777(N19599,R4,N19601);
and and11782(N19606,N19610,in0);
and and11783(N19607,N19611,R0);
and and11784(N19608,R1,N19612);
and and11785(N19609,R3,R4);
and and11790(N19616,N19620,in0);
and and11791(N19617,R0,R1);
and and11792(N19618,N19621,R3);
and and11793(N19619,R4,N19622);
and and11798(N19626,N19630,in0);
and and11799(N19627,N19631,in2);
and and11800(N19628,R2,N19632);
and and11801(N19629,R4,R5);
and and11806(N19636,N19640,in0);
and and11807(N19637,R0,R1);
and and11808(N19638,N19641,R3);
and and11809(N19639,N19642,R5);
and and11814(N19646,N19650,in0);
and and11815(N19647,in1,N19651);
and and11816(N19648,R1,N19652);
and and11817(N19649,R3,R5);
and and11822(N19656,N19660,in1);
and and11823(N19657,in2,R0);
and and11824(N19658,R1,R2);
and and11825(N19659,N19661,R4);
and and11830(N19666,N19670,in1);
and and11831(N19667,in2,R0);
and and11832(N19668,R1,R2);
and and11833(N19669,N19671,N19672);
and and11838(N19676,N19680,in0);
and and11839(N19677,in1,N19681);
and and11840(N19678,R0,R1);
and and11841(N19679,R2,N19682);
and and11846(N19686,N19690,in0);
and and11847(N19687,in1,in2);
and and11848(N19688,R0,R1);
and and11849(N19689,R2,N19691);
and and11854(N19696,N19700,in0);
and and11855(N19697,in1,in2);
and and11856(N19698,R0,R1);
and and11857(N19699,R2,R3);
and and11862(N19706,N19710,N19711);
and and11863(N19707,R0,R1);
and and11864(N19708,N19712,R3);
and and11865(N19709,R4,R5);
and and11870(N19716,N19720,in0);
and and11871(N19717,in1,N19721);
and and11872(N19718,R1,R2);
and and11873(N19719,R4,R5);
and and11878(N19726,N19730,in0);
and and11879(N19727,in1,in2);
and and11880(N19728,N19731,R2);
and and11881(N19729,R3,R4);
and and11886(N19736,N19740,in0);
and and11887(N19737,N19741,in2);
and and11888(N19738,R0,R1);
and and11889(N19739,R2,R4);
and and11894(N19746,N19750,in0);
and and11895(N19747,N19751,R0);
and and11896(N19748,R1,R2);
and and11897(N19749,R3,N19752);
and and11902(N19756,N19760,in0);
and and11903(N19757,R0,R1);
and and11904(N19758,R2,N19761);
and and11905(N19759,N19762,R5);
and and11910(N19766,N19770,N19771);
and and11911(N19767,in1,in2);
and and11912(N19768,R2,R3);
and and11913(N19769,R4,R5);
and and11918(N19775,N19779,in0);
and and11919(N19776,in2,R0);
and and11920(N19777,R1,R2);
and and11921(N19778,R4,N19780);
and and11926(N19784,N19788,in0);
and and11927(N19785,in1,R0);
and and11928(N19786,R1,R2);
and and11929(N19787,N19789,R4);
and and11934(N19793,N19797,in0);
and and11935(N19794,N19798,R0);
and and11936(N19795,R2,R3);
and and11937(N19796,R4,R5);
and and11942(N19802,N19806,N19807);
and and11943(N19803,in2,R0);
and and11944(N19804,R2,R3);
and and11945(N19805,R4,R5);
and and11950(N19811,N19815,in0);
and and11951(N19812,in1,in2);
and and11952(N19813,R2,R3);
and and11953(N19814,R4,R5);
and and11958(N19820,N19824,in0);
and and11959(N19821,N19825,in2);
and and11960(N19822,R1,R2);
and and11961(N19823,R4,R5);
and and11966(N19829,N19833,in0);
and and11967(N19830,in2,R1);
and and11968(N19831,R2,N19834);
and and11969(N19832,R4,R5);
and and11974(N19838,N19842,in0);
and and11975(N19839,in1,R0);
and and11976(N19840,R1,N19843);
and and11977(N19841,R3,R4);
and and11982(N19847,N19851,in0);
and and11983(N19848,in1,in2);
and and11984(N19849,R0,R2);
and and11985(N19850,R3,R5);
and and11990(N19855,N19859,R0);
and and11991(N19856,N19860,N19861);
and and11992(N19857,N19862,N19863);
and and11993(N19858,N19864,N19865);
and and11997(N19869,N19873,N19874);
and and11998(N19870,N19875,N19876);
and and11999(N19871,N19877,N19878);
and and12000(N19872,R6,N19879);
and and12004(N19883,in0,N19887);
and and12005(N19884,N19888,N19889);
and and12006(N19885,N19890,N19891);
and and12007(N19886,N19892,N19893);
and and12011(N19897,N19901,N19902);
and and12012(N19898,N19903,N19904);
and and12013(N19899,N19905,R5);
and and12014(N19900,N19906,N19907);
and and12018(N19911,in0,N19915);
and and12019(N19912,N19916,N19917);
and and12020(N19913,N19918,N19919);
and and12021(N19914,N19920,N19921);
and and12025(N19925,in0,N19929);
and and12026(N19926,N19930,N19931);
and and12027(N19927,N19932,R4);
and and12028(N19928,N19933,N19934);
and and12032(N19938,N19942,R0);
and and12033(N19939,N19943,N19944);
and and12034(N19940,R4,N19945);
and and12035(N19941,N19946,N19947);
and and12039(N19951,N19955,N19956);
and and12040(N19952,N19957,N19958);
and and12041(N19953,R3,R5);
and and12042(N19954,N19959,N19960);
and and12046(N19964,in0,in1);
and and12047(N19965,R0,N19968);
and and12048(N19966,N19969,N19970);
and and12049(N19967,N19971,N19972);
and and12053(N19976,in0,N19980);
and and12054(N19977,N19981,R2);
and and12055(N19978,N19982,N19983);
and and12056(N19979,N19984,R7);
and and12060(N19988,in0,N19992);
and and12061(N19989,R1,R2);
and and12062(N19990,N19993,N19994);
and and12063(N19991,N19995,N19996);
and and12067(N20000,in0,N20004);
and and12068(N20001,N20005,R2);
and and12069(N20002,N20006,R5);
and and12070(N20003,N20007,N20008);
and and12074(N20012,N20016,N20017);
and and12075(N20013,R1,N20018);
and and12076(N20014,R3,R4);
and and12077(N20015,N20019,N20020);
and and12081(N20024,in0,N20028);
and and12082(N20025,N20029,R1);
and and12083(N20026,N20030,N20031);
and and12084(N20027,R5,N20032);
and and12088(N20036,in1,N20040);
and and12089(N20037,N20041,R1);
and and12090(N20038,N20042,N20043);
and and12091(N20039,R5,N20044);
and and12095(N20048,N20052,N20053);
and and12096(N20049,N20054,R2);
and and12097(N20050,N20055,R4);
and and12098(N20051,R6,N20056);
and and12102(N20060,in0,N20064);
and and12103(N20061,N20065,R2);
and and12104(N20062,N20066,R5);
and and12105(N20063,N20067,N20068);
and and12109(N20072,in0,N20076);
and and12110(N20073,N20077,N20078);
and and12111(N20074,R3,R4);
and and12112(N20075,N20079,N20080);
and and12116(N20084,in0,N20088);
and and12117(N20085,R0,R1);
and and12118(N20086,N20089,N20090);
and and12119(N20087,N20091,R7);
and and12123(N20095,in0,in2);
and and12124(N20096,N20099,N20100);
and and12125(N20097,N20101,R5);
and and12126(N20098,N20102,R7);
and and12130(N20106,in0,N20110);
and and12131(N20107,N20111,R2);
and and12132(N20108,N20112,N20113);
and and12133(N20109,R6,R7);
and and12137(N20117,in1,R0);
and and12138(N20118,N20121,N20122);
and and12139(N20119,R4,N20123);
and and12140(N20120,R6,N20124);
and and12144(N20128,in0,R0);
and and12145(N20129,N20132,N20133);
and and12146(N20130,R4,N20134);
and and12147(N20131,R6,N20135);
and and12151(N20139,N20143,R0);
and and12152(N20140,R1,N20144);
and and12153(N20141,N20145,R4);
and and12154(N20142,N20146,R7);
and and12158(N20150,in0,R0);
and and12159(N20151,N20154,R3);
and and12160(N20152,N20155,N20156);
and and12161(N20153,N20157,R7);
and and12165(N20161,in0,R0);
and and12166(N20162,N20165,N20166);
and and12167(N20163,N20167,N20168);
and and12168(N20164,R6,R7);
and and12172(N20172,N20176,N20177);
and and12173(N20173,N20178,R2);
and and12174(N20174,R4,N20179);
and and12175(N20175,R6,R7);
and and12179(N20183,in0,N20187);
and and12180(N20184,R0,N20188);
and and12181(N20185,N20189,R4);
and and12182(N20186,R5,N20190);
and and12186(N20194,in0,R0);
and and12187(N20195,R1,N20198);
and and12188(N20196,N20199,R5);
and and12189(N20197,N20200,N20201);
and and12193(N20205,in0,N20209);
and and12194(N20206,R1,R3);
and and12195(N20207,N20210,N20211);
and and12196(N20208,N20212,R7);
and and12200(N20216,in0,N20220);
and and12201(N20217,N20221,N20222);
and and12202(N20218,R2,R4);
and and12203(N20219,N20223,R7);
and and12207(N20227,in0,N20231);
and and12208(N20228,R1,R2);
and and12209(N20229,R3,N20232);
and and12210(N20230,R6,N20233);
and and12214(N20237,in0,R0);
and and12215(N20238,N20241,R3);
and and12216(N20239,R4,N20242);
and and12217(N20240,N20243,R7);
and and12221(N20247,N20251,in2);
and and12222(N20248,R1,R3);
and and12223(N20249,R4,R5);
and and12224(N20250,N20252,N20253);
and and12228(N20257,in0,R1);
and and12229(N20258,R2,R3);
and and12230(N20259,N20261,R5);
and and12231(N20260,N20262,N20263);
and and12235(N20267,in0,N20271);
and and12236(N20268,R0,N20272);
and and12237(N20269,R3,N20273);
and and12238(N20270,R6,R7);
and and12242(N20277,in1,N20281);
and and12243(N20278,N20282,N20283);
and and12244(N20279,R3,R4);
and and12245(N20280,R5,R6);
and and12249(N20287,in0,R0);
and and12250(N20288,R1,N20291);
and and12251(N20289,R3,N20292);
and and12252(N20290,N20293,R7);
and and12256(N20297,N20301,in1);
and and12257(N20298,R0,N20302);
and and12258(N20299,R2,R4);
and and12259(N20300,N20303,R7);
and and12263(N20307,in0,in1);
and and12264(N20308,N20311,N20312);
and and12265(N20309,N20313,R2);
and and12266(N20310,R4,R7);
and and12270(N20317,in0,N20321);
and and12271(N20318,R0,N20322);
and and12272(N20319,R3,N20323);
and and12273(N20320,R6,R7);
and and12277(N20327,in0,in1);
and and12278(N20328,R0,N20331);
and and12279(N20329,N20332,R4);
and and12280(N20330,R5,N20333);
and and12284(N20337,in1,in2);
and and12285(N20338,R0,R2);
and and12286(N20339,R3,N20341);
and and12287(N20340,N20342,R6);
and and12291(N20346,R0,R1);
and and12292(N20347,R2,R3);
and and12293(N20348,N20350,R5);
and and12294(N20349,R6,N20351);
and and12298(N20355,in0,N20359);
and and12299(N20356,R2,R3);
and and12300(N20357,R4,R5);
and and12301(N20358,R6,N20360);
and and12305(N20364,in0,in1);
and and12306(N20365,in2,R2);
and and12307(N20366,R3,R4);
and and12308(N20367,N20368,N20369);
and and12312(N20373,in0,R0);
and and12313(N20374,R1,R2);
and and12314(N20375,R3,N20377);
and and12315(N20376,R5,R7);
and and12319(N20381,in0,in1);
and and12320(N20382,R0,R1);
and and12321(N20383,R3,R4);
and and12322(N20384,R6,N20385);
and and12326(N20389,in0,R0);
and and12327(N20390,R1,R3);
and and12328(N20391,R4,R5);
and and12329(N20392,R6,N20393);
and and12333(N20397,R1,R3);
and and12334(N20398,R4,R5);
and and12335(N20399,N20400,N20401);
and and8884(N15153,N15160,N15161);
and and8885(N15154,N15162,N15163);
and and8893(N15171,R4,N15178);
and and8894(N15172,N15179,N15180);
and and8902(N15188,N15195,N15196);
and and8903(N15189,N15197,R7);
and and8911(N15205,N15210,N15211);
and and8912(N15206,N15212,N15213);
and and8920(N15221,N15226,N15227);
and and8921(N15222,N15228,N15229);
and and8929(N15237,N15242,N15243);
and and8930(N15238,N15244,N15245);
and and8938(N15253,N15259,N15260);
and and8939(N15254,R6,N15261);
and and8947(N15269,R3,N15275);
and and8948(N15270,N15276,N15277);
and and8956(N15285,N15292,R4);
and and8957(N15286,R5,N15293);
and and8965(N15301,N15308,N15309);
and and8966(N15302,R6,R7);
and and8974(N15317,R3,N15324);
and and8975(N15318,N15325,R7);
and and8983(N15333,R3,N15340);
and and8984(N15334,R5,N15341);
and and8992(N15349,R4,R5);
and and8993(N15350,N15356,R7);
and and9001(N15364,N15368,N15369);
and and9002(N15365,N15370,N15371);
and and9010(N15379,N15385,R5);
and and9011(N15380,N15386,R7);
and and9019(N15394,R4,R5);
and and9020(N15395,N15401,R7);
and and9028(N15409,R4,N15414);
and and9029(N15410,N15415,N15416);
and and9037(N15424,N15430,R5);
and and9038(N15425,N15431,R7);
and and9046(N15439,N15444,N15445);
and and9047(N15440,R5,N15446);
and and9055(N15454,R4,N15460);
and and9056(N15455,R6,N15461);
and and9064(N15469,R4,R5);
and and9065(N15470,N15475,N15476);
and and9073(N15484,R4,N15489);
and and9074(N15485,N15490,N15491);
and and9082(N15499,R4,N15504);
and and9083(N15500,N15505,N15506);
and and9091(N15514,N15519,N15520);
and and9092(N15515,R6,N15521);
and and9100(N15529,N15534,N15535);
and and9101(N15530,N15536,R7);
and and9109(N15544,N15550,R4);
and and9110(N15545,N15551,R7);
and and9118(N15559,N15562,N15563);
and and9119(N15560,N15564,N15565);
and and9127(N15573,R4,R5);
and and9128(N15574,N15578,N15579);
and and9136(N15587,N15592,R5);
and and9137(N15588,R6,N15593);
and and9145(N15601,N15605,N15606);
and and9146(N15602,R6,N15607);
and and9154(N15615,N15621,R4);
and and9155(N15616,R6,R7);
and and9163(N15629,R3,N15634);
and and9164(N15630,N15635,R7);
and and9172(N15643,N15647,N15648);
and and9173(N15644,N15649,R7);
and and9181(N15657,R4,N15662);
and and9182(N15658,N15663,R7);
and and9190(N15671,N15676,R5);
and and9191(N15672,R6,N15677);
and and9199(N15685,N15690,R5);
and and9200(N15686,R6,N15691);
and and9208(N15699,N15704,R5);
and and9209(N15700,R6,N15705);
and and9217(N15713,R3,R5);
and and9218(N15714,R6,R7);
and and9226(N15727,R4,N15731);
and and9227(N15728,N15732,N15733);
and and9235(N15741,R4,R5);
and and9236(N15742,R6,R7);
and and9244(N15755,N15759,N15760);
and and9245(N15756,R5,N15761);
and and9253(N15769,R3,N15774);
and and9254(N15770,N15775,R7);
and and9262(N15783,R4,N15787);
and and9263(N15784,N15788,N15789);
and and9271(N15797,N15802,R5);
and and9272(N15798,N15803,R7);
and and9280(N15811,N15816,N15817);
and and9281(N15812,R6,R7);
and and9289(N15825,R3,N15831);
and and9290(N15826,R5,R6);
and and9298(N15839,N15844,N15845);
and and9299(N15840,R5,R6);
and and9307(N15853,R3,R4);
and and9308(N15854,N15858,N15859);
and and9316(N15867,R4,R5);
and and9317(N15868,R6,R7);
and and9325(N15881,R4,N15885);
and and9326(N15882,N15886,N15887);
and and9334(N15895,R4,R5);
and and9335(N15896,R6,N15901);
and and9343(N15909,R4,N15913);
and and9344(N15910,N15914,N15915);
and and9352(N15923,N15928,N15929);
and and9353(N15924,R6,R7);
and and9361(N15937,N15941,N15942);
and and9362(N15938,R6,N15943);
and and9370(N15951,R4,R5);
and and9371(N15952,R6,N15957);
and and9379(N15965,N15970,R4);
and and9380(N15966,R5,N15971);
and and9388(N15979,N15984,R4);
and and9389(N15980,R5,N15985);
and and9397(N15993,R3,R4);
and and9398(N15994,N15999,R6);
and and9406(N16007,N16013,R5);
and and9407(N16008,R6,R7);
and and9415(N16021,R4,N16026);
and and9416(N16022,R6,N16027);
and and9424(N16035,R3,N16041);
and and9425(N16036,R5,R6);
and and9433(N16049,R3,N16055);
and and9434(N16050,R5,R7);
and and9442(N16063,N16068,N16069);
and and9443(N16064,R6,R7);
and and9451(N16077,R3,N16082);
and and9452(N16078,R5,N16083);
and and9460(N16091,N16096,R5);
and and9461(N16092,N16097,R7);
and and9469(N16105,R4,R5);
and and9470(N16106,N16109,N16110);
and and9478(N16118,R4,R5);
and and9479(N16119,N16122,N16123);
and and9487(N16131,R3,R4);
and and9488(N16132,N16136,R7);
and and9496(N16144,R4,R5);
and and9497(N16145,N16149,R7);
and and9505(N16157,N16161,R5);
and and9506(N16158,N16162,R7);
and and9514(N16170,N16175,R5);
and and9515(N16171,R6,R7);
and and9523(N16183,R4,N16187);
and and9524(N16184,R6,N16188);
and and9532(N16196,N16201,R5);
and and9533(N16197,R6,R7);
and and9541(N16209,N16213,R5);
and and9542(N16210,R6,N16214);
and and9550(N16222,N16226,R5);
and and9551(N16223,R6,N16227);
and and9559(N16235,R3,R5);
and and9560(N16236,N16239,N16240);
and and9568(N16248,R4,N16253);
and and9569(N16249,R6,R7);
and and9577(N16261,R4,N16265);
and and9578(N16262,R6,N16266);
and and9586(N16274,R3,R4);
and and9587(N16275,R5,N16279);
and and9595(N16287,R4,N16290);
and and9596(N16288,N16291,N16292);
and and9604(N16300,N16305,R4);
and and9605(N16301,R5,R6);
and and9613(N16313,N16317,R4);
and and9614(N16314,R5,N16318);
and and9622(N16326,R3,R4);
and and9623(N16327,R5,R7);
and and9631(N16339,R3,R5);
and and9632(N16340,R6,R7);
and and9640(N16352,R3,R4);
and and9641(N16353,R5,R6);
and and9649(N16365,N16368,N16369);
and and9650(N16366,R6,N16370);
and and9658(N16378,R3,R4);
and and9659(N16379,N16383,R7);
and and9667(N16391,R4,R5);
and and9668(N16392,R6,N16396);
and and9676(N16404,R3,N16409);
and and9677(N16405,R5,R6);
and and9685(N16417,R4,R5);
and and9686(N16418,N16420,N16421);
and and9694(N16429,R3,R4);
and and9695(N16430,R5,N16433);
and and9703(N16441,N16444,R5);
and and9704(N16442,N16445,R7);
and and9712(N16453,N16456,R5);
and and9713(N16454,N16457,R7);
and and9721(N16465,R4,R5);
and and9722(N16466,N16469,R7);
and and9730(N16477,N16480,R5);
and and9731(N16478,R6,N16481);
and and9739(N16489,N16492,N16493);
and and9740(N16490,R6,R7);
and and9748(N16501,R3,N16505);
and and9749(N16502,R6,R7);
and and9757(N16513,N16517,R5);
and and9758(N16514,R6,R7);
and and9766(N16525,N16529,R5);
and and9767(N16526,R6,R7);
and and9775(N16537,R4,R5);
and and9776(N16538,R6,R7);
and and9784(N16549,N16553,R5);
and and9785(N16550,R6,R7);
and and9793(N16561,N16565,R5);
and and9794(N16562,R6,R7);
and and9802(N16573,N16577,R5);
and and9803(N16574,R6,R7);
and and9811(N16585,R3,R5);
and and9812(N16586,R6,R7);
and and9820(N16597,R3,R5);
and and9821(N16598,R6,R7);
and and9829(N16609,R3,R5);
and and9830(N16610,R6,R7);
and and9838(N16621,R4,R5);
and and9839(N16622,N16625,R7);
and and9847(N16633,R4,R5);
and and9848(N16634,R6,R7);
and and9856(N16645,N16648,R4);
and and9857(N16646,N16649,R7);
and and9865(N16657,R4,R5);
and and9866(N16658,R6,R7);
and and9874(N16669,N16673,R4);
and and9875(N16670,R6,R7);
and and9883(N16681,N16685,R5);
and and9884(N16682,R6,R7);
and and9892(N16693,R3,R4);
and and9893(N16694,N16696,N16697);
and and9901(N16705,R4,N16708);
and and9902(N16706,R6,N16709);
and and9910(N16717,R4,R5);
and and9911(N16718,R6,R7);
and and9919(N16729,R4,R5);
and and9920(N16730,R6,R7);
and and9928(N16741,R3,N16745);
and and9929(N16742,R6,R7);
and and9937(N16753,R3,N16757);
and and9938(N16754,R6,R7);
and and9946(N16765,R4,R5);
and and9947(N16766,N16769,R7);
and and9955(N16777,R4,R5);
and and9956(N16778,N16781,R7);
and and9964(N16789,N16793,R5);
and and9965(N16790,R6,R7);
and and9973(N16801,N16805,R5);
and and9974(N16802,R6,R7);
and and9982(N16813,N16816,R5);
and and9983(N16814,N16817,R7);
and and9991(N16825,R4,N16828);
and and9992(N16826,N16829,R7);
and and10000(N16837,N16840,R5);
and and10001(N16838,N16841,R7);
and and10009(N16849,R3,N16853);
and and10010(N16850,R6,R7);
and and10018(N16861,R4,R5);
and and10019(N16862,R6,N16865);
and and10027(N16873,R4,R5);
and and10028(N16874,R6,N16877);
and and10036(N16885,R3,N16889);
and and10037(N16886,R6,R7);
and and10045(N16897,R4,R5);
and and10046(N16898,R6,R7);
and and10054(N16908,N16911,R5);
and and10055(N16909,R6,R7);
and and10063(N16919,N16922,R5);
and and10064(N16920,R6,R7);
and and10072(N16930,N16933,R4);
and and10073(N16931,R5,R6);
and and10081(N16941,R4,R5);
and and10082(N16942,R6,R7);
and and10090(N16952,R4,R5);
and and10091(N16953,N16954,R7);
and and10099(N16962,R3,R4);
and and10100(N16963,R6,R7);
and and10108(N16972,R4,N16974);
and and10109(N16973,R6,R7);
and and10117(N16982,R4,R5);
and and10118(N16983,R6,R7);
and and10126(N16992,R4,R5);
and and10127(N16993,N16994,R7);
and and10135(N17002,R4,R5);
and and10136(N17003,R6,R7);
and and10144(N17012,R3,R4);
and and10145(N17013,R5,R7);
and and10153(N17022,R4,R5);
and and10154(N17023,N17024,R7);
and and10162(N17032,N17039,N17040);
and and10170(N17048,N17055,N17056);
and and10178(N17064,N17071,R7);
and and10186(N17079,R6,N17086);
and and10194(N17094,N17100,N17101);
and and10202(N17109,N17115,N17116);
and and10210(N17124,R5,N17131);
and and10218(N17139,N17145,N17146);
and and10226(N17154,R5,N17161);
and and10234(N17169,N17176,R7);
and and10242(N17184,N17191,R7);
and and10250(N17199,N17206,R7);
and and10258(N17214,N17220,N17221);
and and10266(N17229,N17235,N17236);
and and10274(N17244,N17251,R7);
and and10282(N17259,R5,N17266);
and and10290(N17274,R5,N17281);
and and10298(N17289,R6,N17296);
and and10306(N17304,N17309,N17310);
and and10314(N17318,N17324,R7);
and and10322(N17332,N17337,N17338);
and and10330(N17346,N17351,N17352);
and and10338(N17360,N17365,N17366);
and and10346(N17374,N17379,N17380);
and and10354(N17388,R6,N17394);
and and10362(N17402,R6,N17408);
and and10370(N17416,R5,R6);
and and10378(N17430,N17435,N17436);
and and10386(N17444,N17449,N17450);
and and10394(N17458,N17464,R7);
and and10402(N17472,R6,R7);
and and10410(N17486,R6,R7);
and and10418(N17500,N17505,N17506);
and and10426(N17514,N17519,N17520);
and and10434(N17528,R6,N17534);
and and10442(N17542,R6,N17548);
and and10450(N17556,N17561,N17562);
and and10458(N17570,R6,N17576);
and and10466(N17584,R6,N17590);
and and10474(N17598,N17604,R7);
and and10482(N17612,N17617,N17618);
and and10490(N17626,R6,N17632);
and and10498(N17640,N17645,N17646);
and and10506(N17654,N17659,N17660);
and and10514(N17668,R6,N17674);
and and10522(N17682,R5,N17688);
and and10530(N17696,R6,N17702);
and and10538(N17710,N17715,N17716);
and and10546(N17724,N17729,N17730);
and and10554(N17738,N17744,R7);
and and10562(N17752,N17757,N17758);
and and10570(N17766,N17771,R7);
and and10578(N17779,N17784,R7);
and and10586(N17792,R6,N17797);
and and10594(N17805,N17809,N17810);
and and10602(N17818,N17823,R7);
and and10610(N17831,N17836,R5);
and and10618(N17844,N17848,N17849);
and and10626(N17857,R6,N17862);
and and10634(N17870,N17874,N17875);
and and10642(N17883,N17888,R7);
and and10650(N17896,N17900,N17901);
and and10658(N17909,N17914,R7);
and and10666(N17922,N17927,R7);
and and10674(N17935,N17940,R7);
and and10682(N17948,N17953,R7);
and and10690(N17961,N17966,R7);
and and10698(N17974,N17979,R7);
and and10706(N17987,R5,R7);
and and10714(N18000,R6,R7);
and and10722(N18013,R6,N18018);
and and10730(N18026,N18030,N18031);
and and10738(N18039,N18043,N18044);
and and10746(N18052,N18056,N18057);
and and10754(N18065,R5,R6);
and and10762(N18078,R6,N18083);
and and10770(N18091,N18096,R7);
and and10778(N18104,N18108,N18109);
and and10786(N18117,N18121,N18122);
and and10794(N18130,N18134,N18135);
and and10802(N18143,N18147,N18148);
and and10810(N18156,R6,R7);
and and10818(N18169,N18173,N18174);
and and10826(N18182,R6,N18187);
and and10834(N18195,R6,N18200);
and and10842(N18208,R6,N18213);
and and10850(N18221,N18225,N18226);
and and10858(N18234,N18239,R7);
and and10866(N18247,N18252,R6);
and and10874(N18260,N18265,R7);
and and10882(N18273,N18278,R7);
and and10890(N18286,R6,N18291);
and and10898(N18299,N18304,R7);
and and10906(N18312,R6,N18317);
and and10914(N18325,R6,N18330);
and and10922(N18338,N18342,N18343);
and and10930(N18351,N18355,N18356);
and and10938(N18364,N18368,N18369);
and and10946(N18377,R6,R7);
and and10954(N18390,N18394,N18395);
and and10962(N18403,N18408,R7);
and and10970(N18416,R6,N18421);
and and10978(N18429,N18433,N18434);
and and10986(N18442,R6,N18447);
and and10994(N18455,N18459,N18460);
and and11002(N18468,N18472,N18473);
and and11010(N18481,N18485,N18486);
and and11018(N18494,R6,R7);
and and11026(N18507,R6,N18512);
and and11034(N18520,N18524,N18525);
and and11042(N18533,N18538,R7);
and and11050(N18546,R6,N18551);
and and11058(N18559,R6,N18564);
and and11066(N18572,R5,R6);
and and11074(N18585,R6,N18590);
and and11082(N18598,N18601,N18602);
and and11090(N18610,N18614,R7);
and and11098(N18622,N18625,N18626);
and and11106(N18634,N18637,N18638);
and and11114(N18646,N18650,R7);
and and11122(N18658,R6,N18662);
and and11130(N18670,N18673,N18674);
and and11138(N18682,N18685,N18686);
and and11146(N18694,N18698,R7);
and and11154(N18706,R6,R7);
and and11162(N18718,R6,N18722);
and and11170(N18730,R6,N18734);
and and11178(N18742,R6,N18746);
and and11186(N18754,N18758,R7);
and and11194(N18766,N18769,N18770);
and and11202(N18778,N18782,R7);
and and11210(N18790,N18793,N18794);
and and11218(N18802,N18805,N18806);
and and11226(N18814,N18817,N18818);
and and11234(N18826,N18829,N18830);
and and11242(N18838,R6,N18842);
and and11250(N18850,R5,R6);
and and11258(N18862,R6,N18866);
and and11266(N18874,R6,N18878);
and and11274(N18886,R6,R7);
and and11282(N18898,R4,N18902);
and and11290(N18910,N18914,R7);
and and11298(N18922,R6,N18926);
and and11306(N18934,N18938,R7);
and and11314(N18946,N18950,R7);
and and11322(N18958,R5,N18962);
and and11330(N18970,N18974,R7);
and and11338(N18982,N18986,R7);
and and11346(N18994,R6,R7);
and and11354(N19006,R5,R6);
and and11362(N19018,N19021,N19022);
and and11370(N19030,R6,R7);
and and11378(N19042,N19045,N19046);
and and11386(N19054,R5,N19058);
and and11394(N19066,R5,R7);
and and11402(N19078,N19082,R7);
and and11410(N19090,N19094,R7);
and and11418(N19102,N19106,R7);
and and11426(N19114,N19117,N19118);
and and11434(N19126,R6,N19130);
and and11442(N19138,R5,N19142);
and and11450(N19150,N19153,N19154);
and and11458(N19162,N19165,R7);
and and11466(N19173,N19176,R7);
and and11474(N19184,R6,R7);
and and11482(N19195,N19198,R7);
and and11490(N19206,R5,N19209);
and and11498(N19217,N19220,R7);
and and11506(N19228,N19231,R7);
and and11514(N19239,N19242,R7);
and and11522(N19250,R6,R7);
and and11530(N19261,R6,R7);
and and11538(N19272,R6,N19275);
and and11546(N19283,R6,N19286);
and and11554(N19294,R6,N19297);
and and11562(N19305,N19307,N19308);
and and11570(N19316,R5,N19319);
and and11578(N19327,R6,R7);
and and11586(N19338,R6,N19341);
and and11594(N19349,R6,R7);
and and11602(N19360,R4,N19363);
and and11610(N19371,R6,R7);
and and11618(N19382,R6,R7);
and and11626(N19393,N19396,R7);
and and11634(N19404,R6,R7);
and and11642(N19415,R5,R7);
and and11650(N19426,N19429,R7);
and and11658(N19437,N19440,R7);
and and11666(N19448,R6,N19451);
and and11674(N19459,R6,N19462);
and and11682(N19470,R6,N19473);
and and11690(N19481,N19484,R7);
and and11698(N19492,N19495,R7);
and and11706(N19503,N19506,R7);
and and11714(N19514,R5,R6);
and and11722(N19525,N19528,R7);
and and11730(N19536,N19539,R7);
and and11738(N19547,N19550,R7);
and and11746(N19558,N19561,R7);
and and11754(N19569,N19571,N19572);
and and11762(N19580,R6,R7);
and and11770(N19590,R6,R7);
and and11778(N19600,R6,N19602);
and and11786(N19610,R5,R7);
and and11794(N19620,R6,R7);
and and11802(N19630,R6,R7);
and and11810(N19640,R6,R7);
and and11818(N19650,R6,R7);
and and11826(N19660,R6,N19662);
and and11834(N19670,R6,R7);
and and11842(N19680,R6,R7);
and and11850(N19690,R4,N19692);
and and11858(N19700,N19701,N19702);
and and11866(N19710,R6,R7);
and and11874(N19720,N19722,R7);
and and11882(N19730,R6,N19732);
and and11890(N19740,N19742,R7);
and and11898(N19750,R6,R7);
and and11906(N19760,R6,R7);
and and11914(N19770,R6,R7);
and and11922(N19779,R6,R7);
and and11930(N19788,R5,R7);
and and11938(N19797,R6,R7);
and and11946(N19806,R6,R7);
and and11954(N19815,R6,N19816);
and and11962(N19824,R6,R7);
and and11970(N19833,R6,R7);
and and11978(N19842,R6,R7);
and and11986(N19851,R6,R7);
and and12336(N20635,N20636,N20637);
and and12346(N20651,N20652,N20653);
and and12355(N20669,N20670,N20671);
and and12364(N20687,N20688,N20689);
and and12373(N20704,N20705,N20706);
and and12382(N20721,N20722,N20723);
and and12391(N20738,N20739,N20740);
and and12400(N20755,N20756,N20757);
and and12409(N20772,N20773,N20774);
and and12418(N20789,N20790,N20791);
and and12427(N20806,N20807,N20808);
and and12436(N20823,N20824,N20825);
and and12445(N20840,N20841,N20842);
and and12454(N20857,N20858,N20859);
and and12463(N20874,N20875,N20876);
and and12472(N20891,N20892,N20893);
and and12481(N20908,N20909,N20910);
and and12490(N20924,N20925,N20926);
and and12499(N20940,N20941,N20942);
and and12508(N20956,N20957,N20958);
and and12517(N20972,N20973,N20974);
and and12526(N20988,N20989,N20990);
and and12535(N21004,N21005,N21006);
and and12544(N21020,N21021,N21022);
and and12553(N21036,N21037,N21038);
and and12562(N21052,N21053,N21054);
and and12571(N21068,N21069,N21070);
and and12580(N21084,N21085,N21086);
and and12589(N21100,N21101,N21102);
and and12598(N21116,N21117,N21118);
and and12607(N21132,N21133,N21134);
and and12616(N21148,N21149,N21150);
and and12625(N21164,N21165,N21166);
and and12634(N21180,N21181,N21182);
and and12643(N21196,N21197,N21198);
and and12652(N21212,N21213,N21214);
and and12661(N21228,N21229,N21230);
and and12670(N21244,N21245,N21246);
and and12679(N21260,N21261,N21262);
and and12688(N21276,N21277,N21278);
and and12697(N21292,N21293,N21294);
and and12706(N21308,N21309,N21310);
and and12715(N21323,N21324,N21325);
and and12724(N21338,N21339,N21340);
and and12733(N21353,N21354,N21355);
and and12742(N21368,N21369,N21370);
and and12751(N21383,N21384,N21385);
and and12760(N21398,N21399,N21400);
and and12769(N21413,N21414,N21415);
and and12778(N21428,N21429,N21430);
and and12787(N21443,N21444,N21445);
and and12796(N21458,N21459,N21460);
and and12805(N21473,N21474,N21475);
and and12814(N21488,N21489,N21490);
and and12823(N21503,N21504,N21505);
and and12832(N21518,N21519,N21520);
and and12841(N21533,N21534,N21535);
and and12850(N21548,N21549,N21550);
and and12859(N21563,N21564,N21565);
and and12868(N21578,N21579,N21580);
and and12877(N21593,N21594,N21595);
and and12886(N21608,N21609,N21610);
and and12895(N21623,N21624,N21625);
and and12904(N21638,N21639,N21640);
and and12913(N21653,N21654,N21655);
and and12922(N21668,N21669,N21670);
and and12931(N21683,N21684,N21685);
and and12940(N21697,N21698,N21699);
and and12949(N21711,N21712,N21713);
and and12958(N21725,N21726,N21727);
and and12967(N21739,N21740,N21741);
and and12976(N21753,N21754,N21755);
and and12985(N21767,N21768,N21769);
and and12994(N21781,N21782,N21783);
and and13003(N21795,N21796,N21797);
and and13012(N21809,N21810,N21811);
and and13021(N21823,N21824,N21825);
and and13030(N21837,N21838,N21839);
and and13039(N21851,N21852,N21853);
and and13048(N21865,N21866,N21867);
and and13057(N21879,N21880,N21881);
and and13066(N21893,N21894,N21895);
and and13075(N21907,N21908,N21909);
and and13084(N21921,N21922,N21923);
and and13093(N21935,N21936,N21937);
and and13102(N21949,N21950,N21951);
and and13111(N21963,N21964,N21965);
and and13120(N21977,N21978,N21979);
and and13129(N21991,N21992,N21993);
and and13138(N22005,N22006,N22007);
and and13147(N22019,N22020,N22021);
and and13156(N22033,N22034,N22035);
and and13165(N22047,N22048,N22049);
and and13174(N22061,N22062,N22063);
and and13183(N22075,N22076,N22077);
and and13192(N22089,N22090,N22091);
and and13201(N22103,N22104,N22105);
and and13210(N22117,N22118,N22119);
and and13219(N22131,N22132,N22133);
and and13228(N22145,N22146,N22147);
and and13237(N22159,N22160,N22161);
and and13246(N22173,N22174,N22175);
and and13255(N22187,N22188,N22189);
and and13264(N22201,N22202,N22203);
and and13273(N22214,N22215,N22216);
and and13282(N22227,N22228,N22229);
and and13291(N22240,N22241,N22242);
and and13300(N22253,N22254,N22255);
and and13309(N22266,N22267,N22268);
and and13318(N22279,N22280,N22281);
and and13327(N22292,N22293,N22294);
and and13336(N22305,N22306,N22307);
and and13345(N22318,N22319,N22320);
and and13354(N22331,N22332,N22333);
and and13363(N22344,N22345,N22346);
and and13372(N22357,N22358,N22359);
and and13381(N22370,N22371,N22372);
and and13390(N22383,N22384,N22385);
and and13399(N22396,N22397,N22398);
and and13408(N22409,N22410,N22411);
and and13417(N22422,N22423,N22424);
and and13426(N22435,N22436,N22437);
and and13435(N22448,N22449,N22450);
and and13444(N22461,N22462,N22463);
and and13453(N22474,N22475,N22476);
and and13462(N22487,N22488,N22489);
and and13471(N22500,N22501,N22502);
and and13480(N22513,N22514,N22515);
and and13489(N22526,N22527,N22528);
and and13498(N22539,N22540,N22541);
and and13507(N22552,N22553,N22554);
and and13516(N22565,N22566,N22567);
and and13525(N22578,N22579,N22580);
and and13534(N22591,N22592,N22593);
and and13543(N22604,N22605,N22606);
and and13552(N22617,N22618,N22619);
and and13561(N22630,N22631,N22632);
and and13570(N22643,N22644,N22645);
and and13579(N22656,N22657,N22658);
and and13588(N22669,N22670,N22671);
and and13597(N22682,N22683,N22684);
and and13606(N22694,N22695,N22696);
and and13615(N22706,N22707,N22708);
and and13624(N22718,N22719,N22720);
and and13633(N22730,N22731,N22732);
and and13642(N22742,N22743,N22744);
and and13651(N22754,N22755,N22756);
and and13660(N22766,N22767,N22768);
and and13669(N22778,N22779,N22780);
and and13678(N22790,N22791,N22792);
and and13687(N22802,N22803,N22804);
and and13696(N22814,N22815,N22816);
and and13705(N22826,N22827,N22828);
and and13714(N22838,N22839,N22840);
and and13723(N22850,N22851,N22852);
and and13732(N22862,N22863,N22864);
and and13741(N22874,N22875,N22876);
and and13750(N22886,N22887,N22888);
and and13759(N22898,N22899,N22900);
and and13768(N22910,N22911,N22912);
and and13777(N22922,N22923,N22924);
and and13786(N22933,N22934,N22935);
and and13795(N22944,N22945,N22946);
and and13804(N22955,N22956,N22957);
and and13813(N22966,N22967,N22968);
and and13822(N22977,N22978,N22979);
and and13831(N22988,N22989,N22990);
and and13840(N22999,N23000,N23001);
and and13849(N23010,N23011,N23012);
and and13858(N23020,N23021,N23022);
and and13867(N23030,N23031,N23032);
and and13875(N23046,N23047,N23048);
and and13883(N23062,N23063,N23064);
and and13891(N23078,N23079,N23080);
and and13899(N23093,N23094,N23095);
and and13907(N23108,N23109,N23110);
and and13915(N23123,N23124,N23125);
and and13923(N23137,N23138,N23139);
and and13931(N23151,N23152,N23153);
and and13939(N23165,N23166,N23167);
and and13947(N23179,N23180,N23181);
and and13955(N23193,N23194,N23195);
and and13963(N23207,N23208,N23209);
and and13971(N23221,N23222,N23223);
and and13979(N23235,N23236,N23237);
and and13987(N23248,N23249,N23250);
and and13995(N23261,N23262,N23263);
and and14003(N23274,N23275,N23276);
and and14011(N23287,N23288,N23289);
and and14019(N23300,N23301,N23302);
and and14027(N23313,N23314,N23315);
and and14035(N23326,N23327,N23328);
and and14043(N23339,N23340,N23341);
and and14051(N23352,N23353,N23354);
and and14059(N23365,N23366,N23367);
and and14067(N23378,N23379,N23380);
and and14075(N23391,N23392,N23393);
and and14083(N23404,N23405,N23406);
and and14091(N23417,N23418,N23419);
and and14099(N23430,N23431,N23432);
and and14107(N23443,N23444,N23445);
and and14115(N23455,N23456,N23457);
and and14123(N23467,N23468,N23469);
and and14131(N23479,N23480,N23481);
and and14139(N23491,N23492,N23493);
and and14147(N23503,N23504,N23505);
and and14155(N23515,N23516,N23517);
and and14163(N23527,N23528,N23529);
and and14171(N23539,N23540,N23541);
and and14179(N23551,N23552,N23553);
and and14187(N23563,N23564,N23565);
and and14195(N23575,N23576,N23577);
and and14203(N23587,N23588,N23589);
and and14211(N23599,N23600,N23601);
and and14219(N23611,N23612,N23613);
and and14227(N23622,N23623,N23624);
and and14235(N23633,N23634,N23635);
and and14243(N23644,N23645,N23646);
and and14251(N23655,N23656,N23657);
and and14259(N23666,N23667,N23668);
and and14267(N23677,N23678,N23679);
and and14275(N23688,N23689,N23690);
and and14283(N23699,N23700,N23701);
and and14291(N23710,N23711,N23712);
and and14299(N23721,N23722,N23723);
and and14307(N23731,N23732,N23733);
and and14315(N23740,N23741,N23742);
and and14322(N23753,N23754,N23755);
and and14329(N23765,N23766,N23767);
and and14336(N23776,N23777,N23778);
and and14343(N23787,N23788,N23789);
and and14350(N23797,N23798,N23799);
and and14357(N23807,N23808,N23809);
and and14364(N23815,N23816,N23817);
and and12337(N20636,N20638,N20639);
and and12338(N20637,N20640,N20641);
and and12347(N20652,N20654,N20655);
and and12348(N20653,N20656,N20657);
and and12356(N20670,N20672,N20673);
and and12357(N20671,N20674,N20675);
and and12365(N20688,N20690,N20691);
and and12366(N20689,N20692,N20693);
and and12374(N20705,N20707,N20708);
and and12375(N20706,N20709,N20710);
and and12383(N20722,N20724,N20725);
and and12384(N20723,N20726,N20727);
and and12392(N20739,N20741,N20742);
and and12393(N20740,N20743,N20744);
and and12401(N20756,N20758,N20759);
and and12402(N20757,N20760,N20761);
and and12410(N20773,N20775,N20776);
and and12411(N20774,N20777,N20778);
and and12419(N20790,N20792,N20793);
and and12420(N20791,N20794,N20795);
and and12428(N20807,N20809,N20810);
and and12429(N20808,N20811,N20812);
and and12437(N20824,N20826,N20827);
and and12438(N20825,N20828,N20829);
and and12446(N20841,N20843,N20844);
and and12447(N20842,N20845,N20846);
and and12455(N20858,N20860,N20861);
and and12456(N20859,N20862,N20863);
and and12464(N20875,N20877,N20878);
and and12465(N20876,N20879,N20880);
and and12473(N20892,N20894,N20895);
and and12474(N20893,N20896,N20897);
and and12482(N20909,N20911,N20912);
and and12483(N20910,N20913,N20914);
and and12491(N20925,N20927,N20928);
and and12492(N20926,N20929,N20930);
and and12500(N20941,N20943,N20944);
and and12501(N20942,N20945,N20946);
and and12509(N20957,N20959,N20960);
and and12510(N20958,N20961,N20962);
and and12518(N20973,N20975,N20976);
and and12519(N20974,N20977,N20978);
and and12527(N20989,N20991,N20992);
and and12528(N20990,N20993,N20994);
and and12536(N21005,N21007,N21008);
and and12537(N21006,N21009,N21010);
and and12545(N21021,N21023,N21024);
and and12546(N21022,N21025,N21026);
and and12554(N21037,N21039,N21040);
and and12555(N21038,N21041,N21042);
and and12563(N21053,N21055,N21056);
and and12564(N21054,N21057,N21058);
and and12572(N21069,N21071,N21072);
and and12573(N21070,N21073,N21074);
and and12581(N21085,N21087,N21088);
and and12582(N21086,N21089,N21090);
and and12590(N21101,N21103,N21104);
and and12591(N21102,N21105,N21106);
and and12599(N21117,N21119,N21120);
and and12600(N21118,N21121,N21122);
and and12608(N21133,N21135,N21136);
and and12609(N21134,N21137,N21138);
and and12617(N21149,N21151,N21152);
and and12618(N21150,N21153,N21154);
and and12626(N21165,N21167,N21168);
and and12627(N21166,N21169,N21170);
and and12635(N21181,N21183,N21184);
and and12636(N21182,N21185,N21186);
and and12644(N21197,N21199,N21200);
and and12645(N21198,N21201,N21202);
and and12653(N21213,N21215,N21216);
and and12654(N21214,N21217,N21218);
and and12662(N21229,N21231,N21232);
and and12663(N21230,N21233,N21234);
and and12671(N21245,N21247,N21248);
and and12672(N21246,N21249,N21250);
and and12680(N21261,N21263,N21264);
and and12681(N21262,N21265,N21266);
and and12689(N21277,N21279,N21280);
and and12690(N21278,N21281,N21282);
and and12698(N21293,N21295,N21296);
and and12699(N21294,N21297,N21298);
and and12707(N21309,N21311,N21312);
and and12708(N21310,N21313,N21314);
and and12716(N21324,N21326,N21327);
and and12717(N21325,N21328,N21329);
and and12725(N21339,N21341,N21342);
and and12726(N21340,N21343,N21344);
and and12734(N21354,N21356,N21357);
and and12735(N21355,N21358,N21359);
and and12743(N21369,N21371,N21372);
and and12744(N21370,N21373,N21374);
and and12752(N21384,N21386,N21387);
and and12753(N21385,N21388,N21389);
and and12761(N21399,N21401,N21402);
and and12762(N21400,N21403,N21404);
and and12770(N21414,N21416,N21417);
and and12771(N21415,N21418,N21419);
and and12779(N21429,N21431,N21432);
and and12780(N21430,N21433,N21434);
and and12788(N21444,N21446,N21447);
and and12789(N21445,N21448,N21449);
and and12797(N21459,N21461,N21462);
and and12798(N21460,N21463,N21464);
and and12806(N21474,N21476,N21477);
and and12807(N21475,N21478,N21479);
and and12815(N21489,N21491,N21492);
and and12816(N21490,N21493,N21494);
and and12824(N21504,N21506,N21507);
and and12825(N21505,N21508,N21509);
and and12833(N21519,N21521,N21522);
and and12834(N21520,N21523,N21524);
and and12842(N21534,N21536,N21537);
and and12843(N21535,N21538,N21539);
and and12851(N21549,N21551,N21552);
and and12852(N21550,N21553,N21554);
and and12860(N21564,N21566,N21567);
and and12861(N21565,N21568,N21569);
and and12869(N21579,N21581,N21582);
and and12870(N21580,N21583,N21584);
and and12878(N21594,N21596,N21597);
and and12879(N21595,N21598,N21599);
and and12887(N21609,N21611,N21612);
and and12888(N21610,N21613,N21614);
and and12896(N21624,N21626,N21627);
and and12897(N21625,N21628,N21629);
and and12905(N21639,N21641,N21642);
and and12906(N21640,N21643,N21644);
and and12914(N21654,N21656,N21657);
and and12915(N21655,N21658,N21659);
and and12923(N21669,N21671,N21672);
and and12924(N21670,N21673,N21674);
and and12932(N21684,N21686,N21687);
and and12933(N21685,N21688,N21689);
and and12941(N21698,N21700,N21701);
and and12942(N21699,N21702,N21703);
and and12950(N21712,N21714,N21715);
and and12951(N21713,N21716,N21717);
and and12959(N21726,N21728,N21729);
and and12960(N21727,N21730,N21731);
and and12968(N21740,N21742,N21743);
and and12969(N21741,N21744,N21745);
and and12977(N21754,N21756,N21757);
and and12978(N21755,N21758,N21759);
and and12986(N21768,N21770,N21771);
and and12987(N21769,N21772,N21773);
and and12995(N21782,N21784,N21785);
and and12996(N21783,N21786,N21787);
and and13004(N21796,N21798,N21799);
and and13005(N21797,N21800,N21801);
and and13013(N21810,N21812,N21813);
and and13014(N21811,N21814,N21815);
and and13022(N21824,N21826,N21827);
and and13023(N21825,N21828,N21829);
and and13031(N21838,N21840,N21841);
and and13032(N21839,N21842,N21843);
and and13040(N21852,N21854,N21855);
and and13041(N21853,N21856,N21857);
and and13049(N21866,N21868,N21869);
and and13050(N21867,N21870,N21871);
and and13058(N21880,N21882,N21883);
and and13059(N21881,N21884,N21885);
and and13067(N21894,N21896,N21897);
and and13068(N21895,N21898,N21899);
and and13076(N21908,N21910,N21911);
and and13077(N21909,N21912,N21913);
and and13085(N21922,N21924,N21925);
and and13086(N21923,N21926,N21927);
and and13094(N21936,N21938,N21939);
and and13095(N21937,N21940,N21941);
and and13103(N21950,N21952,N21953);
and and13104(N21951,N21954,N21955);
and and13112(N21964,N21966,N21967);
and and13113(N21965,N21968,N21969);
and and13121(N21978,N21980,N21981);
and and13122(N21979,N21982,N21983);
and and13130(N21992,N21994,N21995);
and and13131(N21993,N21996,N21997);
and and13139(N22006,N22008,N22009);
and and13140(N22007,N22010,N22011);
and and13148(N22020,N22022,N22023);
and and13149(N22021,N22024,N22025);
and and13157(N22034,N22036,N22037);
and and13158(N22035,N22038,N22039);
and and13166(N22048,N22050,N22051);
and and13167(N22049,N22052,N22053);
and and13175(N22062,N22064,N22065);
and and13176(N22063,N22066,N22067);
and and13184(N22076,N22078,N22079);
and and13185(N22077,N22080,N22081);
and and13193(N22090,N22092,N22093);
and and13194(N22091,N22094,N22095);
and and13202(N22104,N22106,N22107);
and and13203(N22105,N22108,N22109);
and and13211(N22118,N22120,N22121);
and and13212(N22119,N22122,N22123);
and and13220(N22132,N22134,N22135);
and and13221(N22133,N22136,N22137);
and and13229(N22146,N22148,N22149);
and and13230(N22147,N22150,N22151);
and and13238(N22160,N22162,N22163);
and and13239(N22161,N22164,N22165);
and and13247(N22174,N22176,N22177);
and and13248(N22175,N22178,N22179);
and and13256(N22188,N22190,N22191);
and and13257(N22189,N22192,N22193);
and and13265(N22202,N22204,N22205);
and and13266(N22203,N22206,N22207);
and and13274(N22215,N22217,N22218);
and and13275(N22216,N22219,N22220);
and and13283(N22228,N22230,N22231);
and and13284(N22229,N22232,N22233);
and and13292(N22241,N22243,N22244);
and and13293(N22242,N22245,N22246);
and and13301(N22254,N22256,N22257);
and and13302(N22255,N22258,N22259);
and and13310(N22267,N22269,N22270);
and and13311(N22268,N22271,N22272);
and and13319(N22280,N22282,N22283);
and and13320(N22281,N22284,N22285);
and and13328(N22293,N22295,N22296);
and and13329(N22294,N22297,N22298);
and and13337(N22306,N22308,N22309);
and and13338(N22307,N22310,N22311);
and and13346(N22319,N22321,N22322);
and and13347(N22320,N22323,N22324);
and and13355(N22332,N22334,N22335);
and and13356(N22333,N22336,N22337);
and and13364(N22345,N22347,N22348);
and and13365(N22346,N22349,N22350);
and and13373(N22358,N22360,N22361);
and and13374(N22359,N22362,N22363);
and and13382(N22371,N22373,N22374);
and and13383(N22372,N22375,N22376);
and and13391(N22384,N22386,N22387);
and and13392(N22385,N22388,N22389);
and and13400(N22397,N22399,N22400);
and and13401(N22398,N22401,N22402);
and and13409(N22410,N22412,N22413);
and and13410(N22411,N22414,N22415);
and and13418(N22423,N22425,N22426);
and and13419(N22424,N22427,N22428);
and and13427(N22436,N22438,N22439);
and and13428(N22437,N22440,N22441);
and and13436(N22449,N22451,N22452);
and and13437(N22450,N22453,N22454);
and and13445(N22462,N22464,N22465);
and and13446(N22463,N22466,N22467);
and and13454(N22475,N22477,N22478);
and and13455(N22476,N22479,N22480);
and and13463(N22488,N22490,N22491);
and and13464(N22489,N22492,N22493);
and and13472(N22501,N22503,N22504);
and and13473(N22502,N22505,N22506);
and and13481(N22514,N22516,N22517);
and and13482(N22515,N22518,N22519);
and and13490(N22527,N22529,N22530);
and and13491(N22528,N22531,N22532);
and and13499(N22540,N22542,N22543);
and and13500(N22541,N22544,N22545);
and and13508(N22553,N22555,N22556);
and and13509(N22554,N22557,N22558);
and and13517(N22566,N22568,N22569);
and and13518(N22567,N22570,N22571);
and and13526(N22579,N22581,N22582);
and and13527(N22580,N22583,N22584);
and and13535(N22592,N22594,N22595);
and and13536(N22593,N22596,N22597);
and and13544(N22605,N22607,N22608);
and and13545(N22606,N22609,N22610);
and and13553(N22618,N22620,N22621);
and and13554(N22619,N22622,N22623);
and and13562(N22631,N22633,N22634);
and and13563(N22632,N22635,N22636);
and and13571(N22644,N22646,N22647);
and and13572(N22645,N22648,N22649);
and and13580(N22657,N22659,N22660);
and and13581(N22658,N22661,N22662);
and and13589(N22670,N22672,N22673);
and and13590(N22671,N22674,N22675);
and and13598(N22683,N22685,N22686);
and and13599(N22684,N22687,N22688);
and and13607(N22695,N22697,N22698);
and and13608(N22696,N22699,N22700);
and and13616(N22707,N22709,N22710);
and and13617(N22708,N22711,N22712);
and and13625(N22719,N22721,N22722);
and and13626(N22720,N22723,N22724);
and and13634(N22731,N22733,N22734);
and and13635(N22732,N22735,N22736);
and and13643(N22743,N22745,N22746);
and and13644(N22744,N22747,N22748);
and and13652(N22755,N22757,N22758);
and and13653(N22756,N22759,N22760);
and and13661(N22767,N22769,N22770);
and and13662(N22768,N22771,N22772);
and and13670(N22779,N22781,N22782);
and and13671(N22780,N22783,N22784);
and and13679(N22791,N22793,N22794);
and and13680(N22792,N22795,N22796);
and and13688(N22803,N22805,N22806);
and and13689(N22804,N22807,N22808);
and and13697(N22815,N22817,N22818);
and and13698(N22816,N22819,N22820);
and and13706(N22827,N22829,N22830);
and and13707(N22828,N22831,N22832);
and and13715(N22839,N22841,N22842);
and and13716(N22840,N22843,N22844);
and and13724(N22851,N22853,N22854);
and and13725(N22852,N22855,N22856);
and and13733(N22863,N22865,N22866);
and and13734(N22864,N22867,N22868);
and and13742(N22875,N22877,N22878);
and and13743(N22876,N22879,N22880);
and and13751(N22887,N22889,N22890);
and and13752(N22888,N22891,N22892);
and and13760(N22899,N22901,N22902);
and and13761(N22900,N22903,N22904);
and and13769(N22911,N22913,N22914);
and and13770(N22912,N22915,N22916);
and and13778(N22923,N22925,N22926);
and and13779(N22924,N22927,N22928);
and and13787(N22934,N22936,N22937);
and and13788(N22935,N22938,N22939);
and and13796(N22945,N22947,N22948);
and and13797(N22946,N22949,N22950);
and and13805(N22956,N22958,N22959);
and and13806(N22957,N22960,N22961);
and and13814(N22967,N22969,N22970);
and and13815(N22968,N22971,N22972);
and and13823(N22978,N22980,N22981);
and and13824(N22979,N22982,N22983);
and and13832(N22989,N22991,N22992);
and and13833(N22990,N22993,N22994);
and and13841(N23000,N23002,N23003);
and and13842(N23001,N23004,N23005);
and and13850(N23011,N23013,N23014);
and and13851(N23012,N23015,N23016);
and and13859(N23021,N23023,N23024);
and and13860(N23022,N23025,N23026);
and and13868(N23031,N23033,N23034);
and and13869(N23032,N23035,N23036);
and and13876(N23047,N23049,N23050);
and and13877(N23048,N23051,N23052);
and and13884(N23063,N23065,N23066);
and and13885(N23064,N23067,N23068);
and and13892(N23079,N23081,N23082);
and and13893(N23080,N23083,N23084);
and and13900(N23094,N23096,N23097);
and and13901(N23095,N23098,N23099);
and and13908(N23109,N23111,N23112);
and and13909(N23110,N23113,N23114);
and and13916(N23124,N23126,N23127);
and and13917(N23125,N23128,N23129);
and and13924(N23138,N23140,N23141);
and and13925(N23139,N23142,N23143);
and and13932(N23152,N23154,N23155);
and and13933(N23153,N23156,N23157);
and and13940(N23166,N23168,N23169);
and and13941(N23167,N23170,N23171);
and and13948(N23180,N23182,N23183);
and and13949(N23181,N23184,N23185);
and and13956(N23194,N23196,N23197);
and and13957(N23195,N23198,N23199);
and and13964(N23208,N23210,N23211);
and and13965(N23209,N23212,N23213);
and and13972(N23222,N23224,N23225);
and and13973(N23223,N23226,N23227);
and and13980(N23236,N23238,N23239);
and and13981(N23237,N23240,N23241);
and and13988(N23249,N23251,N23252);
and and13989(N23250,N23253,N23254);
and and13996(N23262,N23264,N23265);
and and13997(N23263,N23266,N23267);
and and14004(N23275,N23277,N23278);
and and14005(N23276,N23279,N23280);
and and14012(N23288,N23290,N23291);
and and14013(N23289,N23292,N23293);
and and14020(N23301,N23303,N23304);
and and14021(N23302,N23305,N23306);
and and14028(N23314,N23316,N23317);
and and14029(N23315,N23318,N23319);
and and14036(N23327,N23329,N23330);
and and14037(N23328,N23331,N23332);
and and14044(N23340,N23342,N23343);
and and14045(N23341,N23344,N23345);
and and14052(N23353,N23355,N23356);
and and14053(N23354,N23357,N23358);
and and14060(N23366,N23368,N23369);
and and14061(N23367,N23370,N23371);
and and14068(N23379,N23381,N23382);
and and14069(N23380,N23383,N23384);
and and14076(N23392,N23394,N23395);
and and14077(N23393,N23396,N23397);
and and14084(N23405,N23407,N23408);
and and14085(N23406,N23409,N23410);
and and14092(N23418,N23420,N23421);
and and14093(N23419,N23422,N23423);
and and14100(N23431,N23433,N23434);
and and14101(N23432,N23435,N23436);
and and14108(N23444,N23446,N23447);
and and14109(N23445,N23448,N23449);
and and14116(N23456,N23458,N23459);
and and14117(N23457,N23460,N23461);
and and14124(N23468,N23470,N23471);
and and14125(N23469,N23472,N23473);
and and14132(N23480,N23482,N23483);
and and14133(N23481,N23484,N23485);
and and14140(N23492,N23494,N23495);
and and14141(N23493,N23496,N23497);
and and14148(N23504,N23506,N23507);
and and14149(N23505,N23508,N23509);
and and14156(N23516,N23518,N23519);
and and14157(N23517,N23520,N23521);
and and14164(N23528,N23530,N23531);
and and14165(N23529,N23532,N23533);
and and14172(N23540,N23542,N23543);
and and14173(N23541,N23544,N23545);
and and14180(N23552,N23554,N23555);
and and14181(N23553,N23556,N23557);
and and14188(N23564,N23566,N23567);
and and14189(N23565,N23568,N23569);
and and14196(N23576,N23578,N23579);
and and14197(N23577,N23580,N23581);
and and14204(N23588,N23590,N23591);
and and14205(N23589,N23592,N23593);
and and14212(N23600,N23602,N23603);
and and14213(N23601,N23604,N23605);
and and14220(N23612,N23614,N23615);
and and14221(N23613,N23616,N23617);
and and14228(N23623,N23625,N23626);
and and14229(N23624,N23627,N23628);
and and14236(N23634,N23636,N23637);
and and14237(N23635,N23638,N23639);
and and14244(N23645,N23647,N23648);
and and14245(N23646,N23649,N23650);
and and14252(N23656,N23658,N23659);
and and14253(N23657,N23660,N23661);
and and14260(N23667,N23669,N23670);
and and14261(N23668,N23671,N23672);
and and14268(N23678,N23680,N23681);
and and14269(N23679,N23682,N23683);
and and14276(N23689,N23691,N23692);
and and14277(N23690,N23693,N23694);
and and14284(N23700,N23702,N23703);
and and14285(N23701,N23704,N23705);
and and14292(N23711,N23713,N23714);
and and14293(N23712,N23715,N23716);
and and14300(N23722,N23724,N23725);
and and14301(N23723,N23726,N23727);
and and14308(N23732,N23734,N23735);
and and14309(N23733,N23736,N23737);
and and14316(N23741,N23743,N23744);
and and14317(N23742,N23745,N23746);
and and14323(N23754,N23756,N23757);
and and14324(N23755,N23758,N23759);
and and14330(N23766,N23768,N23769);
and and14331(N23767,N23770,N23771);
and and14337(N23777,N23779,N23780);
and and14338(N23778,N23781,N23782);
and and14344(N23788,N23790,N23791);
and and14345(N23789,N23792,N23793);
and and14351(N23798,N23800,N23801);
and and14352(N23799,N23802,N23803);
and and14358(N23808,N23810,N23811);
and and14359(N23809,N23812,N23813);
and and14365(N23816,N23818,N23819);
and and14366(N23817,N23820,N23821);
and and12339(N20638,N20642,N20643);
and and12340(N20639,N20644,N20645);
and and12341(N20640,N20646,in2);
and and12342(N20641,R0,R1);
and and12349(N20654,N20658,N20659);
and and12350(N20655,N20660,N20661);
and and12351(N20656,N20662,R0);
and and12352(N20657,N20663,N20664);
and and12358(N20672,N20676,N20677);
and and12359(N20673,N20678,N20679);
and and12360(N20674,N20680,N20681);
and and12361(N20675,N20682,N20683);
and and12367(N20690,N20694,N20695);
and and12368(N20691,N20696,in1);
and and12369(N20692,N20697,N20698);
and and12370(N20693,N20699,N20700);
and and12376(N20707,N20711,N20712);
and and12377(N20708,N20713,N20714);
and and12378(N20709,in2,N20715);
and and12379(N20710,N20716,N20717);
and and12385(N20724,N20728,N20729);
and and12386(N20725,N20730,N20731);
and and12387(N20726,N20732,R0);
and and12388(N20727,N20733,R2);
and and12394(N20741,N20745,N20746);
and and12395(N20742,N20747,N20748);
and and12396(N20743,N20749,R0);
and and12397(N20744,N20750,N20751);
and and12403(N20758,N20762,N20763);
and and12404(N20759,N20764,N20765);
and and12405(N20760,N20766,N20767);
and and12406(N20761,N20768,R2);
and and12412(N20775,N20779,N20780);
and and12413(N20776,N20781,N20782);
and and12414(N20777,in2,N20783);
and and12415(N20778,N20784,N20785);
and and12421(N20792,N20796,N20797);
and and12422(N20793,N20798,N20799);
and and12423(N20794,R0,N20800);
and and12424(N20795,N20801,N20802);
and and12430(N20809,N20813,N20814);
and and12431(N20810,N20815,N20816);
and and12432(N20811,N20817,N20818);
and and12433(N20812,N20819,N20820);
and and12439(N20826,N20830,N20831);
and and12440(N20827,N20832,N20833);
and and12441(N20828,N20834,N20835);
and and12442(N20829,N20836,N20837);
and and12448(N20843,N20847,N20848);
and and12449(N20844,N20849,N20850);
and and12450(N20845,N20851,N20852);
and and12451(N20846,N20853,N20854);
and and12457(N20860,N20864,N20865);
and and12458(N20861,N20866,N20867);
and and12459(N20862,N20868,N20869);
and and12460(N20863,N20870,N20871);
and and12466(N20877,N20881,N20882);
and and12467(N20878,N20883,N20884);
and and12468(N20879,N20885,N20886);
and and12469(N20880,N20887,N20888);
and and12475(N20894,N20898,N20899);
and and12476(N20895,N20900,N20901);
and and12477(N20896,in2,N20902);
and and12478(N20897,N20903,N20904);
and and12484(N20911,N20915,N20916);
and and12485(N20912,N20917,N20918);
and and12486(N20913,in2,R0);
and and12487(N20914,R1,N20919);
and and12493(N20927,N20931,N20932);
and and12494(N20928,N20933,in1);
and and12495(N20929,N20934,R0);
and and12496(N20930,R1,N20935);
and and12502(N20943,N20947,N20948);
and and12503(N20944,N20949,in1);
and and12504(N20945,N20950,R0);
and and12505(N20946,N20951,N20952);
and and12511(N20959,N20963,N20964);
and and12512(N20960,N20965,N20966);
and and12513(N20961,in2,R0);
and and12514(N20962,N20967,N20968);
and and12520(N20975,N20979,N20980);
and and12521(N20976,N20981,in2);
and and12522(N20977,R0,N20982);
and and12523(N20978,N20983,N20984);
and and12529(N20991,N20995,N20996);
and and12530(N20992,N20997,N20998);
and and12531(N20993,N20999,R1);
and and12532(N20994,R2,R3);
and and12538(N21007,N21011,N21012);
and and12539(N21008,N21013,N21014);
and and12540(N21009,N21015,N21016);
and and12541(N21010,R2,N21017);
and and12547(N21023,N21027,N21028);
and and12548(N21024,N21029,in1);
and and12549(N21025,N21030,N21031);
and and12550(N21026,N21032,R2);
and and12556(N21039,N21043,N21044);
and and12557(N21040,N21045,N21046);
and and12558(N21041,N21047,R1);
and and12559(N21042,N21048,N21049);
and and12565(N21055,N21059,N21060);
and and12566(N21056,N21061,N21062);
and and12567(N21057,N21063,R0);
and and12568(N21058,N21064,N21065);
and and12574(N21071,N21075,N21076);
and and12575(N21072,N21077,N21078);
and and12576(N21073,in2,N21079);
and and12577(N21074,N21080,N21081);
and and12583(N21087,N21091,N21092);
and and12584(N21088,N21093,N21094);
and and12585(N21089,N21095,R0);
and and12586(N21090,N21096,N21097);
and and12592(N21103,N21107,N21108);
and and12593(N21104,N21109,N21110);
and and12594(N21105,in2,N21111);
and and12595(N21106,N21112,N21113);
and and12601(N21119,N21123,N21124);
and and12602(N21120,N21125,N21126);
and and12603(N21121,N21127,N21128);
and and12604(N21122,R2,R3);
and and12610(N21135,N21139,N21140);
and and12611(N21136,N21141,N21142);
and and12612(N21137,N21143,R0);
and and12613(N21138,N21144,N21145);
and and12619(N21151,N21155,N21156);
and and12620(N21152,N21157,N21158);
and and12621(N21153,N21159,N21160);
and and12622(N21154,N21161,R3);
and and12628(N21167,N21171,N21172);
and and12629(N21168,N21173,N21174);
and and12630(N21169,in2,N21175);
and and12631(N21170,R1,N21176);
and and12637(N21183,N21187,N21188);
and and12638(N21184,N21189,N21190);
and and12639(N21185,N21191,R0);
and and12640(N21186,N21192,N21193);
and and12646(N21199,N21203,N21204);
and and12647(N21200,N21205,N21206);
and and12648(N21201,N21207,R0);
and and12649(N21202,R1,N21208);
and and12655(N21215,N21219,N21220);
and and12656(N21216,N21221,N21222);
and and12657(N21217,N21223,R0);
and and12658(N21218,R1,N21224);
and and12664(N21231,N21235,N21236);
and and12665(N21232,N21237,N21238);
and and12666(N21233,N21239,N21240);
and and12667(N21234,R1,R3);
and and12673(N21247,N21251,N21252);
and and12674(N21248,N21253,N21254);
and and12675(N21249,in2,N21255);
and and12676(N21250,N21256,R3);
and and12682(N21263,N21267,N21268);
and and12683(N21264,N21269,N21270);
and and12684(N21265,R0,N21271);
and and12685(N21266,N21272,N21273);
and and12691(N21279,N21283,N21284);
and and12692(N21280,N21285,N21286);
and and12693(N21281,N21287,N21288);
and and12694(N21282,N21289,R3);
and and12700(N21295,N21299,N21300);
and and12701(N21296,N21301,in1);
and and12702(N21297,N21302,N21303);
and and12703(N21298,R1,N21304);
and and12709(N21311,N21315,N21316);
and and12710(N21312,N21317,N21318);
and and12711(N21313,N21319,N21320);
and and12712(N21314,R2,R3);
and and12718(N21326,N21330,N21331);
and and12719(N21327,N21332,in1);
and and12720(N21328,in2,N21333);
and and12721(N21329,R1,R2);
and and12727(N21341,N21345,N21346);
and and12728(N21342,N21347,N21348);
and and12729(N21343,N21349,R0);
and and12730(N21344,N21350,R2);
and and12736(N21356,N21360,N21361);
and and12737(N21357,N21362,N21363);
and and12738(N21358,N21364,N21365);
and and12739(N21359,N21366,R3);
and and12745(N21371,N21375,N21376);
and and12746(N21372,N21377,N21378);
and and12747(N21373,N21379,R0);
and and12748(N21374,N21380,R2);
and and12754(N21386,N21390,N21391);
and and12755(N21387,N21392,in1);
and and12756(N21388,N21393,R0);
and and12757(N21389,R2,N21394);
and and12763(N21401,N21405,N21406);
and and12764(N21402,N21407,N21408);
and and12765(N21403,in2,N21409);
and and12766(N21404,R1,R3);
and and12772(N21416,N21420,N21421);
and and12773(N21417,N21422,N21423);
and and12774(N21418,N21424,N21425);
and and12775(N21419,R1,R3);
and and12781(N21431,N21435,N21436);
and and12782(N21432,N21437,in1);
and and12783(N21433,N21438,R0);
and and12784(N21434,N21439,N21440);
and and12790(N21446,N21450,N21451);
and and12791(N21447,N21452,N21453);
and and12792(N21448,N21454,R0);
and and12793(N21449,R1,N21455);
and and12799(N21461,N21465,N21466);
and and12800(N21462,N21467,N21468);
and and12801(N21463,in2,R1);
and and12802(N21464,R2,N21469);
and and12808(N21476,N21480,N21481);
and and12809(N21477,N21482,N21483);
and and12810(N21478,in2,N21484);
and and12811(N21479,N21485,R2);
and and12817(N21491,N21495,N21496);
and and12818(N21492,N21497,N21498);
and and12819(N21493,N21499,R1);
and and12820(N21494,R2,R3);
and and12826(N21506,N21510,N21511);
and and12827(N21507,in0,N21512);
and and12828(N21508,R0,N21513);
and and12829(N21509,R2,N21514);
and and12835(N21521,N21525,N21526);
and and12836(N21522,in1,N21527);
and and12837(N21523,R0,N21528);
and and12838(N21524,R2,N21529);
and and12844(N21536,N21540,N21541);
and and12845(N21537,N21542,N21543);
and and12846(N21538,N21544,R0);
and and12847(N21539,N21545,N21546);
and and12853(N21551,N21555,N21556);
and and12854(N21552,N21557,in1);
and and12855(N21553,N21558,N21559);
and and12856(N21554,R1,R3);
and and12862(N21566,N21570,N21571);
and and12863(N21567,N21572,N21573);
and and12864(N21568,N21574,R0);
and and12865(N21569,R1,N21575);
and and12871(N21581,N21585,N21586);
and and12872(N21582,N21587,in1);
and and12873(N21583,in2,N21588);
and and12874(N21584,N21589,R2);
and and12880(N21596,N21600,N21601);
and and12881(N21597,N21602,in1);
and and12882(N21598,N21603,R0);
and and12883(N21599,R1,R3);
and and12889(N21611,N21615,N21616);
and and12890(N21612,N21617,in1);
and and12891(N21613,in2,N21618);
and and12892(N21614,N21619,N21620);
and and12898(N21626,N21630,N21631);
and and12899(N21627,N21632,N21633);
and and12900(N21628,N21634,N21635);
and and12901(N21629,R2,R3);
and and12907(N21641,N21645,N21646);
and and12908(N21642,N21647,N21648);
and and12909(N21643,R0,N21649);
and and12910(N21644,N21650,N21651);
and and12916(N21656,N21660,N21661);
and and12917(N21657,N21662,in2);
and and12918(N21658,R0,N21663);
and and12919(N21659,N21664,N21665);
and and12925(N21671,N21675,N21676);
and and12926(N21672,N21677,in1);
and and12927(N21673,N21678,N21679);
and and12928(N21674,N21680,R2);
and and12934(N21686,N21690,N21691);
and and12935(N21687,N21692,in1);
and and12936(N21688,in2,R0);
and and12937(N21689,N21693,R2);
and and12943(N21700,N21704,N21705);
and and12944(N21701,N21706,N21707);
and and12945(N21702,in2,R0);
and and12946(N21703,N21708,N21709);
and and12952(N21714,N21718,N21719);
and and12953(N21715,N21720,in1);
and and12954(N21716,N21721,N21722);
and and12955(N21717,R2,N21723);
and and12961(N21728,N21732,N21733);
and and12962(N21729,N21734,in2);
and and12963(N21730,N21735,R1);
and and12964(N21731,R2,N21736);
and and12970(N21742,N21746,N21747);
and and12971(N21743,in0,in2);
and and12972(N21744,N21748,R1);
and and12973(N21745,R2,R3);
and and12979(N21756,N21760,N21761);
and and12980(N21757,in0,in1);
and and12981(N21758,N21762,N21763);
and and12982(N21759,R1,R2);
and and12988(N21770,N21774,N21775);
and and12989(N21771,N21776,in1);
and and12990(N21772,N21777,N21778);
and and12991(N21773,R1,R2);
and and12997(N21784,N21788,N21789);
and and12998(N21785,N21790,in2);
and and12999(N21786,R0,N21791);
and and13000(N21787,N21792,R3);
and and13006(N21798,N21802,N21803);
and and13007(N21799,N21804,in1);
and and13008(N21800,N21805,R0);
and and13009(N21801,N21806,R3);
and and13015(N21812,N21816,N21817);
and and13016(N21813,N21818,N21819);
and and13017(N21814,in2,N21820);
and and13018(N21815,R1,R3);
and and13024(N21826,N21830,N21831);
and and13025(N21827,N21832,in1);
and and13026(N21828,in2,N21833);
and and13027(N21829,R2,N21834);
and and13033(N21840,N21844,N21845);
and and13034(N21841,N21846,in1);
and and13035(N21842,N21847,N21848);
and and13036(N21843,R1,R2);
and and13042(N21854,N21858,N21859);
and and13043(N21855,N21860,N21861);
and and13044(N21856,N21862,R0);
and and13045(N21857,R1,R3);
and and13051(N21868,N21872,N21873);
and and13052(N21869,N21874,in1);
and and13053(N21870,in2,N21875);
and and13054(N21871,R2,R3);
and and13060(N21882,N21886,N21887);
and and13061(N21883,N21888,in1);
and and13062(N21884,in2,R1);
and and13063(N21885,N21889,N21890);
and and13069(N21896,N21900,N21901);
and and13070(N21897,N21902,N21903);
and and13071(N21898,in2,R0);
and and13072(N21899,N21904,R3);
and and13078(N21910,N21914,N21915);
and and13079(N21911,N21916,N21917);
and and13080(N21912,N21918,N21919);
and and13081(N21913,R1,R2);
and and13087(N21924,N21928,N21929);
and and13088(N21925,N21930,in1);
and and13089(N21926,in2,N21931);
and and13090(N21927,R2,N21932);
and and13096(N21938,N21942,N21943);
and and13097(N21939,N21944,N21945);
and and13098(N21940,N21946,R0);
and and13099(N21941,R1,R2);
and and13105(N21952,N21956,N21957);
and and13106(N21953,N21958,N21959);
and and13107(N21954,R0,R1);
and and13108(N21955,R2,N21960);
and and13114(N21966,N21970,N21971);
and and13115(N21967,N21972,in1);
and and13116(N21968,in2,R0);
and and13117(N21969,N21973,N21974);
and and13123(N21980,N21984,N21985);
and and13124(N21981,N21986,N21987);
and and13125(N21982,in2,R0);
and and13126(N21983,N21988,R2);
and and13132(N21994,N21998,N21999);
and and13133(N21995,N22000,in2);
and and13134(N21996,R0,R1);
and and13135(N21997,R2,N22001);
and and13141(N22008,N22012,N22013);
and and13142(N22009,N22014,in1);
and and13143(N22010,in2,R0);
and and13144(N22011,N22015,N22016);
and and13150(N22022,N22026,N22027);
and and13151(N22023,N22028,N22029);
and and13152(N22024,in2,R0);
and and13153(N22025,R1,R2);
and and13159(N22036,N22040,N22041);
and and13160(N22037,N22042,N22043);
and and13161(N22038,in2,R0);
and and13162(N22039,R1,N22044);
and and13168(N22050,N22054,N22055);
and and13169(N22051,N22056,in1);
and and13170(N22052,in2,R1);
and and13171(N22053,N22057,R3);
and and13177(N22064,N22068,N22069);
and and13178(N22065,N22070,in1);
and and13179(N22066,N22071,N22072);
and and13180(N22067,R2,R3);
and and13186(N22078,N22082,N22083);
and and13187(N22079,N22084,in1);
and and13188(N22080,in2,R0);
and and13189(N22081,N22085,N22086);
and and13195(N22092,N22096,N22097);
and and13196(N22093,N22098,in1);
and and13197(N22094,in2,R0);
and and13198(N22095,R1,N22099);
and and13204(N22106,N22110,N22111);
and and13205(N22107,N22112,N22113);
and and13206(N22108,in2,N22114);
and and13207(N22109,R2,R3);
and and13213(N22120,N22124,N22125);
and and13214(N22121,N22126,N22127);
and and13215(N22122,in2,N22128);
and and13216(N22123,R1,R2);
and and13222(N22134,N22138,N22139);
and and13223(N22135,N22140,N22141);
and and13224(N22136,in2,N22142);
and and13225(N22137,N22143,R2);
and and13231(N22148,N22152,N22153);
and and13232(N22149,N22154,N22155);
and and13233(N22150,in2,R0);
and and13234(N22151,N22156,N22157);
and and13240(N22162,N22166,N22167);
and and13241(N22163,N22168,in1);
and and13242(N22164,in2,R0);
and and13243(N22165,N22169,N22170);
and and13249(N22176,N22180,N22181);
and and13250(N22177,N22182,N22183);
and and13251(N22178,in2,R1);
and and13252(N22179,N22184,R3);
and and13258(N22190,N22194,N22195);
and and13259(N22191,N22196,N22197);
and and13260(N22192,in2,N22198);
and and13261(N22193,N22199,R2);
and and13267(N22204,N22208,N22209);
and and13268(N22205,N22210,N22211);
and and13269(N22206,N22212,R1);
and and13270(N22207,R2,R3);
and and13276(N22217,N22221,N22222);
and and13277(N22218,N22223,N22224);
and and13278(N22219,N22225,R1);
and and13279(N22220,N22226,R3);
and and13285(N22230,N22234,N22235);
and and13286(N22231,N22236,N22237);
and and13287(N22232,R0,N22238);
and and13288(N22233,R2,R3);
and and13294(N22243,N22247,N22248);
and and13295(N22244,N22249,in1);
and and13296(N22245,R0,R1);
and and13297(N22246,R2,N22250);
and and13303(N22256,N22260,N22261);
and and13304(N22257,N22262,in1);
and and13305(N22258,in2,N22263);
and and13306(N22259,R1,R2);
and and13312(N22269,N22273,N22274);
and and13313(N22270,in1,N22275);
and and13314(N22271,R0,R1);
and and13315(N22272,N22276,R3);
and and13321(N22282,N22286,N22287);
and and13322(N22283,N22288,in1);
and and13323(N22284,R0,N22289);
and and13324(N22285,R2,R3);
and and13330(N22295,N22299,N22300);
and and13331(N22296,N22301,in1);
and and13332(N22297,R0,R1);
and and13333(N22298,R2,R3);
and and13339(N22308,N22312,N22313);
and and13340(N22309,N22314,in1);
and and13341(N22310,N22315,R0);
and and13342(N22311,R1,N22316);
and and13348(N22321,N22325,N22326);
and and13349(N22322,N22327,in1);
and and13350(N22323,N22328,N22329);
and and13351(N22324,N22330,R3);
and and13357(N22334,N22338,N22339);
and and13358(N22335,N22340,N22341);
and and13359(N22336,R0,R1);
and and13360(N22337,N22342,R3);
and and13366(N22347,N22351,N22352);
and and13367(N22348,N22353,N22354);
and and13368(N22349,in2,R1);
and and13369(N22350,R2,N22355);
and and13375(N22360,N22364,N22365);
and and13376(N22361,N22366,in1);
and and13377(N22362,N22367,N22368);
and and13378(N22363,R1,R3);
and and13384(N22373,N22377,N22378);
and and13385(N22374,in1,N22379);
and and13386(N22375,R0,R1);
and and13387(N22376,R2,R3);
and and13393(N22386,N22390,N22391);
and and13394(N22387,N22392,in1);
and and13395(N22388,N22393,R0);
and and13396(N22389,N22394,N22395);
and and13402(N22399,N22403,N22404);
and and13403(N22400,N22405,in1);
and and13404(N22401,N22406,R1);
and and13405(N22402,N22407,R3);
and and13411(N22412,N22416,N22417);
and and13412(N22413,in0,in1);
and and13413(N22414,in2,R0);
and and13414(N22415,N22418,R2);
and and13420(N22425,N22429,N22430);
and and13421(N22426,N22431,N22432);
and and13422(N22427,in2,R0);
and and13423(N22428,R1,R3);
and and13429(N22438,N22442,N22443);
and and13430(N22439,N22444,in1);
and and13431(N22440,N22445,R0);
and and13432(N22441,R1,N22446);
and and13438(N22451,N22455,N22456);
and and13439(N22452,N22457,N22458);
and and13440(N22453,R0,R1);
and and13441(N22454,R2,N22459);
and and13447(N22464,N22468,N22469);
and and13448(N22465,N22470,N22471);
and and13449(N22466,R0,R1);
and and13450(N22467,R2,N22472);
and and13456(N22477,N22481,N22482);
and and13457(N22478,N22483,in2);
and and13458(N22479,N22484,R1);
and and13459(N22480,R2,N22485);
and and13465(N22490,N22494,N22495);
and and13466(N22491,N22496,in1);
and and13467(N22492,N22497,N22498);
and and13468(N22493,R1,R2);
and and13474(N22503,N22507,N22508);
and and13475(N22504,N22509,in1);
and and13476(N22505,N22510,N22511);
and and13477(N22506,N22512,R2);
and and13483(N22516,N22520,N22521);
and and13484(N22517,N22522,N22523);
and and13485(N22518,in2,R0);
and and13486(N22519,R1,R2);
and and13492(N22529,N22533,N22534);
and and13493(N22530,in0,in2);
and and13494(N22531,R0,N22535);
and and13495(N22532,N22536,R3);
and and13501(N22542,N22546,N22547);
and and13502(N22543,N22548,in1);
and and13503(N22544,in2,R0);
and and13504(N22545,N22549,R3);
and and13510(N22555,N22559,N22560);
and and13511(N22556,in1,in2);
and and13512(N22557,N22561,N22562);
and and13513(N22558,R2,R3);
and and13519(N22568,N22572,N22573);
and and13520(N22569,in0,in1);
and and13521(N22570,N22574,N22575);
and and13522(N22571,N22576,R2);
and and13528(N22581,N22585,N22586);
and and13529(N22582,N22587,in1);
and and13530(N22583,in2,R0);
and and13531(N22584,R1,N22588);
and and13537(N22594,N22598,N22599);
and and13538(N22595,N22600,N22601);
and and13539(N22596,R0,R1);
and and13540(N22597,R2,R3);
and and13546(N22607,N22611,N22612);
and and13547(N22608,N22613,in1);
and and13548(N22609,in2,N22614);
and and13549(N22610,R1,R2);
and and13555(N22620,N22624,N22625);
and and13556(N22621,N22626,N22627);
and and13557(N22622,in2,R1);
and and13558(N22623,R2,R3);
and and13564(N22633,N22637,N22638);
and and13565(N22634,N22639,in1);
and and13566(N22635,in2,R0);
and and13567(N22636,N22640,N22641);
and and13573(N22646,N22650,N22651);
and and13574(N22647,N22652,in1);
and and13575(N22648,N22653,R0);
and and13576(N22649,R1,N22654);
and and13582(N22659,N22663,N22664);
and and13583(N22660,N22665,in1);
and and13584(N22661,in2,R0);
and and13585(N22662,N22666,N22667);
and and13591(N22672,N22676,N22677);
and and13592(N22673,in0,in2);
and and13593(N22674,R0,N22678);
and and13594(N22675,N22679,R3);
and and13600(N22685,N22689,N22690);
and and13601(N22686,N22691,in1);
and and13602(N22687,in2,R0);
and and13603(N22688,R2,R3);
and and13609(N22697,N22701,N22702);
and and13610(N22698,N22703,N22704);
and and13611(N22699,in2,R0);
and and13612(N22700,R1,R2);
and and13618(N22709,N22713,N22714);
and and13619(N22710,N22715,N22716);
and and13620(N22711,in2,N22717);
and and13621(N22712,R1,R2);
and and13627(N22721,N22725,N22726);
and and13628(N22722,N22727,N22728);
and and13629(N22723,in2,R0);
and and13630(N22724,R2,N22729);
and and13636(N22733,N22737,N22738);
and and13637(N22734,N22739,in1);
and and13638(N22735,in2,N22740);
and and13639(N22736,N22741,R2);
and and13645(N22745,N22749,N22750);
and and13646(N22746,in0,N22751);
and and13647(N22747,N22752,R1);
and and13648(N22748,R2,R3);
and and13654(N22757,N22761,N22762);
and and13655(N22758,N22763,in1);
and and13656(N22759,in2,R0);
and and13657(N22760,N22764,R2);
and and13663(N22769,N22773,N22774);
and and13664(N22770,in0,in1);
and and13665(N22771,N22775,N22776);
and and13666(N22772,R1,R2);
and and13672(N22781,N22785,N22786);
and and13673(N22782,N22787,in1);
and and13674(N22783,in2,N22788);
and and13675(N22784,R1,R2);
and and13681(N22793,N22797,N22798);
and and13682(N22794,N22799,in2);
and and13683(N22795,N22800,N22801);
and and13684(N22796,R2,R3);
and and13690(N22805,N22809,N22810);
and and13691(N22806,N22811,N22812);
and and13692(N22807,in2,R0);
and and13693(N22808,R1,N22813);
and and13699(N22817,N22821,N22822);
and and13700(N22818,N22823,in1);
and and13701(N22819,in2,N22824);
and and13702(N22820,R2,N22825);
and and13708(N22829,N22833,N22834);
and and13709(N22830,N22835,N22836);
and and13710(N22831,R0,R1);
and and13711(N22832,R2,R3);
and and13717(N22841,N22845,N22846);
and and13718(N22842,N22847,in1);
and and13719(N22843,in2,N22848);
and and13720(N22844,N22849,R3);
and and13726(N22853,N22857,N22858);
and and13727(N22854,N22859,in1);
and and13728(N22855,in2,R0);
and and13729(N22856,N22860,R3);
and and13735(N22865,N22869,N22870);
and and13736(N22866,in1,in2);
and and13737(N22867,R0,N22871);
and and13738(N22868,R2,N22872);
and and13744(N22877,N22881,N22882);
and and13745(N22878,N22883,in1);
and and13746(N22879,in2,R0);
and and13747(N22880,R1,R2);
and and13753(N22889,N22893,N22894);
and and13754(N22890,N22895,in2);
and and13755(N22891,R0,R1);
and and13756(N22892,R2,R3);
and and13762(N22901,N22905,N22906);
and and13763(N22902,in0,in1);
and and13764(N22903,in2,R0);
and and13765(N22904,R1,N22907);
and and13771(N22913,N22917,N22918);
and and13772(N22914,in0,in1);
and and13773(N22915,in2,R0);
and and13774(N22916,R1,R3);
and and13780(N22925,N22929,N22930);
and and13781(N22926,N22931,in1);
and and13782(N22927,in2,R0);
and and13783(N22928,R1,R2);
and and13789(N22936,N22940,N22941);
and and13790(N22937,N22942,in1);
and and13791(N22938,N22943,R1);
and and13792(N22939,R2,R3);
and and13798(N22947,N22951,N22952);
and and13799(N22948,N22953,in1);
and and13800(N22949,R0,R1);
and and13801(N22950,R2,R3);
and and13807(N22958,N22962,N22963);
and and13808(N22959,N22964,in2);
and and13809(N22960,R0,R1);
and and13810(N22961,R2,R3);
and and13816(N22969,N22973,N22974);
and and13817(N22970,in0,in2);
and and13818(N22971,R0,R1);
and and13819(N22972,R2,R3);
and and13825(N22980,N22984,N22985);
and and13826(N22981,in0,in1);
and and13827(N22982,R0,R1);
and and13828(N22983,R2,R3);
and and13834(N22991,N22995,N22996);
and and13835(N22992,N22997,in1);
and and13836(N22993,N22998,R0);
and and13837(N22994,R2,R3);
and and13843(N23002,N23006,N23007);
and and13844(N23003,in0,in2);
and and13845(N23004,N23008,R1);
and and13846(N23005,R2,R3);
and and13852(N23013,N23017,N23018);
and and13853(N23014,N23019,in1);
and and13854(N23015,in2,R0);
and and13855(N23016,R1,R2);
and and13861(N23023,N23027,N23028);
and and13862(N23024,in1,in2);
and and13863(N23025,R0,R1);
and and13864(N23026,R2,R3);
and and13870(N23033,N23037,N23038);
and and13871(N23034,N23039,N23040);
and and13872(N23035,N23041,N23042);
and and13873(N23036,R4,N23043);
and and13878(N23049,N23053,N23054);
and and13879(N23050,in1,N23055);
and and13880(N23051,N23056,N23057);
and and13881(N23052,N23058,N23059);
and and13886(N23065,N23069,N23070);
and and13887(N23066,N23071,N23072);
and and13888(N23067,N23073,N23074);
and and13889(N23068,N23075,N23076);
and and13894(N23081,N23085,N23086);
and and13895(N23082,N23087,N23088);
and and13896(N23083,R1,N23089);
and and13897(N23084,R3,N23090);
and and13902(N23096,N23100,in0);
and and13903(N23097,N23101,N23102);
and and13904(N23098,R2,N23103);
and and13905(N23099,N23104,N23105);
and and13910(N23111,N23115,N23116);
and and13911(N23112,N23117,N23118);
and and13912(N23113,N23119,R2);
and and13913(N23114,N23120,R4);
and and13918(N23126,N23130,N23131);
and and13919(N23127,in1,in2);
and and13920(N23128,N23132,R1);
and and13921(N23129,N23133,N23134);
and and13926(N23140,N23144,N23145);
and and13927(N23141,N23146,in2);
and and13928(N23142,R0,N23147);
and and13929(N23143,R2,N23148);
and and13934(N23154,N23158,N23159);
and and13935(N23155,in1,N23160);
and and13936(N23156,N23161,R2);
and and13937(N23157,N23162,N23163);
and and13942(N23168,N23172,N23173);
and and13943(N23169,in1,R0);
and and13944(N23170,N23174,N23175);
and and13945(N23171,R3,N23176);
and and13950(N23182,N23186,N23187);
and and13951(N23183,N23188,N23189);
and and13952(N23184,N23190,R2);
and and13953(N23185,R3,R5);
and and13958(N23196,N23200,N23201);
and and13959(N23197,N23202,in2);
and and13960(N23198,N23203,R3);
and and13961(N23199,N23204,N23205);
and and13966(N23210,N23214,N23215);
and and13967(N23211,in1,N23216);
and and13968(N23212,N23217,N23218);
and and13969(N23213,N23219,R3);
and and13974(N23224,N23228,N23229);
and and13975(N23225,in2,N23230);
and and13976(N23226,N23231,R3);
and and13977(N23227,N23232,N23233);
and and13982(N23238,N23242,N23243);
and and13983(N23239,in1,N23244);
and and13984(N23240,N23245,R3);
and and13985(N23241,R4,R5);
and and13990(N23251,N23255,in0);
and and13991(N23252,R0,N23256);
and and13992(N23253,N23257,N23258);
and and13993(N23254,N23259,R5);
and and13998(N23264,N23268,in0);
and and13999(N23265,R0,R1);
and and14000(N23266,R2,N23269);
and and14001(N23267,N23270,N23271);
and and14006(N23277,N23281,in0);
and and14007(N23278,N23282,N23283);
and and14008(N23279,R2,R3);
and and14009(N23280,N23284,N23285);
and and14014(N23290,N23294,in0);
and and14015(N23291,N23295,N23296);
and and14016(N23292,R2,N23297);
and and14017(N23293,R4,R5);
and and14022(N23303,N23307,N23308);
and and14023(N23304,in1,N23309);
and and14024(N23305,N23310,R2);
and and14025(N23306,N23311,N23312);
and and14030(N23316,N23320,N23321);
and and14031(N23317,N23322,N23323);
and and14032(N23318,R0,N23324);
and and14033(N23319,R2,N23325);
and and14038(N23329,N23333,N23334);
and and14039(N23330,N23335,in2);
and and14040(N23331,R0,N23336);
and and14041(N23332,R4,N23337);
and and14046(N23342,N23346,N23347);
and and14047(N23343,N23348,N23349);
and and14048(N23344,R0,R1);
and and14049(N23345,R2,N23350);
and and14054(N23355,N23359,N23360);
and and14055(N23356,N23361,N23362);
and and14056(N23357,N23363,R2);
and and14057(N23358,N23364,R4);
and and14062(N23368,N23372,N23373);
and and14063(N23369,N23374,N23375);
and and14064(N23370,N23376,N23377);
and and14065(N23371,R3,R4);
and and14070(N23381,N23385,N23386);
and and14071(N23382,in1,N23387);
and and14072(N23383,N23388,R2);
and and14073(N23384,N23389,R4);
and and14078(N23394,N23398,N23399);
and and14079(N23395,R0,N23400);
and and14080(N23396,N23401,R3);
and and14081(N23397,N23402,R5);
and and14086(N23407,N23411,N23412);
and and14087(N23408,R0,N23413);
and and14088(N23409,N23414,R3);
and and14089(N23410,N23415,R5);
and and14094(N23420,N23424,N23425);
and and14095(N23421,in2,R0);
and and14096(N23422,N23426,R2);
and and14097(N23423,N23427,N23428);
and and14102(N23433,N23437,N23438);
and and14103(N23434,R0,N23439);
and and14104(N23435,N23440,R3);
and and14105(N23436,N23441,R5);
and and14110(N23446,N23450,in0);
and and14111(N23447,R0,R1);
and and14112(N23448,N23451,R3);
and and14113(N23449,N23452,N23453);
and and14118(N23458,N23462,in0);
and and14119(N23459,R0,R1);
and and14120(N23460,N23463,R3);
and and14121(N23461,R4,N23464);
and and14126(N23470,N23474,in0);
and and14127(N23471,N23475,N23476);
and and14128(N23472,R1,R2);
and and14129(N23473,R3,R4);
and and14134(N23482,N23486,N23487);
and and14135(N23483,in1,R1);
and and14136(N23484,R2,N23488);
and and14137(N23485,R4,N23489);
and and14142(N23494,N23498,N23499);
and and14143(N23495,N23500,R0);
and and14144(N23496,N23501,R2);
and and14145(N23497,R3,R4);
and and14150(N23506,N23510,in0);
and and14151(N23507,N23511,R0);
and and14152(N23508,R1,N23512);
and and14153(N23509,R4,N23513);
and and14158(N23518,N23522,N23523);
and and14159(N23519,in1,N23524);
and and14160(N23520,R0,R1);
and and14161(N23521,R2,N23525);
and and14166(N23530,N23534,in0);
and and14167(N23531,N23535,N23536);
and and14168(N23532,N23537,R3);
and and14169(N23533,R4,R5);
and and14174(N23542,N23546,in0);
and and14175(N23543,R0,R1);
and and14176(N23544,N23547,R3);
and and14177(N23545,N23548,N23549);
and and14182(N23554,N23558,in0);
and and14183(N23555,N23559,R0);
and and14184(N23556,N23560,R2);
and and14185(N23557,N23561,R4);
and and14190(N23566,N23570,in0);
and and14191(N23567,N23571,N23572);
and and14192(N23568,N23573,R2);
and and14193(N23569,R3,N23574);
and and14198(N23578,N23582,in0);
and and14199(N23579,N23583,R0);
and and14200(N23580,R1,R3);
and and14201(N23581,R4,N23584);
and and14206(N23590,N23594,in0);
and and14207(N23591,N23595,R0);
and and14208(N23592,N23596,R2);
and and14209(N23593,N23597,R4);
and and14214(N23602,N23606,in0);
and and14215(N23603,N23607,N23608);
and and14216(N23604,N23609,R2);
and and14217(N23605,R3,N23610);
and and14222(N23614,N23618,in0);
and and14223(N23615,N23619,R1);
and and14224(N23616,N23620,R3);
and and14225(N23617,N23621,R5);
and and14230(N23625,N23629,in0);
and and14231(N23626,R0,R1);
and and14232(N23627,R2,N23630);
and and14233(N23628,R4,N23631);
and and14238(N23636,N23640,N23641);
and and14239(N23637,in1,R0);
and and14240(N23638,R1,R2);
and and14241(N23639,R3,N23642);
and and14246(N23647,N23651,in0);
and and14247(N23648,in1,R0);
and and14248(N23649,R1,N23652);
and and14249(N23650,R4,N23653);
and and14254(N23658,N23662,in0);
and and14255(N23659,R0,R1);
and and14256(N23660,R2,N23663);
and and14257(N23661,R4,N23664);
and and14262(N23669,N23673,in1);
and and14263(N23670,R0,N23674);
and and14264(N23671,R2,N23675);
and and14265(N23672,R4,R5);
and and14270(N23680,N23684,in0);
and and14271(N23681,R0,N23685);
and and14272(N23682,R2,N23686);
and and14273(N23683,R4,R5);
and and14278(N23691,N23695,in0);
and and14279(N23692,in2,N23696);
and and14280(N23693,N23697,R2);
and and14281(N23694,R3,N23698);
and and14286(N23702,N23706,in0);
and and14287(N23703,in2,N23707);
and and14288(N23704,R1,R2);
and and14289(N23705,R3,R4);
and and14294(N23713,N23717,N23718);
and and14295(N23714,in1,R0);
and and14296(N23715,N23719,R2);
and and14297(N23716,R3,R4);
and and14302(N23724,N23728,in0);
and and14303(N23725,R0,R1);
and and14304(N23726,R2,R3);
and and14305(N23727,N23729,R5);
and and14310(N23734,N23738,in0);
and and14311(N23735,R0,R1);
and and14312(N23736,R2,R3);
and and14313(N23737,R4,R5);
and and14318(N23743,in0,N23747);
and and14319(N23744,N23748,N23749);
and and14320(N23745,R3,N23750);
and and14321(N23746,N23751,N23752);
and and14325(N23756,in0,N23760);
and and14326(N23757,N23761,R2);
and and14327(N23758,N23762,N23763);
and and14328(N23759,N23764,R7);
and and14332(N23768,in0,N23772);
and and14333(N23769,R1,N23773);
and and14334(N23770,R3,R5);
and and14335(N23771,N23774,N23775);
and and14339(N23779,in0,R0);
and and14340(N23780,N23783,R2);
and and14341(N23781,N23784,N23785);
and and14342(N23782,R5,N23786);
and and14346(N23790,in0,N23794);
and and14347(N23791,N23795,R2);
and and14348(N23792,R3,R4);
and and14349(N23793,N23796,R6);
and and14353(N23800,in0,R0);
and and14354(N23801,R1,N23804);
and and14355(N23802,R3,N23805);
and and14356(N23803,R5,N23806);
and and14360(N23810,in0,R0);
and and14361(N23811,N23814,R2);
and and14362(N23812,R3,R4);
and and14363(N23813,R6,R7);
and and14367(N23818,in0,R0);
and and14368(N23819,N23822,R3);
and and14369(N23820,R4,R5);
and and14370(N23821,R6,R7);
and and12343(N20642,R2,N20647);
and and12344(N20643,N20648,N20649);
and and12345(N20644,R6,N20650);
and and12353(N20658,N20665,N20666);
and and12354(N20659,N20667,N20668);
and and12362(N20676,N20684,R5);
and and12363(N20677,N20685,N20686);
and and12371(N20694,N20701,N20702);
and and12372(N20695,R6,N20703);
and and12380(N20711,R3,N20718);
and and12381(N20712,N20719,N20720);
and and12389(N20728,N20734,N20735);
and and12390(N20729,N20736,N20737);
and and12398(N20745,R3,N20752);
and and12399(N20746,N20753,N20754);
and and12407(N20762,N20769,N20770);
and and12408(N20763,R5,N20771);
and and12416(N20779,N20786,N20787);
and and12417(N20780,N20788,R7);
and and12425(N20796,N20803,N20804);
and and12426(N20797,R6,N20805);
and and12434(N20813,R3,R4);
and and12435(N20814,N20821,N20822);
and and12443(N20830,R4,R5);
and and12444(N20831,N20838,N20839);
and and12452(N20847,R3,N20855);
and and12453(N20848,R6,N20856);
and and12461(N20864,R3,N20872);
and and12462(N20865,N20873,R7);
and and12470(N20881,N20889,R4);
and and12471(N20882,R5,N20890);
and and12479(N20898,R3,N20905);
and and12480(N20899,N20906,N20907);
and and12488(N20915,N20920,N20921);
and and12489(N20916,N20922,N20923);
and and12497(N20931,N20936,N20937);
and and12498(N20932,N20938,N20939);
and and12506(N20947,R4,N20953);
and and12507(N20948,N20954,N20955);
and and12515(N20963,N20969,R4);
and and12516(N20964,N20970,N20971);
and and12524(N20979,N20985,R5);
and and12525(N20980,N20986,N20987);
and and12533(N20995,N21000,N21001);
and and12534(N20996,N21002,N21003);
and and12542(N21011,N21018,R5);
and and12543(N21012,R6,N21019);
and and12551(N21027,R3,N21033);
and and12552(N21028,N21034,N21035);
and and12560(N21043,N21050,R5);
and and12561(N21044,N21051,R7);
and and12569(N21059,R4,N21066);
and and12570(N21060,N21067,R7);
and and12578(N21075,N21082,R5);
and and12579(N21076,N21083,R7);
and and12587(N21091,N21098,N21099);
and and12588(N21092,R5,R6);
and and12596(N21107,R4,R5);
and and12597(N21108,N21114,N21115);
and and12605(N21123,R4,N21129);
and and12606(N21124,N21130,N21131);
and and12614(N21139,N21146,N21147);
and and12615(N21140,R6,R7);
and and12623(N21155,R4,N21162);
and and12624(N21156,R6,N21163);
and and12632(N21171,N21177,R5);
and and12633(N21172,N21178,N21179);
and and12641(N21187,N21194,R4);
and and12642(N21188,R5,N21195);
and and12650(N21203,N21209,R5);
and and12651(N21204,N21210,N21211);
and and12659(N21219,R3,N21225);
and and12660(N21220,N21226,N21227);
and and12668(N21235,N21241,N21242);
and and12669(N21236,N21243,R7);
and and12677(N21251,N21257,R5);
and and12678(N21252,N21258,N21259);
and and12686(N21267,N21274,N21275);
and and12687(N21268,R6,R7);
and and12695(N21283,R4,N21290);
and and12696(N21284,R6,N21291);
and and12704(N21299,R3,N21305);
and and12705(N21300,N21306,N21307);
and and12713(N21315,N21321,R5);
and and12714(N21316,N21322,R7);
and and12722(N21330,N21334,N21335);
and and12723(N21331,N21336,N21337);
and and12731(N21345,R3,N21351);
and and12732(N21346,N21352,R7);
and and12740(N21360,N21367,R5);
and and12741(N21361,R6,R7);
and and12749(N21375,N21381,R4);
and and12750(N21376,N21382,R6);
and and12758(N21390,N21395,N21396);
and and12759(N21391,N21397,R7);
and and12767(N21405,R4,N21410);
and and12768(N21406,N21411,N21412);
and and12776(N21420,N21426,R5);
and and12777(N21421,R6,N21427);
and and12785(N21435,N21441,R5);
and and12786(N21436,R6,N21442);
and and12794(N21450,N21456,R4);
and and12795(N21451,N21457,R7);
and and12803(N21465,R4,N21470);
and and12804(N21466,N21471,N21472);
and and12812(N21480,R3,R4);
and and12813(N21481,N21486,N21487);
and and12821(N21495,N21500,R5);
and and12822(N21496,N21501,N21502);
and and12830(N21510,R4,N21515);
and and12831(N21511,N21516,N21517);
and and12839(N21525,R4,N21530);
and and12840(N21526,N21531,N21532);
and and12848(N21540,R3,N21547);
and and12849(N21541,R6,R7);
and and12857(N21555,N21560,N21561);
and and12858(N21556,R6,N21562);
and and12866(N21570,N21576,R5);
and and12867(N21571,N21577,R7);
and and12875(N21585,N21590,R4);
and and12876(N21586,N21591,N21592);
and and12884(N21600,N21604,N21605);
and and12885(N21601,N21606,N21607);
and and12893(N21615,R3,R5);
and and12894(N21616,N21621,N21622);
and and12902(N21630,N21636,R5);
and and12903(N21631,R6,N21637);
and and12911(N21645,N21652,R5);
and and12912(N21646,R6,R7);
and and12920(N21660,R4,N21666);
and and12921(N21661,R6,N21667);
and and12929(N21675,N21681,N21682);
and and12930(N21676,R6,R7);
and and12938(N21690,R3,N21694);
and and12939(N21691,N21695,N21696);
and and12947(N21704,R4,R5);
and and12948(N21705,N21710,R7);
and and12956(N21718,R4,R5);
and and12957(N21719,N21724,R7);
and and12965(N21732,N21737,N21738);
and and12966(N21733,R6,R7);
and and12974(N21746,N21749,N21750);
and and12975(N21747,N21751,N21752);
and and12983(N21760,R3,N21764);
and and12984(N21761,N21765,N21766);
and and12992(N21774,R3,R4);
and and12993(N21775,N21779,N21780);
and and13001(N21788,R4,R5);
and and13002(N21789,N21793,N21794);
and and13010(N21802,R4,R5);
and and13011(N21803,N21807,N21808);
and and13019(N21816,N21821,R5);
and and13020(N21817,N21822,R7);
and and13028(N21830,N21835,R5);
and and13029(N21831,R6,N21836);
and and13037(N21844,N21849,R5);
and and13038(N21845,N21850,R7);
and and13046(N21858,R4,N21863);
and and13047(N21859,R6,N21864);
and and13055(N21872,N21876,R5);
and and13056(N21873,N21877,N21878);
and and13064(N21886,N21891,R5);
and and13065(N21887,N21892,R7);
and and13073(N21900,R4,N21905);
and and13074(N21901,N21906,R7);
and and13082(N21914,R4,N21920);
and and13083(N21915,R6,R7);
and and13091(N21928,N21933,N21934);
and and13092(N21929,R6,R7);
and and13100(N21942,R3,R4);
and and13101(N21943,N21947,N21948);
and and13109(N21956,N21961,N21962);
and and13110(N21957,R6,R7);
and and13118(N21970,N21975,R5);
and and13119(N21971,R6,N21976);
and and13127(N21984,R3,N21989);
and and13128(N21985,R6,N21990);
and and13136(N21998,N22002,R5);
and and13137(N21999,N22003,N22004);
and and13145(N22012,R3,R4);
and and13146(N22013,N22017,N22018);
and and13154(N22026,R3,N22030);
and and13155(N22027,N22031,N22032);
and and13163(N22040,R4,R5);
and and13164(N22041,N22045,N22046);
and and13172(N22054,N22058,N22059);
and and13173(N22055,R6,N22060);
and and13181(N22068,R4,N22073);
and and13182(N22069,N22074,R7);
and and13190(N22082,R4,R5);
and and13191(N22083,N22087,N22088);
and and13199(N22096,N22100,R5);
and and13200(N22097,N22101,N22102);
and and13208(N22110,R4,N22115);
and and13209(N22111,R6,N22116);
and and13217(N22124,R3,N22129);
and and13218(N22125,N22130,R7);
and and13226(N22138,N22144,R5);
and and13227(N22139,R6,R7);
and and13235(N22152,R3,R5);
and and13236(N22153,N22158,R7);
and and13244(N22166,R3,N22171);
and and13245(N22167,N22172,R6);
and and13253(N22180,R4,N22185);
and and13254(N22181,N22186,R7);
and and13262(N22194,R3,R5);
and and13263(N22195,R6,N22200);
and and13271(N22208,R4,R5);
and and13272(N22209,R6,N22213);
and and13280(N22221,R4,R5);
and and13281(N22222,R6,R7);
and and13289(N22234,R4,R5);
and and13290(N22235,N22239,R7);
and and13298(N22247,N22251,R5);
and and13299(N22248,R6,N22252);
and and13307(N22260,R4,R5);
and and13308(N22261,N22264,N22265);
and and13316(N22273,R4,N22277);
and and13317(N22274,N22278,R7);
and and13325(N22286,N22290,N22291);
and and13326(N22287,R6,R7);
and and13334(N22299,N22302,R5);
and and13335(N22300,N22303,N22304);
and and13343(N22312,R4,R5);
and and13344(N22313,N22317,R7);
and and13352(N22325,R4,R5);
and and13353(N22326,R6,R7);
and and13361(N22338,N22343,R5);
and and13362(N22339,R6,R7);
and and13370(N22351,R4,N22356);
and and13371(N22352,R6,R7);
and and13379(N22364,N22369,R5);
and and13380(N22365,R6,R7);
and and13388(N22377,R4,N22380);
and and13389(N22378,N22381,N22382);
and and13397(N22390,R4,R5);
and and13398(N22391,R6,R7);
and and13406(N22403,R4,R5);
and and13407(N22404,N22408,R7);
and and13415(N22416,N22419,R4);
and and13416(N22417,N22420,N22421);
and and13424(N22429,N22433,N22434);
and and13425(N22430,R6,R7);
and and13433(N22442,R3,N22447);
and and13434(N22443,R6,R7);
and and13442(N22455,R4,R5);
and and13443(N22456,N22460,R7);
and and13451(N22468,N22473,R5);
and and13452(N22469,R6,R7);
and and13460(N22481,R4,R5);
and and13461(N22482,N22486,R7);
and and13469(N22494,N22499,R4);
and and13470(N22495,R5,R7);
and and13478(N22507,R3,R4);
and and13479(N22508,R5,R6);
and and13487(N22520,R4,N22524);
and and13488(N22521,N22525,R7);
and and13496(N22533,N22537,R5);
and and13497(N22534,N22538,R7);
and and13505(N22546,N22550,R5);
and and13506(N22547,N22551,R7);
and and13514(N22559,N22563,N22564);
and and13515(N22560,R6,R7);
and and13523(N22572,R3,N22577);
and and13524(N22573,R5,R6);
and and13532(N22585,R3,N22589);
and and13533(N22586,R5,N22590);
and and13541(N22598,N22602,N22603);
and and13542(N22599,R6,R7);
and and13550(N22611,N22615,R5);
and and13551(N22612,R6,N22616);
and and13559(N22624,N22628,R5);
and and13560(N22625,N22629,R7);
and and13568(N22637,R3,N22642);
and and13569(N22638,R6,R7);
and and13577(N22650,R3,R4);
and and13578(N22651,R5,N22655);
and and13586(N22663,R3,R4);
and and13587(N22664,R5,N22668);
and and13595(N22676,N22680,R5);
and and13596(N22677,R6,N22681);
and and13604(N22689,R4,R5);
and and13605(N22690,N22692,N22693);
and and13613(N22701,R3,R4);
and and13614(N22702,R5,N22705);
and and13622(N22713,R3,R4);
and and13623(N22714,R5,R6);
and and13631(N22725,R4,R5);
and and13632(N22726,R6,R7);
and and13640(N22737,R3,R4);
and and13641(N22738,R5,R7);
and and13649(N22749,R4,N22753);
and and13650(N22750,R6,R7);
and and13658(N22761,N22765,R5);
and and13659(N22762,R6,R7);
and and13667(N22773,R3,R4);
and and13668(N22774,N22777,R7);
and and13676(N22785,R3,R5);
and and13677(N22786,N22789,R7);
and and13685(N22797,R4,R5);
and and13686(N22798,R6,R7);
and and13694(N22809,R3,R4);
and and13695(N22810,R5,R7);
and and13703(N22821,R4,R5);
and and13704(N22822,R6,R7);
and and13712(N22833,R4,R5);
and and13713(N22834,R6,N22837);
and and13721(N22845,R4,R5);
and and13722(N22846,R6,R7);
and and13730(N22857,R4,R5);
and and13731(N22858,R6,N22861);
and and13739(N22869,R4,R5);
and and13740(N22870,N22873,R7);
and and13748(N22881,N22884,N22885);
and and13749(N22882,R6,R7);
and and13757(N22893,N22896,R5);
and and13758(N22894,R6,N22897);
and and13766(N22905,R3,R4);
and and13767(N22906,N22908,N22909);
and and13775(N22917,R4,N22919);
and and13776(N22918,N22920,N22921);
and and13784(N22929,N22932,R4);
and and13785(N22930,R5,R6);
and and13793(N22940,R4,R5);
and and13794(N22941,R6,R7);
and and13802(N22951,R4,N22954);
and and13803(N22952,R6,R7);
and and13811(N22962,R4,N22965);
and and13812(N22963,R6,R7);
and and13820(N22973,N22975,N22976);
and and13821(N22974,R6,R7);
and and13829(N22984,N22986,N22987);
and and13830(N22985,R6,R7);
and and13838(N22995,R4,R5);
and and13839(N22996,R6,R7);
and and13847(N23006,R4,N23009);
and and13848(N23007,R6,R7);
and and13856(N23017,R3,R5);
and and13857(N23018,R6,R7);
and and13865(N23027,R4,R5);
and and13866(N23028,N23029,R7);
and and13874(N23037,N23044,N23045);
and and13882(N23053,N23060,N23061);
and and13890(N23069,N23077,R7);
and and13898(N23085,N23091,N23092);
and and13906(N23100,N23106,N23107);
and and13914(N23115,N23121,N23122);
and and13922(N23130,N23135,N23136);
and and13930(N23144,N23149,N23150);
and and13938(N23158,R6,N23164);
and and13946(N23172,N23177,N23178);
and and13954(N23186,N23191,N23192);
and and13962(N23200,N23206,R7);
and and13970(N23214,N23220,R7);
and and13978(N23228,N23234,R7);
and and13986(N23242,N23246,N23247);
and and13994(N23255,N23260,R7);
and and14002(N23268,N23272,N23273);
and and14010(N23281,R6,N23286);
and and14018(N23294,N23298,N23299);
and and14026(N23307,R6,R7);
and and14034(N23320,R5,R6);
and and14042(N23333,R6,N23338);
and and14050(N23346,R4,N23351);
and and14058(N23359,R5,R6);
and and14066(N23372,R5,R6);
and and14074(N23385,N23390,R6);
and and14082(N23398,R6,N23403);
and and14090(N23411,N23416,R7);
and and14098(N23424,R5,N23429);
and and14106(N23437,R6,N23442);
and and14114(N23450,R6,N23454);
and and14122(N23462,N23465,N23466);
and and14130(N23474,N23477,N23478);
and and14138(N23486,N23490,R7);
and and14146(N23498,R6,N23502);
and and14154(N23510,N23514,R7);
and and14162(N23522,R5,N23526);
and and14170(N23534,N23538,R7);
and and14178(N23546,N23550,R7);
and and14186(N23558,N23562,R7);
and and14194(N23570,R6,R7);
and and14202(N23582,N23585,N23586);
and and14210(N23594,N23598,R7);
and and14218(N23606,R6,R7);
and and14226(N23618,R6,R7);
and and14234(N23629,R6,N23632);
and and14242(N23640,R6,N23643);
and and14250(N23651,N23654,R7);
and and14258(N23662,N23665,R7);
and and14266(N23673,R6,N23676);
and and14274(N23684,R6,N23687);
and and14282(N23695,R5,R6);
and and14290(N23706,N23708,N23709);
and and14298(N23717,R6,N23720);
and and14306(N23728,R6,N23730);
and and14314(N23738,N23739,R7);
and and14371(N24191,N24192,N24193);
and and14380(N24209,N24210,N24211);
and and14389(N24227,N24228,N24229);
and and14398(N24245,N24246,N24247);
and and14407(N24263,N24264,N24265);
and and14416(N24281,N24282,N24283);
and and14425(N24299,N24300,N24301);
and and14434(N24317,N24318,N24319);
and and14443(N24334,N24335,N24336);
and and14452(N24351,N24352,N24353);
and and14461(N24368,N24369,N24370);
and and14470(N24385,N24386,N24387);
and and14479(N24402,N24403,N24404);
and and14488(N24419,N24420,N24421);
and and14497(N24436,N24437,N24438);
and and14506(N24453,N24454,N24455);
and and14515(N24470,N24471,N24472);
and and14524(N24486,N24487,N24488);
and and14533(N24502,N24503,N24504);
and and14542(N24518,N24519,N24520);
and and14551(N24534,N24535,N24536);
and and14560(N24550,N24551,N24552);
and and14569(N24566,N24567,N24568);
and and14578(N24582,N24583,N24584);
and and14587(N24598,N24599,N24600);
and and14596(N24614,N24615,N24616);
and and14605(N24630,N24631,N24632);
and and14614(N24646,N24647,N24648);
and and14623(N24662,N24663,N24664);
and and14632(N24678,N24679,N24680);
and and14641(N24694,N24695,N24696);
and and14650(N24710,N24711,N24712);
and and14659(N24726,N24727,N24728);
and and14668(N24742,N24743,N24744);
and and14677(N24758,N24759,N24760);
and and14686(N24774,N24775,N24776);
and and14695(N24790,N24791,N24792);
and and14704(N24806,N24807,N24808);
and and14713(N24822,N24823,N24824);
and and14722(N24838,N24839,N24840);
and and14731(N24854,N24855,N24856);
and and14740(N24870,N24871,N24872);
and and14749(N24886,N24887,N24888);
and and14758(N24902,N24903,N24904);
and and14767(N24918,N24919,N24920);
and and14776(N24934,N24935,N24936);
and and14785(N24950,N24951,N24952);
and and14794(N24965,N24966,N24967);
and and14803(N24980,N24981,N24982);
and and14812(N24995,N24996,N24997);
and and14821(N25010,N25011,N25012);
and and14830(N25025,N25026,N25027);
and and14839(N25040,N25041,N25042);
and and14848(N25055,N25056,N25057);
and and14857(N25070,N25071,N25072);
and and14866(N25085,N25086,N25087);
and and14875(N25100,N25101,N25102);
and and14884(N25115,N25116,N25117);
and and14893(N25130,N25131,N25132);
and and14902(N25145,N25146,N25147);
and and14911(N25160,N25161,N25162);
and and14920(N25175,N25176,N25177);
and and14929(N25190,N25191,N25192);
and and14938(N25205,N25206,N25207);
and and14947(N25220,N25221,N25222);
and and14956(N25235,N25236,N25237);
and and14965(N25250,N25251,N25252);
and and14974(N25265,N25266,N25267);
and and14983(N25280,N25281,N25282);
and and14992(N25295,N25296,N25297);
and and15001(N25310,N25311,N25312);
and and15010(N25325,N25326,N25327);
and and15019(N25340,N25341,N25342);
and and15028(N25355,N25356,N25357);
and and15037(N25370,N25371,N25372);
and and15046(N25385,N25386,N25387);
and and15055(N25400,N25401,N25402);
and and15064(N25415,N25416,N25417);
and and15073(N25429,N25430,N25431);
and and15082(N25443,N25444,N25445);
and and15091(N25457,N25458,N25459);
and and15100(N25471,N25472,N25473);
and and15109(N25485,N25486,N25487);
and and15118(N25499,N25500,N25501);
and and15127(N25513,N25514,N25515);
and and15136(N25527,N25528,N25529);
and and15145(N25541,N25542,N25543);
and and15154(N25555,N25556,N25557);
and and15163(N25569,N25570,N25571);
and and15172(N25583,N25584,N25585);
and and15181(N25597,N25598,N25599);
and and15190(N25611,N25612,N25613);
and and15199(N25625,N25626,N25627);
and and15208(N25639,N25640,N25641);
and and15217(N25653,N25654,N25655);
and and15226(N25667,N25668,N25669);
and and15235(N25681,N25682,N25683);
and and15244(N25695,N25696,N25697);
and and15253(N25709,N25710,N25711);
and and15262(N25723,N25724,N25725);
and and15271(N25737,N25738,N25739);
and and15280(N25751,N25752,N25753);
and and15289(N25765,N25766,N25767);
and and15298(N25779,N25780,N25781);
and and15307(N25793,N25794,N25795);
and and15316(N25807,N25808,N25809);
and and15325(N25821,N25822,N25823);
and and15334(N25835,N25836,N25837);
and and15343(N25849,N25850,N25851);
and and15352(N25863,N25864,N25865);
and and15361(N25877,N25878,N25879);
and and15370(N25891,N25892,N25893);
and and15379(N25905,N25906,N25907);
and and15388(N25919,N25920,N25921);
and and15397(N25933,N25934,N25935);
and and15406(N25947,N25948,N25949);
and and15415(N25961,N25962,N25963);
and and15424(N25975,N25976,N25977);
and and15433(N25989,N25990,N25991);
and and15442(N26003,N26004,N26005);
and and15451(N26017,N26018,N26019);
and and15460(N26031,N26032,N26033);
and and15469(N26045,N26046,N26047);
and and15478(N26059,N26060,N26061);
and and15487(N26073,N26074,N26075);
and and15496(N26087,N26088,N26089);
and and15505(N26101,N26102,N26103);
and and15514(N26115,N26116,N26117);
and and15523(N26129,N26130,N26131);
and and15532(N26143,N26144,N26145);
and and15541(N26157,N26158,N26159);
and and15550(N26171,N26172,N26173);
and and15559(N26184,N26185,N26186);
and and15568(N26197,N26198,N26199);
and and15577(N26210,N26211,N26212);
and and15586(N26223,N26224,N26225);
and and15595(N26236,N26237,N26238);
and and15604(N26249,N26250,N26251);
and and15613(N26262,N26263,N26264);
and and15622(N26275,N26276,N26277);
and and15631(N26288,N26289,N26290);
and and15640(N26301,N26302,N26303);
and and15649(N26314,N26315,N26316);
and and15658(N26327,N26328,N26329);
and and15667(N26340,N26341,N26342);
and and15676(N26353,N26354,N26355);
and and15685(N26366,N26367,N26368);
and and15694(N26379,N26380,N26381);
and and15703(N26392,N26393,N26394);
and and15712(N26405,N26406,N26407);
and and15721(N26418,N26419,N26420);
and and15730(N26431,N26432,N26433);
and and15739(N26444,N26445,N26446);
and and15748(N26457,N26458,N26459);
and and15757(N26470,N26471,N26472);
and and15766(N26483,N26484,N26485);
and and15775(N26496,N26497,N26498);
and and15784(N26509,N26510,N26511);
and and15793(N26522,N26523,N26524);
and and15802(N26535,N26536,N26537);
and and15811(N26548,N26549,N26550);
and and15820(N26561,N26562,N26563);
and and15829(N26574,N26575,N26576);
and and15838(N26587,N26588,N26589);
and and15847(N26600,N26601,N26602);
and and15856(N26613,N26614,N26615);
and and15865(N26625,N26626,N26627);
and and15874(N26637,N26638,N26639);
and and15883(N26649,N26650,N26651);
and and15892(N26661,N26662,N26663);
and and15901(N26673,N26674,N26675);
and and15910(N26685,N26686,N26687);
and and15919(N26697,N26698,N26699);
and and15928(N26709,N26710,N26711);
and and15937(N26721,N26722,N26723);
and and15946(N26733,N26734,N26735);
and and15955(N26745,N26746,N26747);
and and15964(N26757,N26758,N26759);
and and15973(N26769,N26770,N26771);
and and15982(N26781,N26782,N26783);
and and15991(N26793,N26794,N26795);
and and16000(N26805,N26806,N26807);
and and16009(N26817,N26818,N26819);
and and16018(N26829,N26830,N26831);
and and16027(N26841,N26842,N26843);
and and16036(N26853,N26854,N26855);
and and16045(N26865,N26866,N26867);
and and16054(N26877,N26878,N26879);
and and16063(N26889,N26890,N26891);
and and16072(N26901,N26902,N26903);
and and16081(N26913,N26914,N26915);
and and16090(N26925,N26926,N26927);
and and16099(N26937,N26938,N26939);
and and16108(N26949,N26950,N26951);
and and16117(N26961,N26962,N26963);
and and16126(N26973,N26974,N26975);
and and16135(N26985,N26986,N26987);
and and16144(N26997,N26998,N26999);
and and16153(N27009,N27010,N27011);
and and16162(N27021,N27022,N27023);
and and16171(N27033,N27034,N27035);
and and16180(N27045,N27046,N27047);
and and16189(N27057,N27058,N27059);
and and16198(N27068,N27069,N27070);
and and16207(N27079,N27080,N27081);
and and16216(N27090,N27091,N27092);
and and16225(N27101,N27102,N27103);
and and16234(N27111,N27112,N27113);
and and16243(N27121,N27122,N27123);
and and16252(N27131,N27132,N27133);
and and16261(N27141,N27142,N27143);
and and16270(N27151,N27152,N27153);
and and16279(N27161,N27162,N27163);
and and16288(N27171,N27172,N27173);
and and16297(N27181,N27182,N27183);
and and16306(N27191,N27192,N27193);
and and16315(N27201,N27202,N27203);
and and16323(N27217,N27218,N27219);
and and16331(N27233,N27234,N27235);
and and16339(N27248,N27249,N27250);
and and16347(N27263,N27264,N27265);
and and16355(N27278,N27279,N27280);
and and16363(N27292,N27293,N27294);
and and16371(N27306,N27307,N27308);
and and16379(N27320,N27321,N27322);
and and16387(N27334,N27335,N27336);
and and16395(N27348,N27349,N27350);
and and16403(N27362,N27363,N27364);
and and16411(N27376,N27377,N27378);
and and16419(N27390,N27391,N27392);
and and16427(N27404,N27405,N27406);
and and16435(N27418,N27419,N27420);
and and16443(N27432,N27433,N27434);
and and16451(N27446,N27447,N27448);
and and16459(N27460,N27461,N27462);
and and16467(N27474,N27475,N27476);
and and16475(N27488,N27489,N27490);
and and16483(N27502,N27503,N27504);
and and16491(N27516,N27517,N27518);
and and16499(N27530,N27531,N27532);
and and16507(N27544,N27545,N27546);
and and16515(N27558,N27559,N27560);
and and16523(N27572,N27573,N27574);
and and16531(N27586,N27587,N27588);
and and16539(N27600,N27601,N27602);
and and16547(N27613,N27614,N27615);
and and16555(N27626,N27627,N27628);
and and16563(N27639,N27640,N27641);
and and16571(N27652,N27653,N27654);
and and16579(N27665,N27666,N27667);
and and16587(N27678,N27679,N27680);
and and16595(N27691,N27692,N27693);
and and16603(N27704,N27705,N27706);
and and16611(N27717,N27718,N27719);
and and16619(N27730,N27731,N27732);
and and16627(N27743,N27744,N27745);
and and16635(N27756,N27757,N27758);
and and16643(N27769,N27770,N27771);
and and16651(N27782,N27783,N27784);
and and16659(N27795,N27796,N27797);
and and16667(N27808,N27809,N27810);
and and16675(N27821,N27822,N27823);
and and16683(N27834,N27835,N27836);
and and16691(N27847,N27848,N27849);
and and16699(N27860,N27861,N27862);
and and16707(N27873,N27874,N27875);
and and16715(N27886,N27887,N27888);
and and16723(N27899,N27900,N27901);
and and16731(N27912,N27913,N27914);
and and16739(N27925,N27926,N27927);
and and16747(N27938,N27939,N27940);
and and16755(N27951,N27952,N27953);
and and16763(N27964,N27965,N27966);
and and16771(N27977,N27978,N27979);
and and16779(N27990,N27991,N27992);
and and16787(N28003,N28004,N28005);
and and16795(N28016,N28017,N28018);
and and16803(N28029,N28030,N28031);
and and16811(N28042,N28043,N28044);
and and16819(N28055,N28056,N28057);
and and16827(N28068,N28069,N28070);
and and16835(N28081,N28082,N28083);
and and16843(N28094,N28095,N28096);
and and16851(N28106,N28107,N28108);
and and16859(N28118,N28119,N28120);
and and16867(N28130,N28131,N28132);
and and16875(N28142,N28143,N28144);
and and16883(N28154,N28155,N28156);
and and16891(N28166,N28167,N28168);
and and16899(N28178,N28179,N28180);
and and16907(N28190,N28191,N28192);
and and16915(N28202,N28203,N28204);
and and16923(N28214,N28215,N28216);
and and16931(N28226,N28227,N28228);
and and16939(N28238,N28239,N28240);
and and16947(N28250,N28251,N28252);
and and16955(N28262,N28263,N28264);
and and16963(N28274,N28275,N28276);
and and16971(N28286,N28287,N28288);
and and16979(N28298,N28299,N28300);
and and16987(N28310,N28311,N28312);
and and16995(N28322,N28323,N28324);
and and17003(N28334,N28335,N28336);
and and17011(N28346,N28347,N28348);
and and17019(N28358,N28359,N28360);
and and17027(N28370,N28371,N28372);
and and17035(N28382,N28383,N28384);
and and17043(N28394,N28395,N28396);
and and17051(N28406,N28407,N28408);
and and17059(N28418,N28419,N28420);
and and17067(N28430,N28431,N28432);
and and17075(N28442,N28443,N28444);
and and17083(N28454,N28455,N28456);
and and17091(N28465,N28466,N28467);
and and17099(N28476,N28477,N28478);
and and17107(N28487,N28488,N28489);
and and17115(N28498,N28499,N28500);
and and17123(N28509,N28510,N28511);
and and17131(N28520,N28521,N28522);
and and17139(N28531,N28532,N28533);
and and17147(N28542,N28543,N28544);
and and17155(N28553,N28554,N28555);
and and17163(N28564,N28565,N28566);
and and17171(N28575,N28576,N28577);
and and17179(N28586,N28587,N28588);
and and17187(N28597,N28598,N28599);
and and17195(N28608,N28609,N28610);
and and17203(N28619,N28620,N28621);
and and17211(N28630,N28631,N28632);
and and17219(N28641,N28642,N28643);
and and17227(N28652,N28653,N28654);
and and17235(N28663,N28664,N28665);
and and17243(N28674,N28675,N28676);
and and17251(N28685,N28686,N28687);
and and17259(N28695,N28696,N28697);
and and17267(N28705,N28706,N28707);
and and17275(N28715,N28716,N28717);
and and17283(N28725,N28726,N28727);
and and17291(N28735,N28736,N28737);
and and17299(N28745,N28746,N28747);
and and17307(N28755,N28756,N28757);
and and17315(N28765,N28766,N28767);
and and17323(N28775,N28776,N28777);
and and17331(N28785,N28786,N28787);
and and17339(N28795,N28796,N28797);
and and17347(N28805,N28806,N28807);
and and17355(N28815,N28816,N28817);
and and17363(N28825,N28826,N28827);
and and17371(N28835,N28836,N28837);
and and17379(N28844,N28845,N28846);
and and17387(N28852,N28853,N28854);
and and17395(N28860,N28861,N28862);
and and17402(N28873,N28874,N28875);
and and17409(N28885,N28886,N28887);
and and17416(N28897,N28898,N28899);
and and17423(N28909,N28910,N28911);
and and17430(N28921,N28922,N28923);
and and17437(N28932,N28933,N28934);
and and17444(N28943,N28944,N28945);
and and17451(N28954,N28955,N28956);
and and17458(N28965,N28966,N28967);
and and17465(N28975,N28976,N28977);
and and17472(N28985,N28986,N28987);
and and17479(N28995,N28996,N28997);
and and17486(N29005,N29006,N29007);
and and17493(N29015,N29016,N29017);
and and17500(N29025,N29026,N29027);
and and17507(N29035,N29036,N29037);
and and17514(N29044,N29045,N29046);
and and14372(N24192,N24194,N24195);
and and14373(N24193,N24196,N24197);
and and14381(N24210,N24212,N24213);
and and14382(N24211,N24214,N24215);
and and14390(N24228,N24230,N24231);
and and14391(N24229,N24232,N24233);
and and14399(N24246,N24248,N24249);
and and14400(N24247,N24250,N24251);
and and14408(N24264,N24266,N24267);
and and14409(N24265,N24268,N24269);
and and14417(N24282,N24284,N24285);
and and14418(N24283,N24286,N24287);
and and14426(N24300,N24302,N24303);
and and14427(N24301,N24304,N24305);
and and14435(N24318,N24320,N24321);
and and14436(N24319,N24322,N24323);
and and14444(N24335,N24337,N24338);
and and14445(N24336,N24339,N24340);
and and14453(N24352,N24354,N24355);
and and14454(N24353,N24356,N24357);
and and14462(N24369,N24371,N24372);
and and14463(N24370,N24373,N24374);
and and14471(N24386,N24388,N24389);
and and14472(N24387,N24390,N24391);
and and14480(N24403,N24405,N24406);
and and14481(N24404,N24407,N24408);
and and14489(N24420,N24422,N24423);
and and14490(N24421,N24424,N24425);
and and14498(N24437,N24439,N24440);
and and14499(N24438,N24441,N24442);
and and14507(N24454,N24456,N24457);
and and14508(N24455,N24458,N24459);
and and14516(N24471,N24473,N24474);
and and14517(N24472,N24475,N24476);
and and14525(N24487,N24489,N24490);
and and14526(N24488,N24491,N24492);
and and14534(N24503,N24505,N24506);
and and14535(N24504,N24507,N24508);
and and14543(N24519,N24521,N24522);
and and14544(N24520,N24523,N24524);
and and14552(N24535,N24537,N24538);
and and14553(N24536,N24539,N24540);
and and14561(N24551,N24553,N24554);
and and14562(N24552,N24555,N24556);
and and14570(N24567,N24569,N24570);
and and14571(N24568,N24571,N24572);
and and14579(N24583,N24585,N24586);
and and14580(N24584,N24587,N24588);
and and14588(N24599,N24601,N24602);
and and14589(N24600,N24603,N24604);
and and14597(N24615,N24617,N24618);
and and14598(N24616,N24619,N24620);
and and14606(N24631,N24633,N24634);
and and14607(N24632,N24635,N24636);
and and14615(N24647,N24649,N24650);
and and14616(N24648,N24651,N24652);
and and14624(N24663,N24665,N24666);
and and14625(N24664,N24667,N24668);
and and14633(N24679,N24681,N24682);
and and14634(N24680,N24683,N24684);
and and14642(N24695,N24697,N24698);
and and14643(N24696,N24699,N24700);
and and14651(N24711,N24713,N24714);
and and14652(N24712,N24715,N24716);
and and14660(N24727,N24729,N24730);
and and14661(N24728,N24731,N24732);
and and14669(N24743,N24745,N24746);
and and14670(N24744,N24747,N24748);
and and14678(N24759,N24761,N24762);
and and14679(N24760,N24763,N24764);
and and14687(N24775,N24777,N24778);
and and14688(N24776,N24779,N24780);
and and14696(N24791,N24793,N24794);
and and14697(N24792,N24795,N24796);
and and14705(N24807,N24809,N24810);
and and14706(N24808,N24811,N24812);
and and14714(N24823,N24825,N24826);
and and14715(N24824,N24827,N24828);
and and14723(N24839,N24841,N24842);
and and14724(N24840,N24843,N24844);
and and14732(N24855,N24857,N24858);
and and14733(N24856,N24859,N24860);
and and14741(N24871,N24873,N24874);
and and14742(N24872,N24875,N24876);
and and14750(N24887,N24889,N24890);
and and14751(N24888,N24891,N24892);
and and14759(N24903,N24905,N24906);
and and14760(N24904,N24907,N24908);
and and14768(N24919,N24921,N24922);
and and14769(N24920,N24923,N24924);
and and14777(N24935,N24937,N24938);
and and14778(N24936,N24939,N24940);
and and14786(N24951,N24953,N24954);
and and14787(N24952,N24955,N24956);
and and14795(N24966,N24968,N24969);
and and14796(N24967,N24970,N24971);
and and14804(N24981,N24983,N24984);
and and14805(N24982,N24985,N24986);
and and14813(N24996,N24998,N24999);
and and14814(N24997,N25000,N25001);
and and14822(N25011,N25013,N25014);
and and14823(N25012,N25015,N25016);
and and14831(N25026,N25028,N25029);
and and14832(N25027,N25030,N25031);
and and14840(N25041,N25043,N25044);
and and14841(N25042,N25045,N25046);
and and14849(N25056,N25058,N25059);
and and14850(N25057,N25060,N25061);
and and14858(N25071,N25073,N25074);
and and14859(N25072,N25075,N25076);
and and14867(N25086,N25088,N25089);
and and14868(N25087,N25090,N25091);
and and14876(N25101,N25103,N25104);
and and14877(N25102,N25105,N25106);
and and14885(N25116,N25118,N25119);
and and14886(N25117,N25120,N25121);
and and14894(N25131,N25133,N25134);
and and14895(N25132,N25135,N25136);
and and14903(N25146,N25148,N25149);
and and14904(N25147,N25150,N25151);
and and14912(N25161,N25163,N25164);
and and14913(N25162,N25165,N25166);
and and14921(N25176,N25178,N25179);
and and14922(N25177,N25180,N25181);
and and14930(N25191,N25193,N25194);
and and14931(N25192,N25195,N25196);
and and14939(N25206,N25208,N25209);
and and14940(N25207,N25210,N25211);
and and14948(N25221,N25223,N25224);
and and14949(N25222,N25225,N25226);
and and14957(N25236,N25238,N25239);
and and14958(N25237,N25240,N25241);
and and14966(N25251,N25253,N25254);
and and14967(N25252,N25255,N25256);
and and14975(N25266,N25268,N25269);
and and14976(N25267,N25270,N25271);
and and14984(N25281,N25283,N25284);
and and14985(N25282,N25285,N25286);
and and14993(N25296,N25298,N25299);
and and14994(N25297,N25300,N25301);
and and15002(N25311,N25313,N25314);
and and15003(N25312,N25315,N25316);
and and15011(N25326,N25328,N25329);
and and15012(N25327,N25330,N25331);
and and15020(N25341,N25343,N25344);
and and15021(N25342,N25345,N25346);
and and15029(N25356,N25358,N25359);
and and15030(N25357,N25360,N25361);
and and15038(N25371,N25373,N25374);
and and15039(N25372,N25375,N25376);
and and15047(N25386,N25388,N25389);
and and15048(N25387,N25390,N25391);
and and15056(N25401,N25403,N25404);
and and15057(N25402,N25405,N25406);
and and15065(N25416,N25418,N25419);
and and15066(N25417,N25420,N25421);
and and15074(N25430,N25432,N25433);
and and15075(N25431,N25434,N25435);
and and15083(N25444,N25446,N25447);
and and15084(N25445,N25448,N25449);
and and15092(N25458,N25460,N25461);
and and15093(N25459,N25462,N25463);
and and15101(N25472,N25474,N25475);
and and15102(N25473,N25476,N25477);
and and15110(N25486,N25488,N25489);
and and15111(N25487,N25490,N25491);
and and15119(N25500,N25502,N25503);
and and15120(N25501,N25504,N25505);
and and15128(N25514,N25516,N25517);
and and15129(N25515,N25518,N25519);
and and15137(N25528,N25530,N25531);
and and15138(N25529,N25532,N25533);
and and15146(N25542,N25544,N25545);
and and15147(N25543,N25546,N25547);
and and15155(N25556,N25558,N25559);
and and15156(N25557,N25560,N25561);
and and15164(N25570,N25572,N25573);
and and15165(N25571,N25574,N25575);
and and15173(N25584,N25586,N25587);
and and15174(N25585,N25588,N25589);
and and15182(N25598,N25600,N25601);
and and15183(N25599,N25602,N25603);
and and15191(N25612,N25614,N25615);
and and15192(N25613,N25616,N25617);
and and15200(N25626,N25628,N25629);
and and15201(N25627,N25630,N25631);
and and15209(N25640,N25642,N25643);
and and15210(N25641,N25644,N25645);
and and15218(N25654,N25656,N25657);
and and15219(N25655,N25658,N25659);
and and15227(N25668,N25670,N25671);
and and15228(N25669,N25672,N25673);
and and15236(N25682,N25684,N25685);
and and15237(N25683,N25686,N25687);
and and15245(N25696,N25698,N25699);
and and15246(N25697,N25700,N25701);
and and15254(N25710,N25712,N25713);
and and15255(N25711,N25714,N25715);
and and15263(N25724,N25726,N25727);
and and15264(N25725,N25728,N25729);
and and15272(N25738,N25740,N25741);
and and15273(N25739,N25742,N25743);
and and15281(N25752,N25754,N25755);
and and15282(N25753,N25756,N25757);
and and15290(N25766,N25768,N25769);
and and15291(N25767,N25770,N25771);
and and15299(N25780,N25782,N25783);
and and15300(N25781,N25784,N25785);
and and15308(N25794,N25796,N25797);
and and15309(N25795,N25798,N25799);
and and15317(N25808,N25810,N25811);
and and15318(N25809,N25812,N25813);
and and15326(N25822,N25824,N25825);
and and15327(N25823,N25826,N25827);
and and15335(N25836,N25838,N25839);
and and15336(N25837,N25840,N25841);
and and15344(N25850,N25852,N25853);
and and15345(N25851,N25854,N25855);
and and15353(N25864,N25866,N25867);
and and15354(N25865,N25868,N25869);
and and15362(N25878,N25880,N25881);
and and15363(N25879,N25882,N25883);
and and15371(N25892,N25894,N25895);
and and15372(N25893,N25896,N25897);
and and15380(N25906,N25908,N25909);
and and15381(N25907,N25910,N25911);
and and15389(N25920,N25922,N25923);
and and15390(N25921,N25924,N25925);
and and15398(N25934,N25936,N25937);
and and15399(N25935,N25938,N25939);
and and15407(N25948,N25950,N25951);
and and15408(N25949,N25952,N25953);
and and15416(N25962,N25964,N25965);
and and15417(N25963,N25966,N25967);
and and15425(N25976,N25978,N25979);
and and15426(N25977,N25980,N25981);
and and15434(N25990,N25992,N25993);
and and15435(N25991,N25994,N25995);
and and15443(N26004,N26006,N26007);
and and15444(N26005,N26008,N26009);
and and15452(N26018,N26020,N26021);
and and15453(N26019,N26022,N26023);
and and15461(N26032,N26034,N26035);
and and15462(N26033,N26036,N26037);
and and15470(N26046,N26048,N26049);
and and15471(N26047,N26050,N26051);
and and15479(N26060,N26062,N26063);
and and15480(N26061,N26064,N26065);
and and15488(N26074,N26076,N26077);
and and15489(N26075,N26078,N26079);
and and15497(N26088,N26090,N26091);
and and15498(N26089,N26092,N26093);
and and15506(N26102,N26104,N26105);
and and15507(N26103,N26106,N26107);
and and15515(N26116,N26118,N26119);
and and15516(N26117,N26120,N26121);
and and15524(N26130,N26132,N26133);
and and15525(N26131,N26134,N26135);
and and15533(N26144,N26146,N26147);
and and15534(N26145,N26148,N26149);
and and15542(N26158,N26160,N26161);
and and15543(N26159,N26162,N26163);
and and15551(N26172,N26174,N26175);
and and15552(N26173,N26176,N26177);
and and15560(N26185,N26187,N26188);
and and15561(N26186,N26189,N26190);
and and15569(N26198,N26200,N26201);
and and15570(N26199,N26202,N26203);
and and15578(N26211,N26213,N26214);
and and15579(N26212,N26215,N26216);
and and15587(N26224,N26226,N26227);
and and15588(N26225,N26228,N26229);
and and15596(N26237,N26239,N26240);
and and15597(N26238,N26241,N26242);
and and15605(N26250,N26252,N26253);
and and15606(N26251,N26254,N26255);
and and15614(N26263,N26265,N26266);
and and15615(N26264,N26267,N26268);
and and15623(N26276,N26278,N26279);
and and15624(N26277,N26280,N26281);
and and15632(N26289,N26291,N26292);
and and15633(N26290,N26293,N26294);
and and15641(N26302,N26304,N26305);
and and15642(N26303,N26306,N26307);
and and15650(N26315,N26317,N26318);
and and15651(N26316,N26319,N26320);
and and15659(N26328,N26330,N26331);
and and15660(N26329,N26332,N26333);
and and15668(N26341,N26343,N26344);
and and15669(N26342,N26345,N26346);
and and15677(N26354,N26356,N26357);
and and15678(N26355,N26358,N26359);
and and15686(N26367,N26369,N26370);
and and15687(N26368,N26371,N26372);
and and15695(N26380,N26382,N26383);
and and15696(N26381,N26384,N26385);
and and15704(N26393,N26395,N26396);
and and15705(N26394,N26397,N26398);
and and15713(N26406,N26408,N26409);
and and15714(N26407,N26410,N26411);
and and15722(N26419,N26421,N26422);
and and15723(N26420,N26423,N26424);
and and15731(N26432,N26434,N26435);
and and15732(N26433,N26436,N26437);
and and15740(N26445,N26447,N26448);
and and15741(N26446,N26449,N26450);
and and15749(N26458,N26460,N26461);
and and15750(N26459,N26462,N26463);
and and15758(N26471,N26473,N26474);
and and15759(N26472,N26475,N26476);
and and15767(N26484,N26486,N26487);
and and15768(N26485,N26488,N26489);
and and15776(N26497,N26499,N26500);
and and15777(N26498,N26501,N26502);
and and15785(N26510,N26512,N26513);
and and15786(N26511,N26514,N26515);
and and15794(N26523,N26525,N26526);
and and15795(N26524,N26527,N26528);
and and15803(N26536,N26538,N26539);
and and15804(N26537,N26540,N26541);
and and15812(N26549,N26551,N26552);
and and15813(N26550,N26553,N26554);
and and15821(N26562,N26564,N26565);
and and15822(N26563,N26566,N26567);
and and15830(N26575,N26577,N26578);
and and15831(N26576,N26579,N26580);
and and15839(N26588,N26590,N26591);
and and15840(N26589,N26592,N26593);
and and15848(N26601,N26603,N26604);
and and15849(N26602,N26605,N26606);
and and15857(N26614,N26616,N26617);
and and15858(N26615,N26618,N26619);
and and15866(N26626,N26628,N26629);
and and15867(N26627,N26630,N26631);
and and15875(N26638,N26640,N26641);
and and15876(N26639,N26642,N26643);
and and15884(N26650,N26652,N26653);
and and15885(N26651,N26654,N26655);
and and15893(N26662,N26664,N26665);
and and15894(N26663,N26666,N26667);
and and15902(N26674,N26676,N26677);
and and15903(N26675,N26678,N26679);
and and15911(N26686,N26688,N26689);
and and15912(N26687,N26690,N26691);
and and15920(N26698,N26700,N26701);
and and15921(N26699,N26702,N26703);
and and15929(N26710,N26712,N26713);
and and15930(N26711,N26714,N26715);
and and15938(N26722,N26724,N26725);
and and15939(N26723,N26726,N26727);
and and15947(N26734,N26736,N26737);
and and15948(N26735,N26738,N26739);
and and15956(N26746,N26748,N26749);
and and15957(N26747,N26750,N26751);
and and15965(N26758,N26760,N26761);
and and15966(N26759,N26762,N26763);
and and15974(N26770,N26772,N26773);
and and15975(N26771,N26774,N26775);
and and15983(N26782,N26784,N26785);
and and15984(N26783,N26786,N26787);
and and15992(N26794,N26796,N26797);
and and15993(N26795,N26798,N26799);
and and16001(N26806,N26808,N26809);
and and16002(N26807,N26810,N26811);
and and16010(N26818,N26820,N26821);
and and16011(N26819,N26822,N26823);
and and16019(N26830,N26832,N26833);
and and16020(N26831,N26834,N26835);
and and16028(N26842,N26844,N26845);
and and16029(N26843,N26846,N26847);
and and16037(N26854,N26856,N26857);
and and16038(N26855,N26858,N26859);
and and16046(N26866,N26868,N26869);
and and16047(N26867,N26870,N26871);
and and16055(N26878,N26880,N26881);
and and16056(N26879,N26882,N26883);
and and16064(N26890,N26892,N26893);
and and16065(N26891,N26894,N26895);
and and16073(N26902,N26904,N26905);
and and16074(N26903,N26906,N26907);
and and16082(N26914,N26916,N26917);
and and16083(N26915,N26918,N26919);
and and16091(N26926,N26928,N26929);
and and16092(N26927,N26930,N26931);
and and16100(N26938,N26940,N26941);
and and16101(N26939,N26942,N26943);
and and16109(N26950,N26952,N26953);
and and16110(N26951,N26954,N26955);
and and16118(N26962,N26964,N26965);
and and16119(N26963,N26966,N26967);
and and16127(N26974,N26976,N26977);
and and16128(N26975,N26978,N26979);
and and16136(N26986,N26988,N26989);
and and16137(N26987,N26990,N26991);
and and16145(N26998,N27000,N27001);
and and16146(N26999,N27002,N27003);
and and16154(N27010,N27012,N27013);
and and16155(N27011,N27014,N27015);
and and16163(N27022,N27024,N27025);
and and16164(N27023,N27026,N27027);
and and16172(N27034,N27036,N27037);
and and16173(N27035,N27038,N27039);
and and16181(N27046,N27048,N27049);
and and16182(N27047,N27050,N27051);
and and16190(N27058,N27060,N27061);
and and16191(N27059,N27062,N27063);
and and16199(N27069,N27071,N27072);
and and16200(N27070,N27073,N27074);
and and16208(N27080,N27082,N27083);
and and16209(N27081,N27084,N27085);
and and16217(N27091,N27093,N27094);
and and16218(N27092,N27095,N27096);
and and16226(N27102,N27104,N27105);
and and16227(N27103,N27106,N27107);
and and16235(N27112,N27114,N27115);
and and16236(N27113,N27116,N27117);
and and16244(N27122,N27124,N27125);
and and16245(N27123,N27126,N27127);
and and16253(N27132,N27134,N27135);
and and16254(N27133,N27136,N27137);
and and16262(N27142,N27144,N27145);
and and16263(N27143,N27146,N27147);
and and16271(N27152,N27154,N27155);
and and16272(N27153,N27156,N27157);
and and16280(N27162,N27164,N27165);
and and16281(N27163,N27166,N27167);
and and16289(N27172,N27174,N27175);
and and16290(N27173,N27176,N27177);
and and16298(N27182,N27184,N27185);
and and16299(N27183,N27186,N27187);
and and16307(N27192,N27194,N27195);
and and16308(N27193,N27196,N27197);
and and16316(N27202,N27204,N27205);
and and16317(N27203,N27206,N27207);
and and16324(N27218,N27220,N27221);
and and16325(N27219,N27222,N27223);
and and16332(N27234,N27236,N27237);
and and16333(N27235,N27238,N27239);
and and16340(N27249,N27251,N27252);
and and16341(N27250,N27253,N27254);
and and16348(N27264,N27266,N27267);
and and16349(N27265,N27268,N27269);
and and16356(N27279,N27281,N27282);
and and16357(N27280,N27283,N27284);
and and16364(N27293,N27295,N27296);
and and16365(N27294,N27297,N27298);
and and16372(N27307,N27309,N27310);
and and16373(N27308,N27311,N27312);
and and16380(N27321,N27323,N27324);
and and16381(N27322,N27325,N27326);
and and16388(N27335,N27337,N27338);
and and16389(N27336,N27339,N27340);
and and16396(N27349,N27351,N27352);
and and16397(N27350,N27353,N27354);
and and16404(N27363,N27365,N27366);
and and16405(N27364,N27367,N27368);
and and16412(N27377,N27379,N27380);
and and16413(N27378,N27381,N27382);
and and16420(N27391,N27393,N27394);
and and16421(N27392,N27395,N27396);
and and16428(N27405,N27407,N27408);
and and16429(N27406,N27409,N27410);
and and16436(N27419,N27421,N27422);
and and16437(N27420,N27423,N27424);
and and16444(N27433,N27435,N27436);
and and16445(N27434,N27437,N27438);
and and16452(N27447,N27449,N27450);
and and16453(N27448,N27451,N27452);
and and16460(N27461,N27463,N27464);
and and16461(N27462,N27465,N27466);
and and16468(N27475,N27477,N27478);
and and16469(N27476,N27479,N27480);
and and16476(N27489,N27491,N27492);
and and16477(N27490,N27493,N27494);
and and16484(N27503,N27505,N27506);
and and16485(N27504,N27507,N27508);
and and16492(N27517,N27519,N27520);
and and16493(N27518,N27521,N27522);
and and16500(N27531,N27533,N27534);
and and16501(N27532,N27535,N27536);
and and16508(N27545,N27547,N27548);
and and16509(N27546,N27549,N27550);
and and16516(N27559,N27561,N27562);
and and16517(N27560,N27563,N27564);
and and16524(N27573,N27575,N27576);
and and16525(N27574,N27577,N27578);
and and16532(N27587,N27589,N27590);
and and16533(N27588,N27591,N27592);
and and16540(N27601,N27603,N27604);
and and16541(N27602,N27605,N27606);
and and16548(N27614,N27616,N27617);
and and16549(N27615,N27618,N27619);
and and16556(N27627,N27629,N27630);
and and16557(N27628,N27631,N27632);
and and16564(N27640,N27642,N27643);
and and16565(N27641,N27644,N27645);
and and16572(N27653,N27655,N27656);
and and16573(N27654,N27657,N27658);
and and16580(N27666,N27668,N27669);
and and16581(N27667,N27670,N27671);
and and16588(N27679,N27681,N27682);
and and16589(N27680,N27683,N27684);
and and16596(N27692,N27694,N27695);
and and16597(N27693,N27696,N27697);
and and16604(N27705,N27707,N27708);
and and16605(N27706,N27709,N27710);
and and16612(N27718,N27720,N27721);
and and16613(N27719,N27722,N27723);
and and16620(N27731,N27733,N27734);
and and16621(N27732,N27735,N27736);
and and16628(N27744,N27746,N27747);
and and16629(N27745,N27748,N27749);
and and16636(N27757,N27759,N27760);
and and16637(N27758,N27761,N27762);
and and16644(N27770,N27772,N27773);
and and16645(N27771,N27774,N27775);
and and16652(N27783,N27785,N27786);
and and16653(N27784,N27787,N27788);
and and16660(N27796,N27798,N27799);
and and16661(N27797,N27800,N27801);
and and16668(N27809,N27811,N27812);
and and16669(N27810,N27813,N27814);
and and16676(N27822,N27824,N27825);
and and16677(N27823,N27826,N27827);
and and16684(N27835,N27837,N27838);
and and16685(N27836,N27839,N27840);
and and16692(N27848,N27850,N27851);
and and16693(N27849,N27852,N27853);
and and16700(N27861,N27863,N27864);
and and16701(N27862,N27865,N27866);
and and16708(N27874,N27876,N27877);
and and16709(N27875,N27878,N27879);
and and16716(N27887,N27889,N27890);
and and16717(N27888,N27891,N27892);
and and16724(N27900,N27902,N27903);
and and16725(N27901,N27904,N27905);
and and16732(N27913,N27915,N27916);
and and16733(N27914,N27917,N27918);
and and16740(N27926,N27928,N27929);
and and16741(N27927,N27930,N27931);
and and16748(N27939,N27941,N27942);
and and16749(N27940,N27943,N27944);
and and16756(N27952,N27954,N27955);
and and16757(N27953,N27956,N27957);
and and16764(N27965,N27967,N27968);
and and16765(N27966,N27969,N27970);
and and16772(N27978,N27980,N27981);
and and16773(N27979,N27982,N27983);
and and16780(N27991,N27993,N27994);
and and16781(N27992,N27995,N27996);
and and16788(N28004,N28006,N28007);
and and16789(N28005,N28008,N28009);
and and16796(N28017,N28019,N28020);
and and16797(N28018,N28021,N28022);
and and16804(N28030,N28032,N28033);
and and16805(N28031,N28034,N28035);
and and16812(N28043,N28045,N28046);
and and16813(N28044,N28047,N28048);
and and16820(N28056,N28058,N28059);
and and16821(N28057,N28060,N28061);
and and16828(N28069,N28071,N28072);
and and16829(N28070,N28073,N28074);
and and16836(N28082,N28084,N28085);
and and16837(N28083,N28086,N28087);
and and16844(N28095,N28097,N28098);
and and16845(N28096,N28099,N28100);
and and16852(N28107,N28109,N28110);
and and16853(N28108,N28111,N28112);
and and16860(N28119,N28121,N28122);
and and16861(N28120,N28123,N28124);
and and16868(N28131,N28133,N28134);
and and16869(N28132,N28135,N28136);
and and16876(N28143,N28145,N28146);
and and16877(N28144,N28147,N28148);
and and16884(N28155,N28157,N28158);
and and16885(N28156,N28159,N28160);
and and16892(N28167,N28169,N28170);
and and16893(N28168,N28171,N28172);
and and16900(N28179,N28181,N28182);
and and16901(N28180,N28183,N28184);
and and16908(N28191,N28193,N28194);
and and16909(N28192,N28195,N28196);
and and16916(N28203,N28205,N28206);
and and16917(N28204,N28207,N28208);
and and16924(N28215,N28217,N28218);
and and16925(N28216,N28219,N28220);
and and16932(N28227,N28229,N28230);
and and16933(N28228,N28231,N28232);
and and16940(N28239,N28241,N28242);
and and16941(N28240,N28243,N28244);
and and16948(N28251,N28253,N28254);
and and16949(N28252,N28255,N28256);
and and16956(N28263,N28265,N28266);
and and16957(N28264,N28267,N28268);
and and16964(N28275,N28277,N28278);
and and16965(N28276,N28279,N28280);
and and16972(N28287,N28289,N28290);
and and16973(N28288,N28291,N28292);
and and16980(N28299,N28301,N28302);
and and16981(N28300,N28303,N28304);
and and16988(N28311,N28313,N28314);
and and16989(N28312,N28315,N28316);
and and16996(N28323,N28325,N28326);
and and16997(N28324,N28327,N28328);
and and17004(N28335,N28337,N28338);
and and17005(N28336,N28339,N28340);
and and17012(N28347,N28349,N28350);
and and17013(N28348,N28351,N28352);
and and17020(N28359,N28361,N28362);
and and17021(N28360,N28363,N28364);
and and17028(N28371,N28373,N28374);
and and17029(N28372,N28375,N28376);
and and17036(N28383,N28385,N28386);
and and17037(N28384,N28387,N28388);
and and17044(N28395,N28397,N28398);
and and17045(N28396,N28399,N28400);
and and17052(N28407,N28409,N28410);
and and17053(N28408,N28411,N28412);
and and17060(N28419,N28421,N28422);
and and17061(N28420,N28423,N28424);
and and17068(N28431,N28433,N28434);
and and17069(N28432,N28435,N28436);
and and17076(N28443,N28445,N28446);
and and17077(N28444,N28447,N28448);
and and17084(N28455,N28457,N28458);
and and17085(N28456,N28459,N28460);
and and17092(N28466,N28468,N28469);
and and17093(N28467,N28470,N28471);
and and17100(N28477,N28479,N28480);
and and17101(N28478,N28481,N28482);
and and17108(N28488,N28490,N28491);
and and17109(N28489,N28492,N28493);
and and17116(N28499,N28501,N28502);
and and17117(N28500,N28503,N28504);
and and17124(N28510,N28512,N28513);
and and17125(N28511,N28514,N28515);
and and17132(N28521,N28523,N28524);
and and17133(N28522,N28525,N28526);
and and17140(N28532,N28534,N28535);
and and17141(N28533,N28536,N28537);
and and17148(N28543,N28545,N28546);
and and17149(N28544,N28547,N28548);
and and17156(N28554,N28556,N28557);
and and17157(N28555,N28558,N28559);
and and17164(N28565,N28567,N28568);
and and17165(N28566,N28569,N28570);
and and17172(N28576,N28578,N28579);
and and17173(N28577,N28580,N28581);
and and17180(N28587,N28589,N28590);
and and17181(N28588,N28591,N28592);
and and17188(N28598,N28600,N28601);
and and17189(N28599,N28602,N28603);
and and17196(N28609,N28611,N28612);
and and17197(N28610,N28613,N28614);
and and17204(N28620,N28622,N28623);
and and17205(N28621,N28624,N28625);
and and17212(N28631,N28633,N28634);
and and17213(N28632,N28635,N28636);
and and17220(N28642,N28644,N28645);
and and17221(N28643,N28646,N28647);
and and17228(N28653,N28655,N28656);
and and17229(N28654,N28657,N28658);
and and17236(N28664,N28666,N28667);
and and17237(N28665,N28668,N28669);
and and17244(N28675,N28677,N28678);
and and17245(N28676,N28679,N28680);
and and17252(N28686,N28688,N28689);
and and17253(N28687,N28690,N28691);
and and17260(N28696,N28698,N28699);
and and17261(N28697,N28700,N28701);
and and17268(N28706,N28708,N28709);
and and17269(N28707,N28710,N28711);
and and17276(N28716,N28718,N28719);
and and17277(N28717,N28720,N28721);
and and17284(N28726,N28728,N28729);
and and17285(N28727,N28730,N28731);
and and17292(N28736,N28738,N28739);
and and17293(N28737,N28740,N28741);
and and17300(N28746,N28748,N28749);
and and17301(N28747,N28750,N28751);
and and17308(N28756,N28758,N28759);
and and17309(N28757,N28760,N28761);
and and17316(N28766,N28768,N28769);
and and17317(N28767,N28770,N28771);
and and17324(N28776,N28778,N28779);
and and17325(N28777,N28780,N28781);
and and17332(N28786,N28788,N28789);
and and17333(N28787,N28790,N28791);
and and17340(N28796,N28798,N28799);
and and17341(N28797,N28800,N28801);
and and17348(N28806,N28808,N28809);
and and17349(N28807,N28810,N28811);
and and17356(N28816,N28818,N28819);
and and17357(N28817,N28820,N28821);
and and17364(N28826,N28828,N28829);
and and17365(N28827,N28830,N28831);
and and17372(N28836,N28838,N28839);
and and17373(N28837,N28840,N28841);
and and17380(N28845,N28847,N28848);
and and17381(N28846,N28849,N28850);
and and17388(N28853,N28855,N28856);
and and17389(N28854,N28857,N28858);
and and17396(N28861,N28863,N28864);
and and17397(N28862,N28865,N28866);
and and17403(N28874,N28876,N28877);
and and17404(N28875,N28878,N28879);
and and17410(N28886,N28888,N28889);
and and17411(N28887,N28890,N28891);
and and17417(N28898,N28900,N28901);
and and17418(N28899,N28902,N28903);
and and17424(N28910,N28912,N28913);
and and17425(N28911,N28914,N28915);
and and17431(N28922,N28924,N28925);
and and17432(N28923,N28926,N28927);
and and17438(N28933,N28935,N28936);
and and17439(N28934,N28937,N28938);
and and17445(N28944,N28946,N28947);
and and17446(N28945,N28948,N28949);
and and17452(N28955,N28957,N28958);
and and17453(N28956,N28959,N28960);
and and17459(N28966,N28968,N28969);
and and17460(N28967,N28970,N28971);
and and17466(N28976,N28978,N28979);
and and17467(N28977,N28980,N28981);
and and17473(N28986,N28988,N28989);
and and17474(N28987,N28990,N28991);
and and17480(N28996,N28998,N28999);
and and17481(N28997,N29000,N29001);
and and17487(N29006,N29008,N29009);
and and17488(N29007,N29010,N29011);
and and17494(N29016,N29018,N29019);
and and17495(N29017,N29020,N29021);
and and17501(N29026,N29028,N29029);
and and17502(N29027,N29030,N29031);
and and17508(N29036,N29038,N29039);
and and17509(N29037,N29040,N29041);
and and17515(N29045,N29047,N29048);
and and17516(N29046,N29049,N29050);
and and14374(N24194,N24198,N24199);
and and14375(N24195,N24200,N24201);
and and14376(N24196,N24202,R1);
and and14377(N24197,N24203,N24204);
and and14383(N24212,N24216,N24217);
and and14384(N24213,N24218,N24219);
and and14385(N24214,R0,N24220);
and and14386(N24215,N24221,N24222);
and and14392(N24230,N24234,N24235);
and and14393(N24231,N24236,N24237);
and and14394(N24232,N24238,N24239);
and and14395(N24233,N24240,N24241);
and and14401(N24248,N24252,N24253);
and and14402(N24249,N24254,N24255);
and and14403(N24250,N24256,N24257);
and and14404(N24251,N24258,N24259);
and and14410(N24266,N24270,N24271);
and and14411(N24267,N24272,in2);
and and14412(N24268,N24273,N24274);
and and14413(N24269,N24275,N24276);
and and14419(N24284,N24288,N24289);
and and14420(N24285,N24290,in1);
and and14421(N24286,N24291,N24292);
and and14422(N24287,N24293,N24294);
and and14428(N24302,N24306,N24307);
and and14429(N24303,N24308,N24309);
and and14430(N24304,N24310,N24311);
and and14431(N24305,N24312,R3);
and and14437(N24320,N24324,N24325);
and and14438(N24321,N24326,N24327);
and and14439(N24322,N24328,R1);
and and14440(N24323,N24329,N24330);
and and14446(N24337,N24341,N24342);
and and14447(N24338,N24343,N24344);
and and14448(N24339,R0,N24345);
and and14449(N24340,N24346,N24347);
and and14455(N24354,N24358,N24359);
and and14456(N24355,N24360,in1);
and and14457(N24356,in2,N24361);
and and14458(N24357,N24362,N24363);
and and14464(N24371,N24375,N24376);
and and14465(N24372,in0,N24377);
and and14466(N24373,N24378,N24379);
and and14467(N24374,R2,N24380);
and and14473(N24388,N24392,N24393);
and and14474(N24389,N24394,N24395);
and and14475(N24390,N24396,N24397);
and and14476(N24391,R2,N24398);
and and14482(N24405,N24409,N24410);
and and14483(N24406,N24411,in2);
and and14484(N24407,N24412,N24413);
and and14485(N24408,N24414,N24415);
and and14491(N24422,N24426,N24427);
and and14492(N24423,N24428,N24429);
and and14493(N24424,N24430,N24431);
and and14494(N24425,N24432,N24433);
and and14500(N24439,N24443,N24444);
and and14501(N24440,N24445,N24446);
and and14502(N24441,N24447,N24448);
and and14503(N24442,N24449,N24450);
and and14509(N24456,N24460,N24461);
and and14510(N24457,N24462,N24463);
and and14511(N24458,N24464,N24465);
and and14512(N24459,N24466,N24467);
and and14518(N24473,N24477,N24478);
and and14519(N24474,N24479,in1);
and and14520(N24475,N24480,R1);
and and14521(N24476,N24481,R3);
and and14527(N24489,N24493,N24494);
and and14528(N24490,N24495,N24496);
and and14529(N24491,in2,N24497);
and and14530(N24492,R1,R3);
and and14536(N24505,N24509,N24510);
and and14537(N24506,in0,in2);
and and14538(N24507,N24511,N24512);
and and14539(N24508,N24513,N24514);
and and14545(N24521,N24525,N24526);
and and14546(N24522,in0,in1);
and and14547(N24523,N24527,N24528);
and and14548(N24524,N24529,N24530);
and and14554(N24537,N24541,N24542);
and and14555(N24538,in0,in1);
and and14556(N24539,in2,N24543);
and and14557(N24540,N24544,N24545);
and and14563(N24553,N24557,N24558);
and and14564(N24554,N24559,in1);
and and14565(N24555,in2,N24560);
and and14566(N24556,R2,N24561);
and and14572(N24569,N24573,N24574);
and and14573(N24570,in1,in2);
and and14574(N24571,N24575,N24576);
and and14575(N24572,N24577,N24578);
and and14581(N24585,N24589,N24590);
and and14582(N24586,in0,in1);
and and14583(N24587,N24591,N24592);
and and14584(N24588,N24593,N24594);
and and14590(N24601,N24605,N24606);
and and14591(N24602,in0,in2);
and and14592(N24603,N24607,N24608);
and and14593(N24604,N24609,R3);
and and14599(N24617,N24621,N24622);
and and14600(N24618,in0,in1);
and and14601(N24619,N24623,N24624);
and and14602(N24620,N24625,R3);
and and14608(N24633,N24637,N24638);
and and14609(N24634,N24639,N24640);
and and14610(N24635,N24641,N24642);
and and14611(N24636,R2,N24643);
and and14617(N24649,N24653,N24654);
and and14618(N24650,N24655,in1);
and and14619(N24651,N24656,R0);
and and14620(N24652,R2,N24657);
and and14626(N24665,N24669,N24670);
and and14627(N24666,N24671,N24672);
and and14628(N24667,in2,N24673);
and and14629(N24668,N24674,R2);
and and14635(N24681,N24685,N24686);
and and14636(N24682,N24687,N24688);
and and14637(N24683,R0,R1);
and and14638(N24684,N24689,N24690);
and and14644(N24697,N24701,N24702);
and and14645(N24698,N24703,N24704);
and and14646(N24699,N24705,N24706);
and and14647(N24700,R2,R3);
and and14653(N24713,N24717,N24718);
and and14654(N24714,N24719,in1);
and and14655(N24715,N24720,N24721);
and and14656(N24716,R2,R3);
and and14662(N24729,N24733,N24734);
and and14663(N24730,N24735,N24736);
and and14664(N24731,N24737,R0);
and and14665(N24732,N24738,N24739);
and and14671(N24745,N24749,N24750);
and and14672(N24746,N24751,in1);
and and14673(N24747,N24752,N24753);
and and14674(N24748,N24754,R2);
and and14680(N24761,N24765,N24766);
and and14681(N24762,N24767,N24768);
and and14682(N24763,N24769,N24770);
and and14683(N24764,R1,R3);
and and14689(N24777,N24781,N24782);
and and14690(N24778,N24783,in1);
and and14691(N24779,N24784,N24785);
and and14692(N24780,N24786,N24787);
and and14698(N24793,N24797,N24798);
and and14699(N24794,N24799,N24800);
and and14700(N24795,N24801,N24802);
and and14701(N24796,R2,N24803);
and and14707(N24809,N24813,N24814);
and and14708(N24810,N24815,in1);
and and14709(N24811,R0,N24816);
and and14710(N24812,N24817,N24818);
and and14716(N24825,N24829,N24830);
and and14717(N24826,N24831,N24832);
and and14718(N24827,N24833,R0);
and and14719(N24828,N24834,N24835);
and and14725(N24841,N24845,N24846);
and and14726(N24842,N24847,N24848);
and and14727(N24843,N24849,N24850);
and and14728(N24844,R2,R3);
and and14734(N24857,N24861,N24862);
and and14735(N24858,N24863,N24864);
and and14736(N24859,R0,N24865);
and and14737(N24860,N24866,R3);
and and14743(N24873,N24877,N24878);
and and14744(N24874,N24879,N24880);
and and14745(N24875,N24881,N24882);
and and14746(N24876,R1,N24883);
and and14752(N24889,N24893,N24894);
and and14753(N24890,N24895,N24896);
and and14754(N24891,in2,N24897);
and and14755(N24892,N24898,N24899);
and and14761(N24905,N24909,N24910);
and and14762(N24906,N24911,in1);
and and14763(N24907,N24912,N24913);
and and14764(N24908,N24914,N24915);
and and14770(N24921,N24925,N24926);
and and14771(N24922,N24927,in1);
and and14772(N24923,N24928,N24929);
and and14773(N24924,N24930,N24931);
and and14779(N24937,N24941,N24942);
and and14780(N24938,N24943,N24944);
and and14781(N24939,R0,N24945);
and and14782(N24940,N24946,N24947);
and and14788(N24953,N24957,N24958);
and and14789(N24954,N24959,in2);
and and14790(N24955,R0,N24960);
and and14791(N24956,R2,R3);
and and14797(N24968,N24972,N24973);
and and14798(N24969,N24974,N24975);
and and14799(N24970,N24976,R0);
and and14800(N24971,N24977,R2);
and and14806(N24983,N24987,N24988);
and and14807(N24984,in0,N24989);
and and14808(N24985,in2,R1);
and and14809(N24986,N24990,N24991);
and and14815(N24998,N25002,N25003);
and and14816(N24999,in0,in1);
and and14817(N25000,N25004,R1);
and and14818(N25001,N25005,N25006);
and and14824(N25013,N25017,N25018);
and and14825(N25014,in0,in2);
and and14826(N25015,R0,N25019);
and and14827(N25016,N25020,N25021);
and and14833(N25028,N25032,N25033);
and and14834(N25029,in0,in1);
and and14835(N25030,N25034,R0);
and and14836(N25031,N25035,N25036);
and and14842(N25043,N25047,N25048);
and and14843(N25044,N25049,N25050);
and and14844(N25045,in2,R0);
and and14845(N25046,N25051,N25052);
and and14851(N25058,N25062,N25063);
and and14852(N25059,N25064,in2);
and and14853(N25060,N25065,N25066);
and and14854(N25061,R2,R3);
and and14860(N25073,N25077,N25078);
and and14861(N25074,N25079,N25080);
and and14862(N25075,N25081,N25082);
and and14863(N25076,N25083,R3);
and and14869(N25088,N25092,N25093);
and and14870(N25089,N25094,N25095);
and and14871(N25090,N25096,R1);
and and14872(N25091,R2,N25097);
and and14878(N25103,N25107,N25108);
and and14879(N25104,N25109,N25110);
and and14880(N25105,N25111,N25112);
and and14881(N25106,R1,R2);
and and14887(N25118,N25122,N25123);
and and14888(N25119,N25124,N25125);
and and14889(N25120,in2,N25126);
and and14890(N25121,R1,R2);
and and14896(N25133,N25137,N25138);
and and14897(N25134,in0,N25139);
and and14898(N25135,N25140,R0);
and and14899(N25136,R1,N25141);
and and14905(N25148,N25152,N25153);
and and14906(N25149,N25154,N25155);
and and14907(N25150,in2,N25156);
and and14908(N25151,R1,N25157);
and and14914(N25163,N25167,N25168);
and and14915(N25164,N25169,in1);
and and14916(N25165,N25170,N25171);
and and14917(N25166,R1,N25172);
and and14923(N25178,N25182,N25183);
and and14924(N25179,N25184,N25185);
and and14925(N25180,N25186,R1);
and and14926(N25181,R2,N25187);
and and14932(N25193,N25197,N25198);
and and14933(N25194,N25199,N25200);
and and14934(N25195,in2,N25201);
and and14935(N25196,N25202,R3);
and and14941(N25208,N25212,N25213);
and and14942(N25209,N25214,N25215);
and and14943(N25210,N25216,R0);
and and14944(N25211,N25217,N25218);
and and14950(N25223,N25227,N25228);
and and14951(N25224,N25229,N25230);
and and14952(N25225,R0,N25231);
and and14953(N25226,N25232,N25233);
and and14959(N25238,N25242,N25243);
and and14960(N25239,N25244,N25245);
and and14961(N25240,in2,R0);
and and14962(N25241,N25246,N25247);
and and14968(N25253,N25257,N25258);
and and14969(N25254,N25259,in1);
and and14970(N25255,in2,N25260);
and and14971(N25256,N25261,N25262);
and and14977(N25268,N25272,N25273);
and and14978(N25269,in0,N25274);
and and14979(N25270,N25275,R0);
and and14980(N25271,N25276,R2);
and and14986(N25283,N25287,N25288);
and and14987(N25284,N25289,N25290);
and and14988(N25285,N25291,R0);
and and14989(N25286,R1,R2);
and and14995(N25298,N25302,N25303);
and and14996(N25299,N25304,N25305);
and and14997(N25300,in2,R0);
and and14998(N25301,N25306,N25307);
and and15004(N25313,N25317,N25318);
and and15005(N25314,in1,N25319);
and and15006(N25315,R0,N25320);
and and15007(N25316,N25321,N25322);
and and15013(N25328,N25332,N25333);
and and15014(N25329,in0,in1);
and and15015(N25330,N25334,R1);
and and15016(N25331,N25335,N25336);
and and15022(N25343,N25347,N25348);
and and15023(N25344,N25349,in1);
and and15024(N25345,N25350,R0);
and and15025(N25346,N25351,N25352);
and and15031(N25358,N25362,N25363);
and and15032(N25359,N25364,N25365);
and and15033(N25360,N25366,N25367);
and and15034(N25361,N25368,R2);
and and15040(N25373,N25377,N25378);
and and15041(N25374,in0,N25379);
and and15042(N25375,N25380,R0);
and and15043(N25376,R1,N25381);
and and15049(N25388,N25392,N25393);
and and15050(N25389,N25394,N25395);
and and15051(N25390,in2,R1);
and and15052(N25391,N25396,R3);
and and15058(N25403,N25407,N25408);
and and15059(N25404,N25409,in1);
and and15060(N25405,N25410,N25411);
and and15061(N25406,R1,N25412);
and and15067(N25418,N25422,N25423);
and and15068(N25419,N25424,in1);
and and15069(N25420,N25425,N25426);
and and15070(N25421,R2,R3);
and and15076(N25432,N25436,N25437);
and and15077(N25433,N25438,in2);
and and15078(N25434,N25439,N25440);
and and15079(N25435,R2,N25441);
and and15085(N25446,N25450,N25451);
and and15086(N25447,N25452,in1);
and and15087(N25448,in2,R1);
and and15088(N25449,R2,N25453);
and and15094(N25460,N25464,N25465);
and and15095(N25461,N25466,N25467);
and and15096(N25462,in2,N25468);
and and15097(N25463,R1,R2);
and and15103(N25474,N25478,N25479);
and and15104(N25475,N25480,in1);
and and15105(N25476,N25481,N25482);
and and15106(N25477,R1,R2);
and and15112(N25488,N25492,N25493);
and and15113(N25489,N25494,in1);
and and15114(N25490,N25495,R0);
and and15115(N25491,R1,R2);
and and15121(N25502,N25506,N25507);
and and15122(N25503,N25508,N25509);
and and15123(N25504,N25510,N25511);
and and15124(N25505,R2,R3);
and and15130(N25516,N25520,N25521);
and and15131(N25517,in0,in1);
and and15132(N25518,N25522,N25523);
and and15133(N25519,N25524,N25525);
and and15139(N25530,N25534,N25535);
and and15140(N25531,N25536,in1);
and and15141(N25532,N25537,R0);
and and15142(N25533,N25538,R3);
and and15148(N25544,N25548,N25549);
and and15149(N25545,N25550,N25551);
and and15150(N25546,R0,N25552);
and and15151(N25547,R2,R3);
and and15157(N25558,N25562,N25563);
and and15158(N25559,N25564,in1);
and and15159(N25560,N25565,R1);
and and15160(N25561,R2,R3);
and and15166(N25572,N25576,N25577);
and and15167(N25573,N25578,N25579);
and and15168(N25574,N25580,R0);
and and15169(N25575,R1,N25581);
and and15175(N25586,N25590,N25591);
and and15176(N25587,N25592,in1);
and and15177(N25588,in2,N25593);
and and15178(N25589,N25594,N25595);
and and15184(N25600,N25604,N25605);
and and15185(N25601,in0,in1);
and and15186(N25602,in2,R0);
and and15187(N25603,N25606,N25607);
and and15193(N25614,N25618,N25619);
and and15194(N25615,N25620,in1);
and and15195(N25616,in2,R0);
and and15196(N25617,N25621,R2);
and and15202(N25628,N25632,N25633);
and and15203(N25629,N25634,in1);
and and15204(N25630,in2,N25635);
and and15205(N25631,R2,R3);
and and15211(N25642,N25646,N25647);
and and15212(N25643,N25648,in1);
and and15213(N25644,R0,N25649);
and and15214(N25645,R2,N25650);
and and15220(N25656,N25660,N25661);
and and15221(N25657,N25662,N25663);
and and15222(N25658,R0,R1);
and and15223(N25659,N25664,R3);
and and15229(N25670,N25674,N25675);
and and15230(N25671,N25676,N25677);
and and15231(N25672,N25678,N25679);
and and15232(N25673,N25680,R3);
and and15238(N25684,N25688,N25689);
and and15239(N25685,in0,in1);
and and15240(N25686,N25690,N25691);
and and15241(N25687,R2,N25692);
and and15247(N25698,N25702,N25703);
and and15248(N25699,in0,N25704);
and and15249(N25700,in2,N25705);
and and15250(N25701,N25706,R2);
and and15256(N25712,N25716,N25717);
and and15257(N25713,in0,in1);
and and15258(N25714,in2,R0);
and and15259(N25715,N25718,N25719);
and and15265(N25726,N25730,N25731);
and and15266(N25727,N25732,N25733);
and and15267(N25728,N25734,N25735);
and and15268(N25729,R1,R2);
and and15274(N25740,N25744,N25745);
and and15275(N25741,N25746,N25747);
and and15276(N25742,R0,R1);
and and15277(N25743,R2,R3);
and and15283(N25754,N25758,N25759);
and and15284(N25755,N25760,N25761);
and and15285(N25756,N25762,R0);
and and15286(N25757,R1,R2);
and and15292(N25768,N25772,N25773);
and and15293(N25769,in1,in2);
and and15294(N25770,R0,N25774);
and and15295(N25771,R2,N25775);
and and15301(N25782,N25786,N25787);
and and15302(N25783,N25788,N25789);
and and15303(N25784,N25790,R0);
and and15304(N25785,R1,R2);
and and15310(N25796,N25800,N25801);
and and15311(N25797,N25802,in1);
and and15312(N25798,in2,R0);
and and15313(N25799,N25803,N25804);
and and15319(N25810,N25814,N25815);
and and15320(N25811,in0,in1);
and and15321(N25812,N25816,R0);
and and15322(N25813,N25817,N25818);
and and15328(N25824,N25828,N25829);
and and15329(N25825,N25830,in1);
and and15330(N25826,in2,R0);
and and15331(N25827,N25831,N25832);
and and15337(N25838,N25842,N25843);
and and15338(N25839,N25844,in1);
and and15339(N25840,N25845,R0);
and and15340(N25841,R2,R3);
and and15346(N25852,N25856,N25857);
and and15347(N25853,N25858,N25859);
and and15348(N25854,in2,R0);
and and15349(N25855,N25860,R2);
and and15355(N25866,N25870,N25871);
and and15356(N25867,N25872,N25873);
and and15357(N25868,in2,R0);
and and15358(N25869,R1,R2);
and and15364(N25880,N25884,N25885);
and and15365(N25881,in0,in2);
and and15366(N25882,R0,N25886);
and and15367(N25883,N25887,R3);
and and15373(N25894,N25898,N25899);
and and15374(N25895,in0,in1);
and and15375(N25896,N25900,R0);
and and15376(N25897,N25901,R3);
and and15382(N25908,N25912,N25913);
and and15383(N25909,in0,in2);
and and15384(N25910,R0,N25914);
and and15385(N25911,R2,N25915);
and and15391(N25922,N25926,N25927);
and and15392(N25923,in0,in1);
and and15393(N25924,N25928,R0);
and and15394(N25925,N25929,R2);
and and15400(N25936,N25940,N25941);
and and15401(N25937,N25942,in1);
and and15402(N25938,in2,R0);
and and15403(N25939,R2,N25943);
and and15409(N25950,N25954,N25955);
and and15410(N25951,in0,N25956);
and and15411(N25952,N25957,R0);
and and15412(N25953,R1,R2);
and and15418(N25964,N25968,N25969);
and and15419(N25965,N25970,in1);
and and15420(N25966,N25971,R0);
and and15421(N25967,R1,N25972);
and and15427(N25978,N25982,N25983);
and and15428(N25979,N25984,N25985);
and and15429(N25980,in2,R0);
and and15430(N25981,R1,N25986);
and and15436(N25992,N25996,N25997);
and and15437(N25993,N25998,N25999);
and and15438(N25994,in2,N26000);
and and15439(N25995,R2,R3);
and and15445(N26006,N26010,N26011);
and and15446(N26007,N26012,in1);
and and15447(N26008,in2,R0);
and and15448(N26009,R1,N26013);
and and15454(N26020,N26024,N26025);
and and15455(N26021,N26026,in1);
and and15456(N26022,N26027,N26028);
and and15457(N26023,R1,R2);
and and15463(N26034,N26038,N26039);
and and15464(N26035,N26040,in2);
and and15465(N26036,N26041,N26042);
and and15466(N26037,R2,N26043);
and and15472(N26048,N26052,N26053);
and and15473(N26049,N26054,N26055);
and and15474(N26050,in2,R0);
and and15475(N26051,R1,N26056);
and and15481(N26062,N26066,N26067);
and and15482(N26063,N26068,N26069);
and and15483(N26064,N26070,N26071);
and and15484(N26065,R2,R3);
and and15490(N26076,N26080,N26081);
and and15491(N26077,in0,N26082);
and and15492(N26078,R0,N26083);
and and15493(N26079,N26084,R3);
and and15499(N26090,N26094,N26095);
and and15500(N26091,N26096,N26097);
and and15501(N26092,in2,R0);
and and15502(N26093,N26098,N26099);
and and15508(N26104,N26108,N26109);
and and15509(N26105,in0,N26110);
and and15510(N26106,in2,R0);
and and15511(N26107,R1,R3);
and and15517(N26118,N26122,N26123);
and and15518(N26119,N26124,in2);
and and15519(N26120,N26125,N26126);
and and15520(N26121,R2,R3);
and and15526(N26132,N26136,N26137);
and and15527(N26133,in0,N26138);
and and15528(N26134,in2,N26139);
and and15529(N26135,R2,N26140);
and and15535(N26146,N26150,N26151);
and and15536(N26147,N26152,N26153);
and and15537(N26148,R0,N26154);
and and15538(N26149,R2,N26155);
and and15544(N26160,N26164,N26165);
and and15545(N26161,N26166,N26167);
and and15546(N26162,in2,R0);
and and15547(N26163,R1,N26168);
and and15553(N26174,N26178,N26179);
and and15554(N26175,N26180,in1);
and and15555(N26176,in2,R0);
and and15556(N26177,N26181,N26182);
and and15562(N26187,N26191,N26192);
and and15563(N26188,N26193,N26194);
and and15564(N26189,in2,N26195);
and and15565(N26190,R1,R2);
and and15571(N26200,N26204,N26205);
and and15572(N26201,N26206,in2);
and and15573(N26202,R0,N26207);
and and15574(N26203,R2,R3);
and and15580(N26213,N26217,N26218);
and and15581(N26214,in1,in2);
and and15582(N26215,R0,N26219);
and and15583(N26216,R2,N26220);
and and15589(N26226,N26230,N26231);
and and15590(N26227,in0,in1);
and and15591(N26228,N26232,R0);
and and15592(N26229,R1,R2);
and and15598(N26239,N26243,N26244);
and and15599(N26240,in0,in2);
and and15600(N26241,R0,N26245);
and and15601(N26242,R2,R3);
and and15607(N26252,N26256,N26257);
and and15608(N26253,in0,in1);
and and15609(N26254,in2,N26258);
and and15610(N26255,R1,N26259);
and and15616(N26265,N26269,N26270);
and and15617(N26266,N26271,N26272);
and and15618(N26267,N26273,R1);
and and15619(N26268,R2,R3);
and and15625(N26278,N26282,N26283);
and and15626(N26279,N26284,in1);
and and15627(N26280,R0,N26285);
and and15628(N26281,N26286,R3);
and and15634(N26291,N26295,N26296);
and and15635(N26292,N26297,N26298);
and and15636(N26293,in2,R0);
and and15637(N26294,N26299,N26300);
and and15643(N26304,N26308,N26309);
and and15644(N26305,in0,in1);
and and15645(N26306,in2,R0);
and and15646(N26307,N26310,R2);
and and15652(N26317,N26321,N26322);
and and15653(N26318,N26323,in1);
and and15654(N26319,N26324,N26325);
and and15655(N26320,R2,N26326);
and and15661(N26330,N26334,N26335);
and and15662(N26331,N26336,in1);
and and15663(N26332,R0,R1);
and and15664(N26333,R2,R3);
and and15670(N26343,N26347,N26348);
and and15671(N26344,N26349,N26350);
and and15672(N26345,in2,N26351);
and and15673(N26346,N26352,R3);
and and15679(N26356,N26360,N26361);
and and15680(N26357,in1,in2);
and and15681(N26358,R0,N26362);
and and15682(N26359,N26363,N26364);
and and15688(N26369,N26373,N26374);
and and15689(N26370,in0,in1);
and and15690(N26371,N26375,R0);
and and15691(N26372,N26376,N26377);
and and15697(N26382,N26386,N26387);
and and15698(N26383,N26388,in2);
and and15699(N26384,N26389,R1);
and and15700(N26385,N26390,R3);
and and15706(N26395,N26399,N26400);
and and15707(N26396,in0,N26401);
and and15708(N26397,N26402,R1);
and and15709(N26398,R2,R3);
and and15715(N26408,N26412,N26413);
and and15716(N26409,in1,N26414);
and and15717(N26410,N26415,R1);
and and15718(N26411,R2,R3);
and and15724(N26421,N26425,N26426);
and and15725(N26422,N26427,in2);
and and15726(N26423,R0,N26428);
and and15727(N26424,R2,N26429);
and and15733(N26434,N26438,N26439);
and and15734(N26435,N26440,N26441);
and and15735(N26436,in2,N26442);
and and15736(N26437,R1,R3);
and and15742(N26447,N26451,N26452);
and and15743(N26448,N26453,N26454);
and and15744(N26449,R0,R1);
and and15745(N26450,R2,R3);
and and15751(N26460,N26464,N26465);
and and15752(N26461,in0,in1);
and and15753(N26462,in2,R0);
and and15754(N26463,N26466,N26467);
and and15760(N26473,N26477,N26478);
and and15761(N26474,in0,in1);
and and15762(N26475,N26479,N26480);
and and15763(N26476,N26481,R3);
and and15769(N26486,N26490,N26491);
and and15770(N26487,N26492,in1);
and and15771(N26488,N26493,R0);
and and15772(N26489,N26494,R3);
and and15778(N26499,N26503,N26504);
and and15779(N26500,N26505,in1);
and and15780(N26501,in2,N26506);
and and15781(N26502,R1,R2);
and and15787(N26512,N26516,N26517);
and and15788(N26513,in0,in1);
and and15789(N26514,N26518,N26519);
and and15790(N26515,N26520,R2);
and and15796(N26525,N26529,N26530);
and and15797(N26526,in0,in1);
and and15798(N26527,N26531,R0);
and and15799(N26528,R1,N26532);
and and15805(N26538,N26542,N26543);
and and15806(N26539,N26544,in1);
and and15807(N26540,in2,R0);
and and15808(N26541,N26545,R3);
and and15814(N26551,N26555,N26556);
and and15815(N26552,in0,in1);
and and15816(N26553,in2,R0);
and and15817(N26554,R1,N26557);
and and15823(N26564,N26568,N26569);
and and15824(N26565,in0,in1);
and and15825(N26566,N26570,N26571);
and and15826(N26567,N26572,R2);
and and15832(N26577,N26581,N26582);
and and15833(N26578,N26583,in1);
and and15834(N26579,in2,N26584);
and and15835(N26580,R2,R3);
and and15841(N26590,N26594,N26595);
and and15842(N26591,N26596,in1);
and and15843(N26592,in2,R0);
and and15844(N26593,N26597,R3);
and and15850(N26603,N26607,N26608);
and and15851(N26604,N26609,N26610);
and and15852(N26605,in2,R0);
and and15853(N26606,R1,N26611);
and and15859(N26616,N26620,N26621);
and and15860(N26617,N26622,in1);
and and15861(N26618,in2,R0);
and and15862(N26619,R2,R3);
and and15868(N26628,N26632,N26633);
and and15869(N26629,N26634,in1);
and and15870(N26630,in2,R0);
and and15871(N26631,R1,R2);
and and15877(N26640,N26644,N26645);
and and15878(N26641,N26646,in2);
and and15879(N26642,N26647,R1);
and and15880(N26643,R2,R3);
and and15886(N26652,N26656,N26657);
and and15887(N26653,in0,in2);
and and15888(N26654,N26658,R1);
and and15889(N26655,R2,R3);
and and15895(N26664,N26668,N26669);
and and15896(N26665,N26670,in1);
and and15897(N26666,in2,N26671);
and and15898(N26667,R2,R3);
and and15904(N26676,N26680,N26681);
and and15905(N26677,in0,in1);
and and15906(N26678,N26682,R1);
and and15907(N26679,R2,R3);
and and15913(N26688,N26692,N26693);
and and15914(N26689,N26694,in1);
and and15915(N26690,R0,R1);
and and15916(N26691,R2,N26695);
and and15922(N26700,N26704,N26705);
and and15923(N26701,N26706,in1);
and and15924(N26702,N26707,R0);
and and15925(N26703,R2,R3);
and and15931(N26712,N26716,N26717);
and and15932(N26713,in1,in2);
and and15933(N26714,R0,R1);
and and15934(N26715,N26718,R3);
and and15940(N26724,N26728,N26729);
and and15941(N26725,N26730,in1);
and and15942(N26726,N26731,R1);
and and15943(N26727,R2,R3);
and and15949(N26736,N26740,N26741);
and and15950(N26737,in0,in1);
and and15951(N26738,in2,R0);
and and15952(N26739,N26742,R2);
and and15958(N26748,N26752,N26753);
and and15959(N26749,in0,N26754);
and and15960(N26750,in2,R0);
and and15961(N26751,R1,R2);
and and15967(N26760,N26764,N26765);
and and15968(N26761,N26766,N26767);
and and15969(N26762,in2,N26768);
and and15970(N26763,R1,R2);
and and15976(N26772,N26776,N26777);
and and15977(N26773,in1,in2);
and and15978(N26774,N26778,R1);
and and15979(N26775,R2,N26779);
and and15985(N26784,N26788,N26789);
and and15986(N26785,in0,N26790);
and and15987(N26786,in2,R1);
and and15988(N26787,R2,N26791);
and and15994(N26796,N26800,N26801);
and and15995(N26797,in0,in1);
and and15996(N26798,N26802,R1);
and and15997(N26799,N26803,R3);
and and16003(N26808,N26812,N26813);
and and16004(N26809,N26814,in1);
and and16005(N26810,in2,R0);
and and16006(N26811,R1,R2);
and and16012(N26820,N26824,N26825);
and and16013(N26821,N26826,in1);
and and16014(N26822,in2,N26827);
and and16015(N26823,R1,R2);
and and16021(N26832,N26836,N26837);
and and16022(N26833,in0,in1);
and and16023(N26834,N26838,R0);
and and16024(N26835,R1,R2);
and and16030(N26844,N26848,N26849);
and and16031(N26845,in0,in1);
and and16032(N26846,N26850,R0);
and and16033(N26847,R2,N26851);
and and16039(N26856,N26860,N26861);
and and16040(N26857,N26862,in1);
and and16041(N26858,in2,R0);
and and16042(N26859,R1,R2);
and and16048(N26868,N26872,N26873);
and and16049(N26869,in1,in2);
and and16050(N26870,R0,N26874);
and and16051(N26871,R2,R3);
and and16057(N26880,N26884,N26885);
and and16058(N26881,in0,in2);
and and16059(N26882,R0,N26886);
and and16060(N26883,N26887,N26888);
and and16066(N26892,N26896,N26897);
and and16067(N26893,in0,N26898);
and and16068(N26894,R0,R1);
and and16069(N26895,R2,R3);
and and16075(N26904,N26908,N26909);
and and16076(N26905,N26910,N26911);
and and16077(N26906,R0,R1);
and and16078(N26907,R2,R3);
and and16084(N26916,N26920,N26921);
and and16085(N26917,in0,in1);
and and16086(N26918,in2,R0);
and and16087(N26919,R1,R2);
and and16093(N26928,N26932,N26933);
and and16094(N26929,in0,N26934);
and and16095(N26930,R0,R1);
and and16096(N26931,R2,N26935);
and and16102(N26940,N26944,N26945);
and and16103(N26941,N26946,in2);
and and16104(N26942,R0,R1);
and and16105(N26943,R2,N26947);
and and16111(N26952,N26956,N26957);
and and16112(N26953,in1,N26958);
and and16113(N26954,R0,R1);
and and16114(N26955,R2,N26959);
and and16120(N26964,N26968,N26969);
and and16121(N26965,in0,N26970);
and and16122(N26966,N26971,R0);
and and16123(N26967,R1,R2);
and and16129(N26976,N26980,N26981);
and and16130(N26977,N26982,in1);
and and16131(N26978,in2,R0);
and and16132(N26979,N26983,N26984);
and and16138(N26988,N26992,N26993);
and and16139(N26989,in0,in1);
and and16140(N26990,in2,N26994);
and and16141(N26991,N26995,R2);
and and16147(N27000,N27004,N27005);
and and16148(N27001,in0,in2);
and and16149(N27002,R0,N27006);
and and16150(N27003,R2,N27007);
and and16156(N27012,N27016,N27017);
and and16157(N27013,in0,in1);
and and16158(N27014,N27018,R0);
and and16159(N27015,N27019,R2);
and and16165(N27024,N27028,N27029);
and and16166(N27025,in0,in1);
and and16167(N27026,in2,N27030);
and and16168(N27027,R2,R3);
and and16174(N27036,N27040,N27041);
and and16175(N27037,in0,N27042);
and and16176(N27038,R0,R1);
and and16177(N27039,R2,R3);
and and16183(N27048,N27052,N27053);
and and16184(N27049,in1,N27054);
and and16185(N27050,R0,R1);
and and16186(N27051,R2,R3);
and and16192(N27060,N27064,N27065);
and and16193(N27061,N27066,in1);
and and16194(N27062,in2,N27067);
and and16195(N27063,R1,R3);
and and16201(N27071,N27075,N27076);
and and16202(N27072,N27077,in2);
and and16203(N27073,R0,R1);
and and16204(N27074,R2,R3);
and and16210(N27082,N27086,N27087);
and and16211(N27083,N27088,N27089);
and and16212(N27084,R0,R1);
and and16213(N27085,R2,R3);
and and16219(N27093,N27097,N27098);
and and16220(N27094,in0,in1);
and and16221(N27095,in2,R0);
and and16222(N27096,R2,N27099);
and and16228(N27104,N27108,N27109);
and and16229(N27105,in0,in1);
and and16230(N27106,in2,R0);
and and16231(N27107,N27110,R2);
and and16237(N27114,N27118,N27119);
and and16238(N27115,in0,in2);
and and16239(N27116,R0,R1);
and and16240(N27117,R2,R3);
and and16246(N27124,N27128,N27129);
and and16247(N27125,N27130,in1);
and and16248(N27126,in2,R0);
and and16249(N27127,R1,R2);
and and16255(N27134,N27138,N27139);
and and16256(N27135,in0,in1);
and and16257(N27136,in2,R0);
and and16258(N27137,R1,N27140);
and and16264(N27144,N27148,N27149);
and and16265(N27145,in0,in1);
and and16266(N27146,in2,R0);
and and16267(N27147,R1,R2);
and and16273(N27154,N27158,N27159);
and and16274(N27155,in0,N27160);
and and16275(N27156,in2,R0);
and and16276(N27157,R1,R2);
and and16282(N27164,N27168,N27169);
and and16283(N27165,N27170,in1);
and and16284(N27166,in2,R0);
and and16285(N27167,R1,R2);
and and16291(N27174,N27178,N27179);
and and16292(N27175,in0,in1);
and and16293(N27176,in2,R0);
and and16294(N27177,R1,R2);
and and16300(N27184,N27188,N27189);
and and16301(N27185,in0,in1);
and and16302(N27186,in2,R0);
and and16303(N27187,R1,R2);
and and16309(N27194,N27198,N27199);
and and16310(N27195,in0,in1);
and and16311(N27196,in2,R0);
and and16312(N27197,R1,R2);
and and16318(N27204,N27208,in0);
and and16319(N27205,N27209,N27210);
and and16320(N27206,N27211,N27212);
and and16321(N27207,N27213,N27214);
and and16326(N27220,N27224,N27225);
and and16327(N27221,N27226,N27227);
and and16328(N27222,N27228,N27229);
and and16329(N27223,N27230,R5);
and and16334(N27236,N27240,N27241);
and and16335(N27237,N27242,N27243);
and and16336(N27238,R0,N27244);
and and16337(N27239,R3,N27245);
and and16342(N27251,N27255,N27256);
and and16343(N27252,N27257,N27258);
and and16344(N27253,R1,N27259);
and and16345(N27254,N27260,R5);
and and16350(N27266,N27270,N27271);
and and16351(N27267,N27272,N27273);
and and16352(N27268,N27274,N27275);
and and16353(N27269,R3,N27276);
and and16358(N27281,N27285,in0);
and and16359(N27282,in1,N27286);
and and16360(N27283,N27287,N27288);
and and16361(N27284,R2,N27289);
and and16366(N27295,N27299,in0);
and and16367(N27296,R0,N27300);
and and16368(N27297,N27301,N27302);
and and16369(N27298,R4,N27303);
and and16374(N27309,N27313,in0);
and and16375(N27310,N27314,N27315);
and and16376(N27311,N27316,R2);
and and16377(N27312,N27317,N27318);
and and16382(N27323,N27327,in0);
and and16383(N27324,N27328,R0);
and and16384(N27325,N27329,N27330);
and and16385(N27326,N27331,N27332);
and and16390(N27337,N27341,in0);
and and16391(N27338,N27342,R1);
and and16392(N27339,R2,N27343);
and and16393(N27340,N27344,N27345);
and and16398(N27351,N27355,in1);
and and16399(N27352,N27356,R1);
and and16400(N27353,R2,N27357);
and and16401(N27354,N27358,N27359);
and and16406(N27365,N27369,N27370);
and and16407(N27366,in1,N27371);
and and16408(N27367,N27372,N27373);
and and16409(N27368,R2,N27374);
and and16414(N27379,N27383,N27384);
and and16415(N27380,in1,R0);
and and16416(N27381,N27385,N27386);
and and16417(N27382,R3,N27387);
and and16422(N27393,N27397,N27398);
and and16423(N27394,in2,N27399);
and and16424(N27395,N27400,R2);
and and16425(N27396,N27401,N27402);
and and16430(N27407,N27411,in0);
and and16431(N27408,N27412,R0);
and and16432(N27409,N27413,N27414);
and and16433(N27410,N27415,N27416);
and and16438(N27421,N27425,N27426);
and and16439(N27422,in1,N27427);
and and16440(N27423,N27428,N27429);
and and16441(N27424,R3,R4);
and and16446(N27435,N27439,in0);
and and16447(N27436,N27440,N27441);
and and16448(N27437,N27442,N27443);
and and16449(N27438,N27444,R4);
and and16454(N27449,N27453,in0);
and and16455(N27450,N27454,N27455);
and and16456(N27451,R1,N27456);
and and16457(N27452,N27457,R5);
and and16462(N27463,N27467,N27468);
and and16463(N27464,N27469,R0);
and and16464(N27465,N27470,N27471);
and and16465(N27466,R4,R5);
and and16470(N27477,N27481,in0);
and and16471(N27478,N27482,N27483);
and and16472(N27479,N27484,N27485);
and and16473(N27480,R3,N27486);
and and16478(N27491,N27495,N27496);
and and16479(N27492,N27497,N27498);
and and16480(N27493,R2,N27499);
and and16481(N27494,R4,N27500);
and and16486(N27505,N27509,in0);
and and16487(N27506,N27510,N27511);
and and16488(N27507,R2,N27512);
and and16489(N27508,R4,N27513);
and and16494(N27519,N27523,N27524);
and and16495(N27520,N27525,in2);
and and16496(N27521,N27526,R2);
and and16497(N27522,N27527,R4);
and and16502(N27533,N27537,in1);
and and16503(N27534,N27538,N27539);
and and16504(N27535,R2,N27540);
and and16505(N27536,R4,N27541);
and and16510(N27547,N27551,N27552);
and and16511(N27548,N27553,N27554);
and and16512(N27549,R0,R2);
and and16513(N27550,N27555,N27556);
and and16518(N27561,N27565,N27566);
and and16519(N27562,N27567,N27568);
and and16520(N27563,R1,R3);
and and16521(N27564,N27569,N27570);
and and16526(N27575,N27579,in0);
and and16527(N27576,N27580,N27581);
and and16528(N27577,N27582,R3);
and and16529(N27578,N27583,R5);
and and16534(N27589,N27593,N27594);
and and16535(N27590,N27595,in2);
and and16536(N27591,N27596,N27597);
and and16537(N27592,R3,R5);
and and16542(N27603,N27607,in1);
and and16543(N27604,in2,R1);
and and16544(N27605,N27608,N27609);
and and16545(N27606,N27610,N27611);
and and16550(N27616,N27620,in0);
and and16551(N27617,N27621,R1);
and and16552(N27618,R2,R3);
and and16553(N27619,N27622,N27623);
and and16558(N27629,N27633,N27634);
and and16559(N27630,R0,N27635);
and and16560(N27631,R2,R3);
and and16561(N27632,N27636,N27637);
and and16566(N27642,N27646,in1);
and and16567(N27643,N27647,N27648);
and and16568(N27644,R1,N27649);
and and16569(N27645,R3,N27650);
and and16574(N27655,N27659,N27660);
and and16575(N27656,in1,N27661);
and and16576(N27657,N27662,N27663);
and and16577(N27658,R4,R5);
and and16582(N27668,N27672,N27673);
and and16583(N27669,in2,R0);
and and16584(N27670,R1,N27674);
and and16585(N27671,R4,N27675);
and and16590(N27681,N27685,in0);
and and16591(N27682,N27686,R0);
and and16592(N27683,N27687,R2);
and and16593(N27684,N27688,N27689);
and and16598(N27694,N27698,N27699);
and and16599(N27695,N27700,in2);
and and16600(N27696,R0,R2);
and and16601(N27697,N27701,R5);
and and16606(N27707,N27711,N27712);
and and16607(N27708,in1,N27713);
and and16608(N27709,R0,N27714);
and and16609(N27710,N27715,N27716);
and and16614(N27720,N27724,in0);
and and16615(N27721,in1,N27725);
and and16616(N27722,N27726,N27727);
and and16617(N27723,R4,R5);
and and16622(N27733,N27737,N27738);
and and16623(N27734,in2,R0);
and and16624(N27735,N27739,N27740);
and and16625(N27736,R3,R4);
and and16630(N27746,N27750,in0);
and and16631(N27747,N27751,R0);
and and16632(N27748,N27752,N27753);
and and16633(N27749,N27754,N27755);
and and16638(N27759,N27763,in0);
and and16639(N27760,N27764,N27765);
and and16640(N27761,N27766,R3);
and and16641(N27762,R4,N27767);
and and16646(N27772,N27776,N27777);
and and16647(N27773,in1,in2);
and and16648(N27774,N27778,R1);
and and16649(N27775,N27779,N27780);
and and16654(N27785,N27789,N27790);
and and16655(N27786,in1,N27791);
and and16656(N27787,R0,R1);
and and16657(N27788,N27792,N27793);
and and16662(N27798,N27802,N27803);
and and16663(N27799,N27804,R0);
and and16664(N27800,R1,N27805);
and and16665(N27801,N27806,R5);
and and16670(N27811,N27815,in1);
and and16671(N27812,in2,N27816);
and and16672(N27813,N27817,R3);
and and16673(N27814,N27818,N27819);
and and16678(N27824,N27828,in0);
and and16679(N27825,in1,N27829);
and and16680(N27826,N27830,N27831);
and and16681(N27827,R3,N27832);
and and16686(N27837,N27841,N27842);
and and16687(N27838,in1,in2);
and and16688(N27839,N27843,N27844);
and and16689(N27840,R2,R4);
and and16694(N27850,N27854,N27855);
and and16695(N27851,in2,R0);
and and16696(N27852,R2,N27856);
and and16697(N27853,N27857,N27858);
and and16702(N27863,N27867,N27868);
and and16703(N27864,N27869,R0);
and and16704(N27865,N27870,R2);
and and16705(N27866,R4,N27871);
and and16710(N27876,N27880,N27881);
and and16711(N27877,N27882,R0);
and and16712(N27878,N27883,N27884);
and and16713(N27879,R3,N27885);
and and16718(N27889,N27893,N27894);
and and16719(N27890,N27895,in2);
and and16720(N27891,R0,N27896);
and and16721(N27892,R3,N27897);
and and16726(N27902,N27906,N27907);
and and16727(N27903,in1,R0);
and and16728(N27904,R1,R3);
and and16729(N27905,N27908,N27909);
and and16734(N27915,N27919,in0);
and and16735(N27916,N27920,N27921);
and and16736(N27917,N27922,R2);
and and16737(N27918,N27923,R4);
and and16742(N27928,N27932,N27933);
and and16743(N27929,in1,N27934);
and and16744(N27930,N27935,R2);
and and16745(N27931,R4,N27936);
and and16750(N27941,N27945,in0);
and and16751(N27942,in2,N27946);
and and16752(N27943,N27947,R2);
and and16753(N27944,N27948,N27949);
and and16758(N27954,N27958,in0);
and and16759(N27955,in2,R0);
and and16760(N27956,N27959,N27960);
and and16761(N27957,N27961,N27962);
and and16766(N27967,N27971,in1);
and and16767(N27968,R0,R1);
and and16768(N27969,N27972,N27973);
and and16769(N27970,R4,N27974);
and and16774(N27980,N27984,in0);
and and16775(N27981,N27985,R0);
and and16776(N27982,N27986,R2);
and and16777(N27983,N27987,N27988);
and and16782(N27993,N27997,in0);
and and16783(N27994,in2,N27998);
and and16784(N27995,N27999,R2);
and and16785(N27996,N28000,R5);
and and16790(N28006,N28010,in0);
and and16791(N28007,N28011,R0);
and and16792(N28008,N28012,R2);
and and16793(N28009,N28013,R5);
and and16798(N28019,N28023,in1);
and and16799(N28020,N28024,N28025);
and and16800(N28021,R1,R3);
and and16801(N28022,N28026,R5);
and and16806(N28032,N28036,N28037);
and and16807(N28033,N28038,in2);
and and16808(N28034,N28039,R2);
and and16809(N28035,N28040,R4);
and and16814(N28045,N28049,N28050);
and and16815(N28046,N28051,in2);
and and16816(N28047,N28052,R2);
and and16817(N28048,R4,N28053);
and and16822(N28058,N28062,in0);
and and16823(N28059,in2,N28063);
and and16824(N28060,N28064,N28065);
and and16825(N28061,R3,N28066);
and and16830(N28071,N28075,in0);
and and16831(N28072,in2,N28076);
and and16832(N28073,R2,N28077);
and and16833(N28074,R4,N28078);
and and16838(N28084,N28088,in1);
and and16839(N28085,N28089,R0);
and and16840(N28086,R1,R3);
and and16841(N28087,N28090,N28091);
and and16846(N28097,N28101,N28102);
and and16847(N28098,N28103,R0);
and and16848(N28099,N28104,R2);
and and16849(N28100,R3,R4);
and and16854(N28109,N28113,N28114);
and and16855(N28110,in1,R1);
and and16856(N28111,R2,N28115);
and and16857(N28112,R4,R5);
and and16862(N28121,N28125,in0);
and and16863(N28122,R0,N28126);
and and16864(N28123,N28127,R3);
and and16865(N28124,R4,R5);
and and16870(N28133,N28137,N28138);
and and16871(N28134,in1,in2);
and and16872(N28135,N28139,R3);
and and16873(N28136,R4,N28140);
and and16878(N28145,N28149,in1);
and and16879(N28146,N28150,R1);
and and16880(N28147,R2,N28151);
and and16881(N28148,N28152,R5);
and and16886(N28157,N28161,in0);
and and16887(N28158,N28162,R1);
and and16888(N28159,R2,N28163);
and and16889(N28160,N28164,R5);
and and16894(N28169,N28173,in0);
and and16895(N28170,N28174,N28175);
and and16896(N28171,R1,N28176);
and and16897(N28172,R3,N28177);
and and16902(N28181,N28185,N28186);
and and16903(N28182,N28187,R0);
and and16904(N28183,N28188,R2);
and and16905(N28184,R3,R4);
and and16910(N28193,N28197,N28198);
and and16911(N28194,N28199,in2);
and and16912(N28195,R1,R3);
and and16913(N28196,R4,R5);
and and16918(N28205,N28209,N28210);
and and16919(N28206,N28211,in2);
and and16920(N28207,R0,R1);
and and16921(N28208,N28212,R4);
and and16926(N28217,N28221,in0);
and and16927(N28218,N28222,R0);
and and16928(N28219,N28223,N28224);
and and16929(N28220,R4,R5);
and and16934(N28229,N28233,N28234);
and and16935(N28230,R0,N28235);
and and16936(N28231,N28236,N28237);
and and16937(N28232,R4,R5);
and and16942(N28241,N28245,in0);
and and16943(N28242,R0,R1);
and and16944(N28243,R2,N28246);
and and16945(N28244,N28247,R5);
and and16950(N28253,N28257,in0);
and and16951(N28254,in2,N28258);
and and16952(N28255,R2,R3);
and and16953(N28256,R4,N28259);
and and16958(N28265,N28269,in0);
and and16959(N28266,in1,N28270);
and and16960(N28267,R2,R3);
and and16961(N28268,R4,N28271);
and and16966(N28277,N28281,in0);
and and16967(N28278,N28282,N28283);
and and16968(N28279,R1,R2);
and and16969(N28280,R3,N28284);
and and16974(N28289,N28293,N28294);
and and16975(N28290,N28295,R0);
and and16976(N28291,R1,N28296);
and and16977(N28292,R3,N28297);
and and16982(N28301,N28305,in0);
and and16983(N28302,R0,R1);
and and16984(N28303,N28306,N28307);
and and16985(N28304,R4,R5);
and and16990(N28313,N28317,in0);
and and16991(N28314,N28318,N28319);
and and16992(N28315,N28320,R3);
and and16993(N28316,R4,R5);
and and16998(N28325,N28329,N28330);
and and16999(N28326,N28331,N28332);
and and17000(N28327,R1,R2);
and and17001(N28328,N28333,R4);
and and17006(N28337,N28341,in0);
and and17007(N28338,N28342,N28343);
and and17008(N28339,R2,N28344);
and and17009(N28340,N28345,R5);
and and17014(N28349,N28353,in0);
and and17015(N28350,R0,R1);
and and17016(N28351,N28354,R3);
and and17017(N28352,N28355,N28356);
and and17022(N28361,N28365,in0);
and and17023(N28362,in1,R0);
and and17024(N28363,N28366,N28367);
and and17025(N28364,R3,N28368);
and and17030(N28373,N28377,in0);
and and17031(N28374,N28378,N28379);
and and17032(N28375,R2,R3);
and and17033(N28376,N28380,N28381);
and and17038(N28385,N28389,in0);
and and17039(N28386,N28390,R1);
and and17040(N28387,N28391,R3);
and and17041(N28388,R4,N28392);
and and17046(N28397,N28401,in0);
and and17047(N28398,in1,N28402);
and and17048(N28399,N28403,R2);
and and17049(N28400,N28404,R4);
and and17054(N28409,N28413,in0);
and and17055(N28410,N28414,N28415);
and and17056(N28411,N28416,R2);
and and17057(N28412,R3,N28417);
and and17062(N28421,N28425,in0);
and and17063(N28422,R0,R1);
and and17064(N28423,N28426,R3);
and and17065(N28424,N28427,R5);
and and17070(N28433,N28437,in0);
and and17071(N28434,N28438,N28439);
and and17072(N28435,R0,N28440);
and and17073(N28436,R2,N28441);
and and17078(N28445,N28449,N28450);
and and17079(N28446,in1,N28451);
and and17080(N28447,N28452,R3);
and and17081(N28448,R4,R5);
and and17086(N28457,N28461,in0);
and and17087(N28458,in2,R0);
and and17088(N28459,R1,R2);
and and17089(N28460,N28462,N28463);
and and17094(N28468,N28472,in0);
and and17095(N28469,N28473,R0);
and and17096(N28470,R1,R3);
and and17097(N28471,R4,N28474);
and and17102(N28479,N28483,N28484);
and and17103(N28480,in1,N28485);
and and17104(N28481,R0,R2);
and and17105(N28482,R3,R4);
and and17110(N28490,N28494,in0);
and and17111(N28491,N28495,N28496);
and and17112(N28492,R1,R2);
and and17113(N28493,R4,N28497);
and and17118(N28501,N28505,in0);
and and17119(N28502,R0,R1);
and and17120(N28503,R2,N28506);
and and17121(N28504,R4,N28507);
and and17126(N28512,N28516,in0);
and and17127(N28513,R0,R1);
and and17128(N28514,R2,R3);
and and17129(N28515,R4,N28517);
and and17134(N28523,N28527,N28528);
and and17135(N28524,in1,N28529);
and and17136(N28525,R0,R1);
and and17137(N28526,R2,R3);
and and17142(N28534,N28538,in1);
and and17143(N28535,in2,N28539);
and and17144(N28536,R1,R3);
and and17145(N28537,R4,R5);
and and17150(N28545,N28549,in1);
and and17151(N28546,in2,R0);
and and17152(N28547,R1,N28550);
and and17153(N28548,R4,N28551);
and and17158(N28556,N28560,in1);
and and17159(N28557,in2,N28561);
and and17160(N28558,N28562,R3);
and and17161(N28559,R4,R5);
and and17166(N28567,N28571,N28572);
and and17167(N28568,in1,N28573);
and and17168(N28569,R1,R2);
and and17169(N28570,R4,R5);
and and17174(N28578,N28582,N28583);
and and17175(N28579,in1,N28584);
and and17176(N28580,N28585,R2);
and and17177(N28581,R3,R5);
and and17182(N28589,N28593,in0);
and and17183(N28590,in2,R0);
and and17184(N28591,R1,N28594);
and and17185(N28592,N28595,R5);
and and17190(N28600,N28604,in0);
and and17191(N28601,N28605,R0);
and and17192(N28602,R1,R2);
and and17193(N28603,N28606,R4);
and and17198(N28611,N28615,in0);
and and17199(N28612,N28616,R0);
and and17200(N28613,R1,R3);
and and17201(N28614,R4,N28617);
and and17206(N28622,N28626,in0);
and and17207(N28623,N28627,R0);
and and17208(N28624,N28628,R2);
and and17209(N28625,R3,R4);
and and17214(N28633,N28637,in0);
and and17215(N28634,N28638,R0);
and and17216(N28635,N28639,R2);
and and17217(N28636,R3,R4);
and and17222(N28644,N28648,in0);
and and17223(N28645,in2,R0);
and and17224(N28646,N28649,N28650);
and and17225(N28647,R4,R5);
and and17230(N28655,N28659,in0);
and and17231(N28656,in2,N28660);
and and17232(N28657,R1,R2);
and and17233(N28658,R3,N28661);
and and17238(N28666,N28670,in0);
and and17239(N28667,in2,N28671);
and and17240(N28668,R2,N28672);
and and17241(N28669,N28673,R5);
and and17246(N28677,N28681,N28682);
and and17247(N28678,in2,R0);
and and17248(N28679,R1,R2);
and and17249(N28680,N28683,R4);
and and17254(N28688,N28692,in1);
and and17255(N28689,N28693,R0);
and and17256(N28690,N28694,R2);
and and17257(N28691,R3,R4);
and and17262(N28698,N28702,in0);
and and17263(N28699,in2,R0);
and and17264(N28700,N28703,R2);
and and17265(N28701,N28704,R4);
and and17270(N28708,N28712,in0);
and and17271(N28709,in1,R0);
and and17272(N28710,N28713,R2);
and and17273(N28711,N28714,R4);
and and17278(N28718,N28722,in0);
and and17279(N28719,N28723,R0);
and and17280(N28720,R1,R2);
and and17281(N28721,R3,N28724);
and and17286(N28728,N28732,in0);
and and17287(N28729,R0,N28733);
and and17288(N28730,N28734,R3);
and and17289(N28731,R4,R5);
and and17294(N28738,N28742,in0);
and and17295(N28739,R0,N28743);
and and17296(N28740,R2,R3);
and and17297(N28741,N28744,R5);
and and17302(N28748,N28752,in0);
and and17303(N28749,R0,R1);
and and17304(N28750,N28753,R3);
and and17305(N28751,R4,N28754);
and and17310(N28758,N28762,in1);
and and17311(N28759,in2,R0);
and and17312(N28760,N28763,R2);
and and17313(N28761,R3,R4);
and and17318(N28768,N28772,in0);
and and17319(N28769,N28773,R0);
and and17320(N28770,R1,N28774);
and and17321(N28771,R3,R5);
and and17326(N28778,N28782,in1);
and and17327(N28779,N28783,R0);
and and17328(N28780,R1,N28784);
and and17329(N28781,R3,R5);
and and17334(N28788,N28792,in0);
and and17335(N28789,N28793,R1);
and and17336(N28790,R2,N28794);
and and17337(N28791,R4,R5);
and and17342(N28798,N28802,in1);
and and17343(N28799,N28803,R0);
and and17344(N28800,R1,N28804);
and and17345(N28801,R3,R4);
and and17350(N28808,N28812,in0);
and and17351(N28809,N28813,R0);
and and17352(N28810,R1,N28814);
and and17353(N28811,R3,R4);
and and17358(N28818,N28822,in0);
and and17359(N28819,in2,R0);
and and17360(N28820,R1,R2);
and and17361(N28821,R3,N28823);
and and17366(N28828,N28832,in0);
and and17367(N28829,in1,in2);
and and17368(N28830,N28833,R1);
and and17369(N28831,R2,R3);
and and17374(N28838,N28842,in0);
and and17375(N28839,N28843,R0);
and and17376(N28840,R2,R3);
and and17377(N28841,R4,R5);
and and17382(N28847,N28851,in1);
and and17383(N28848,in2,R0);
and and17384(N28849,R1,R2);
and and17385(N28850,R3,R5);
and and17390(N28855,N28859,in0);
and and17391(N28856,in1,in2);
and and17392(N28857,R0,R1);
and and17393(N28858,R3,R5);
and and17398(N28863,N28867,R0);
and and17399(N28864,R1,N28868);
and and17400(N28865,N28869,N28870);
and and17401(N28866,N28871,N28872);
and and17405(N28876,in0,in2);
and and17406(N28877,R1,N28880);
and and17407(N28878,N28881,N28882);
and and17408(N28879,N28883,N28884);
and and17412(N28888,in0,N28892);
and and17413(N28889,R0,N28893);
and and17414(N28890,N28894,R3);
and and17415(N28891,N28895,N28896);
and and17419(N28900,in0,N28904);
and and17420(N28901,N28905,R2);
and and17421(N28902,N28906,R5);
and and17422(N28903,N28907,N28908);
and and17426(N28912,in0,N28916);
and and17427(N28913,N28917,R3);
and and17428(N28914,N28918,N28919);
and and17429(N28915,R6,N28920);
and and17433(N28924,in0,R1);
and and17434(N28925,N28928,R3);
and and17435(N28926,N28929,N28930);
and and17436(N28927,R6,N28931);
and and17440(N28935,in0,N28939);
and and17441(N28936,N28940,R2);
and and17442(N28937,N28941,R4);
and and17443(N28938,R6,N28942);
and and17447(N28946,in0,R0);
and and17448(N28947,R2,N28950);
and and17449(N28948,N28951,N28952);
and and17450(N28949,R6,N28953);
and and17454(N28957,in0,N28961);
and and17455(N28958,R1,R3);
and and17456(N28959,N28962,N28963);
and and17457(N28960,N28964,R7);
and and17461(N28968,in0,N28972);
and and17462(N28969,R1,R2);
and and17463(N28970,R3,R4);
and and17464(N28971,N28973,N28974);
and and17468(N28978,in0,R0);
and and17469(N28979,N28982,R2);
and and17470(N28980,N28983,R5);
and and17471(N28981,R6,N28984);
and and17475(N28988,in0,N28992);
and and17476(N28989,R1,R3);
and and17477(N28990,R4,R5);
and and17478(N28991,N28993,N28994);
and and17482(N28998,in0,R0);
and and17483(N28999,R1,N29002);
and and17484(N29000,R4,N29003);
and and17485(N29001,N29004,R7);
and and17489(N29008,in0,N29012);
and and17490(N29009,N29013,R2);
and and17491(N29010,R3,R4);
and and17492(N29011,N29014,R6);
and and17496(N29018,in0,N29022);
and and17497(N29019,N29023,R3);
and and17498(N29020,R4,R5);
and and17499(N29021,N29024,R7);
and and17503(N29028,in0,R0);
and and17504(N29029,N29032,N29033);
and and17505(N29030,R3,R5);
and and17506(N29031,N29034,R7);
and and17510(N29038,in0,R0);
and and17511(N29039,N29042,R2);
and and17512(N29040,R3,R4);
and and17513(N29041,N29043,R7);
and and17517(N29047,in0,in1);
and and17518(N29048,R0,R1);
and and17519(N29049,R2,R3);
and and17520(N29050,R5,R7);
and and14378(N24198,N24205,N24206);
and and14379(N24199,N24207,N24208);
and and14387(N24216,N24223,N24224);
and and14388(N24217,N24225,N24226);
and and14396(N24234,N24242,N24243);
and and14397(N24235,R6,N24244);
and and14405(N24252,R4,N24260);
and and14406(N24253,N24261,N24262);
and and14414(N24270,N24277,N24278);
and and14415(N24271,N24279,N24280);
and and14423(N24288,N24295,N24296);
and and14424(N24289,N24297,N24298);
and and14432(N24306,N24313,N24314);
and and14433(N24307,N24315,N24316);
and and14441(N24324,N24331,N24332);
and and14442(N24325,N24333,R7);
and and14450(N24341,N24348,N24349);
and and14451(N24342,N24350,R7);
and and14459(N24358,N24364,N24365);
and and14460(N24359,N24366,N24367);
and and14468(N24375,N24381,N24382);
and and14469(N24376,N24383,N24384);
and and14477(N24392,N24399,N24400);
and and14478(N24393,N24401,R7);
and and14486(N24409,N24416,N24417);
and and14487(N24410,N24418,R7);
and and14495(N24426,N24434,R5);
and and14496(N24427,N24435,R7);
and and14504(N24443,R3,R4);
and and14505(N24444,N24451,N24452);
and and14513(N24460,R3,N24468);
and and14514(N24461,R5,N24469);
and and14522(N24477,N24482,N24483);
and and14523(N24478,N24484,N24485);
and and14531(N24493,N24498,N24499);
and and14532(N24494,N24500,N24501);
and and14540(N24509,N24515,N24516);
and and14541(N24510,R6,N24517);
and and14549(N24525,N24531,N24532);
and and14550(N24526,R6,N24533);
and and14558(N24541,N24546,N24547);
and and14559(N24542,N24548,N24549);
and and14567(N24557,N24562,N24563);
and and14568(N24558,N24564,N24565);
and and14576(N24573,N24579,R5);
and and14577(N24574,N24580,N24581);
and and14585(N24589,N24595,R5);
and and14586(N24590,N24596,N24597);
and and14594(N24605,N24610,N24611);
and and14595(N24606,N24612,N24613);
and and14603(N24621,N24626,N24627);
and and14604(N24622,N24628,N24629);
and and14612(N24637,N24644,R5);
and and14613(N24638,R6,N24645);
and and14621(N24653,N24658,N24659);
and and14622(N24654,N24660,N24661);
and and14630(N24669,N24675,N24676);
and and14631(N24670,N24677,R6);
and and14639(N24685,N24691,N24692);
and and14640(N24686,N24693,R7);
and and14648(N24701,N24707,R5);
and and14649(N24702,N24708,N24709);
and and14657(N24717,N24722,N24723);
and and14658(N24718,N24724,N24725);
and and14666(N24733,N24740,R4);
and and14667(N24734,N24741,R7);
and and14675(N24749,N24755,R5);
and and14676(N24750,N24756,N24757);
and and14684(N24765,R4,N24771);
and and14685(N24766,N24772,N24773);
and and14693(N24781,N24788,R5);
and and14694(N24782,N24789,R7);
and and14702(N24797,N24804,N24805);
and and14703(N24798,R6,R7);
and and14711(N24813,N24819,N24820);
and and14712(N24814,R6,N24821);
and and14720(N24829,R4,N24836);
and and14721(N24830,R6,N24837);
and and14729(N24845,R4,N24851);
and and14730(N24846,N24852,N24853);
and and14738(N24861,R4,N24867);
and and14739(N24862,N24868,N24869);
and and14747(N24877,R3,N24884);
and and14748(N24878,R6,N24885);
and and14756(N24893,R3,N24900);
and and14757(N24894,R6,N24901);
and and14765(N24909,R3,N24916);
and and14766(N24910,R6,N24917);
and and14774(N24925,R3,N24932);
and and14775(N24926,N24933,R7);
and and14783(N24941,R4,N24948);
and and14784(N24942,N24949,R7);
and and14792(N24957,N24961,N24962);
and and14793(N24958,N24963,N24964);
and and14801(N24972,N24978,R5);
and and14802(N24973,N24979,R7);
and and14810(N24987,N24992,N24993);
and and14811(N24988,N24994,R7);
and and14819(N25002,N25007,N25008);
and and14820(N25003,N25009,R7);
and and14828(N25017,N25022,N25023);
and and14829(N25018,N25024,R7);
and and14837(N25032,N25037,N25038);
and and14838(N25033,N25039,R7);
and and14846(N25047,N25053,R5);
and and14847(N25048,N25054,R7);
and and14855(N25062,N25067,N25068);
and and14856(N25063,N25069,R7);
and and14864(N25077,N25084,R5);
and and14865(N25078,R6,R7);
and and14873(N25092,N25098,R5);
and and14874(N25093,N25099,R7);
and and14882(N25107,N25113,R5);
and and14883(N25108,R6,N25114);
and and14891(N25122,N25127,N25128);
and and14892(N25123,R5,N25129);
and and14900(N25137,N25142,N25143);
and and14901(N25138,N25144,R7);
and and14909(N25152,N25158,R5);
and and14910(N25153,N25159,R7);
and and14918(N25167,R3,R4);
and and14919(N25168,N25173,N25174);
and and14927(N25182,R4,N25188);
and and14928(N25183,N25189,R7);
and and14936(N25197,N25203,R5);
and and14937(N25198,N25204,R7);
and and14945(N25212,N25219,R5);
and and14946(N25213,R6,R7);
and and14954(N25227,R4,R5);
and and14955(N25228,R6,N25234);
and and14963(N25242,R3,N25248);
and and14964(N25243,N25249,R7);
and and14972(N25257,R4,R5);
and and14973(N25258,N25263,N25264);
and and14981(N25272,R4,N25277);
and and14982(N25273,N25278,N25279);
and and14990(N25287,R3,N25292);
and and14991(N25288,N25293,N25294);
and and14999(N25302,N25308,N25309);
and and15000(N25303,R6,R7);
and and15008(N25317,N25323,N25324);
and and15009(N25318,R6,R7);
and and15017(N25332,N25337,R5);
and and15018(N25333,N25338,N25339);
and and15026(N25347,R4,R5);
and and15027(N25348,N25353,N25354);
and and15035(N25362,N25369,R5);
and and15036(N25363,R6,R7);
and and15044(N25377,R3,N25382);
and and15045(N25378,N25383,N25384);
and and15053(N25392,N25397,N25398);
and and15054(N25393,N25399,R7);
and and15062(N25407,R3,N25413);
and and15063(N25408,R5,N25414);
and and15071(N25422,N25427,R5);
and and15072(N25423,N25428,R7);
and and15080(N25436,R4,R5);
and and15081(N25437,N25442,R7);
and and15089(N25450,N25454,N25455);
and and15090(N25451,N25456,R7);
and and15098(N25464,N25469,N25470);
and and15099(N25465,R6,R7);
and and15107(N25478,N25483,N25484);
and and15108(N25479,R6,R7);
and and15116(N25492,N25496,N25497);
and and15117(N25493,R6,N25498);
and and15125(N25506,R4,N25512);
and and15126(N25507,R6,R7);
and and15134(N25520,R4,R5);
and and15135(N25521,N25526,R7);
and and15143(N25534,R4,N25539);
and and15144(N25535,R6,N25540);
and and15152(N25548,N25553,N25554);
and and15153(N25549,R6,R7);
and and15161(N25562,N25566,N25567);
and and15162(N25563,R6,N25568);
and and15170(N25576,R3,R5);
and and15171(N25577,R6,N25582);
and and15179(N25590,R3,N25596);
and and15180(N25591,R5,R6);
and and15188(N25604,R3,N25608);
and and15189(N25605,N25609,N25610);
and and15197(N25618,N25622,N25623);
and and15198(N25619,N25624,R7);
and and15206(N25632,N25636,R5);
and and15207(N25633,N25637,N25638);
and and15215(N25646,R4,R5);
and and15216(N25647,N25651,N25652);
and and15224(N25660,R4,R5);
and and15225(N25661,N25665,N25666);
and and15233(N25674,R4,R5);
and and15234(N25675,R6,R7);
and and15242(N25688,N25693,N25694);
and and15243(N25689,R6,R7);
and and15251(N25702,N25707,N25708);
and and15252(N25703,R6,R7);
and and15260(N25716,N25720,N25721);
and and15261(N25717,R6,N25722);
and and15269(N25730,R3,R4);
and and15270(N25731,R6,N25736);
and and15278(N25744,N25748,N25749);
and and15279(N25745,R6,N25750);
and and15287(N25758,R3,R4);
and and15288(N25759,N25763,N25764);
and and15296(N25772,N25776,R5);
and and15297(N25773,N25777,N25778);
and and15305(N25786,N25791,N25792);
and and15306(N25787,R6,R7);
and and15314(N25800,R4,N25805);
and and15315(N25801,R6,N25806);
and and15323(N25814,N25819,R4);
and and15324(N25815,R6,N25820);
and and15332(N25828,R3,N25833);
and and15333(N25829,N25834,R7);
and and15341(N25842,N25846,N25847);
and and15342(N25843,R6,N25848);
and and15350(N25856,R3,N25861);
and and15351(N25857,R6,N25862);
and and15359(N25870,N25874,R4);
and and15360(N25871,N25875,N25876);
and and15368(N25884,R4,N25888);
and and15369(N25885,N25889,N25890);
and and15377(N25898,R4,N25902);
and and15378(N25899,N25903,N25904);
and and15386(N25912,R4,N25916);
and and15387(N25913,N25917,N25918);
and and15395(N25926,N25930,R4);
and and15396(N25927,N25931,N25932);
and and15404(N25940,R4,N25944);
and and15405(N25941,N25945,N25946);
and and15413(N25954,R3,N25958);
and and15414(N25955,N25959,N25960);
and and15422(N25968,N25973,R4);
and and15423(N25969,R5,N25974);
and and15431(N25982,N25987,R4);
and and15432(N25983,R5,N25988);
and and15440(N25996,R4,N26001);
and and15441(N25997,N26002,R7);
and and15449(N26010,N26014,R5);
and and15450(N26011,N26015,N26016);
and and15458(N26024,R3,N26029);
and and15459(N26025,N26030,R7);
and and15467(N26038,N26044,R5);
and and15468(N26039,R6,R7);
and and15476(N26052,N26057,R5);
and and15477(N26053,N26058,R7);
and and15485(N26066,R4,R5);
and and15486(N26067,R6,N26072);
and and15494(N26080,N26085,R5);
and and15495(N26081,R6,N26086);
and and15503(N26094,R3,N26100);
and and15504(N26095,R5,R6);
and and15512(N26108,N26111,N26112);
and and15513(N26109,N26113,N26114);
and and15521(N26122,N26127,N26128);
and and15522(N26123,R6,R7);
and and15530(N26136,R4,N26141);
and and15531(N26137,N26142,R7);
and and15539(N26150,R4,R5);
and and15540(N26151,R6,N26156);
and and15548(N26164,R3,N26169);
and and15549(N26165,N26170,R6);
and and15557(N26178,R4,R5);
and and15558(N26179,N26183,R7);
and and15566(N26191,R3,R5);
and and15567(N26192,R6,N26196);
and and15575(N26204,N26208,R5);
and and15576(N26205,N26209,R7);
and and15584(N26217,N26221,N26222);
and and15585(N26218,R6,R7);
and and15593(N26230,N26233,N26234);
and and15594(N26231,N26235,R7);
and and15602(N26243,N26246,N26247);
and and15603(N26244,N26248,R7);
and and15611(N26256,R3,N26260);
and and15612(N26257,R5,N26261);
and and15620(N26269,N26274,R5);
and and15621(N26270,R6,R7);
and and15629(N26282,R4,N26287);
and and15630(N26283,R6,R7);
and and15638(N26295,R3,R4);
and and15639(N26296,R6,R7);
and and15647(N26308,N26311,N26312);
and and15648(N26309,N26313,R7);
and and15656(N26321,R4,R5);
and and15657(N26322,R6,R7);
and and15665(N26334,N26337,N26338);
and and15666(N26335,N26339,R7);
and and15674(N26347,R4,R5);
and and15675(N26348,R6,R7);
and and15683(N26360,N26365,R5);
and and15684(N26361,R6,R7);
and and15692(N26373,N26378,R5);
and and15693(N26374,R6,R7);
and and15701(N26386,N26391,R5);
and and15702(N26387,R6,R7);
and and15710(N26399,R4,N26403);
and and15711(N26400,R6,N26404);
and and15719(N26412,R4,N26416);
and and15720(N26413,R6,N26417);
and and15728(N26425,R4,R5);
and and15729(N26426,N26430,R7);
and and15737(N26438,R4,R5);
and and15738(N26439,N26443,R7);
and and15746(N26451,N26455,R5);
and and15747(N26452,R6,N26456);
and and15755(N26464,N26468,N26469);
and and15756(N26465,R6,R7);
and and15764(N26477,R4,R5);
and and15765(N26478,R6,N26482);
and and15773(N26490,R4,R5);
and and15774(N26491,N26495,R7);
and and15782(N26503,R3,N26507);
and and15783(N26504,N26508,R7);
and and15791(N26516,N26521,R5);
and and15792(N26517,R6,R7);
and and15800(N26529,N26533,R5);
and and15801(N26530,N26534,R7);
and and15809(N26542,N26546,R5);
and and15810(N26543,R6,N26547);
and and15818(N26555,R3,N26558);
and and15819(N26556,N26559,N26560);
and and15827(N26568,R3,R5);
and and15828(N26569,R6,N26573);
and and15836(N26581,N26585,R5);
and and15837(N26582,R6,N26586);
and and15845(N26594,N26598,R5);
and and15846(N26595,R6,N26599);
and and15854(N26607,R4,R5);
and and15855(N26608,N26612,R7);
and and15863(N26620,R4,R5);
and and15864(N26621,N26623,N26624);
and and15872(N26632,N26635,R5);
and and15873(N26633,R6,N26636);
and and15881(N26644,R4,N26648);
and and15882(N26645,R6,R7);
and and15890(N26656,N26659,N26660);
and and15891(N26657,R6,R7);
and and15899(N26668,R4,N26672);
and and15900(N26669,R6,R7);
and and15908(N26680,N26683,R5);
and and15909(N26681,N26684,R7);
and and15917(N26692,R4,R5);
and and15918(N26693,R6,N26696);
and and15926(N26704,N26708,R5);
and and15927(N26705,R6,R7);
and and15935(N26716,R4,N26719);
and and15936(N26717,R6,N26720);
and and15944(N26728,N26732,R5);
and and15945(N26729,R6,R7);
and and15953(N26740,N26743,R4);
and and15954(N26741,R5,N26744);
and and15962(N26752,R3,N26755);
and and15963(N26753,N26756,R7);
and and15971(N26764,R4,R5);
and and15972(N26765,R6,R7);
and and15980(N26776,R4,N26780);
and and15981(N26777,R6,R7);
and and15989(N26788,R4,N26792);
and and15990(N26789,R6,R7);
and and15998(N26800,N26804,R5);
and and15999(N26801,R6,R7);
and and16007(N26812,N26815,R4);
and and16008(N26813,N26816,R6);
and and16016(N26824,R3,R4);
and and16017(N26825,R6,N26828);
and and16025(N26836,R3,N26839);
and and16026(N26837,R6,N26840);
and and16034(N26848,R4,R5);
and and16035(N26849,N26852,R7);
and and16043(N26860,N26863,N26864);
and and16044(N26861,R6,R7);
and and16052(N26872,R4,N26875);
and and16053(N26873,R6,N26876);
and and16061(N26884,R4,R5);
and and16062(N26885,R6,R7);
and and16070(N26896,N26899,R5);
and and16071(N26897,R6,N26900);
and and16079(N26908,R4,R5);
and and16080(N26909,N26912,R7);
and and16088(N26920,R3,N26922);
and and16089(N26921,N26923,N26924);
and and16097(N26932,R4,R5);
and and16098(N26933,N26936,R7);
and and16106(N26944,N26948,R5);
and and16107(N26945,R6,R7);
and and16115(N26956,N26960,R5);
and and16116(N26957,R6,R7);
and and16124(N26968,N26972,R5);
and and16125(N26969,R6,R7);
and and16133(N26980,R3,R4);
and and16134(N26981,R5,R7);
and and16142(N26992,R3,N26996);
and and16143(N26993,R6,R7);
and and16151(N27004,R4,R5);
and and16152(N27005,R6,N27008);
and and16160(N27016,N27020,R4);
and and16161(N27017,R5,R6);
and and16169(N27028,N27031,R5);
and and16170(N27029,R6,N27032);
and and16178(N27040,N27043,N27044);
and and16179(N27041,R6,R7);
and and16187(N27052,N27055,N27056);
and and16188(N27053,R6,R7);
and and16196(N27064,R4,R5);
and and16197(N27065,R6,R7);
and and16205(N27075,R4,R5);
and and16206(N27076,R6,N27078);
and and16214(N27086,R4,R5);
and and16215(N27087,R6,R7);
and and16223(N27097,R4,N27100);
and and16224(N27098,R6,R7);
and and16232(N27108,R3,R4);
and and16233(N27109,R5,R6);
and and16241(N27118,N27120,R5);
and and16242(N27119,R6,R7);
and and16250(N27128,R4,R5);
and and16251(N27129,R6,R7);
and and16259(N27138,R3,R4);
and and16260(N27139,R5,R6);
and and16268(N27148,R3,N27150);
and and16269(N27149,R5,R6);
and and16277(N27158,R3,R4);
and and16278(N27159,R5,R7);
and and16286(N27168,R3,R4);
and and16287(N27169,R6,R7);
and and16295(N27178,R4,R5);
and and16296(N27179,N27180,R7);
and and16304(N27188,N27190,R5);
and and16305(N27189,R6,R7);
and and16313(N27198,R3,N27200);
and and16314(N27199,R6,R7);
and and16322(N27208,N27215,N27216);
and and16330(N27224,N27231,N27232);
and and16338(N27240,N27246,N27247);
and and16346(N27255,N27261,N27262);
and and16354(N27270,N27277,R7);
and and16362(N27285,N27290,N27291);
and and16370(N27299,N27304,N27305);
and and16378(N27313,N27319,R7);
and and16386(N27327,R5,N27333);
and and16394(N27341,N27346,N27347);
and and16402(N27355,N27360,N27361);
and and16410(N27369,R6,N27375);
and and16418(N27383,N27388,N27389);
and and16426(N27397,R5,N27403);
and and16434(N27411,R6,N27417);
and and16442(N27425,N27430,N27431);
and and16450(N27439,R5,N27445);
and and16458(N27453,N27458,N27459);
and and16466(N27467,N27472,N27473);
and and16474(N27481,N27487,R7);
and and16482(N27495,R6,N27501);
and and16490(N27509,N27514,N27515);
and and16498(N27523,N27528,N27529);
and and16506(N27537,N27542,N27543);
and and16514(N27551,R6,N27557);
and and16522(N27565,N27571,R7);
and and16530(N27579,N27584,N27585);
and and16538(N27593,N27598,N27599);
and and16546(N27607,N27612,R7);
and and16554(N27620,N27624,N27625);
and and16562(N27633,N27638,R7);
and and16570(N27646,R5,N27651);
and and16578(N27659,N27664,R7);
and and16586(N27672,N27676,N27677);
and and16594(N27685,N27690,R7);
and and16602(N27698,N27702,N27703);
and and16610(N27711,R5,R6);
and and16618(N27724,N27728,N27729);
and and16626(N27737,N27741,N27742);
and and16634(N27750,R6,R7);
and and16642(N27763,R6,N27768);
and and16650(N27776,R5,N27781);
and and16658(N27789,R5,N27794);
and and16666(N27802,N27807,R7);
and and16674(N27815,R6,N27820);
and and16682(N27828,N27833,R7);
and and16690(N27841,N27845,N27846);
and and16698(N27854,R6,N27859);
and and16706(N27867,N27872,R7);
and and16714(N27880,R5,R7);
and and16722(N27893,R6,N27898);
and and16730(N27906,N27910,N27911);
and and16738(N27919,N27924,R7);
and and16746(N27932,N27937,R7);
and and16754(N27945,N27950,R7);
and and16762(N27958,R5,N27963);
and and16770(N27971,N27975,N27976);
and and16778(N27984,N27989,R7);
and and16786(N27997,N28001,N28002);
and and16794(N28010,N28014,N28015);
and and16802(N28023,N28027,N28028);
and and16810(N28036,N28041,R6);
and and16818(N28049,R6,N28054);
and and16826(N28062,N28067,R7);
and and16834(N28075,N28079,N28080);
and and16842(N28088,N28092,N28093);
and and16850(N28101,R5,N28105);
and and16858(N28113,N28116,N28117);
and and16866(N28125,N28128,N28129);
and and16874(N28137,N28141,R7);
and and16882(N28149,R6,N28153);
and and16890(N28161,R6,N28165);
and and16898(N28173,R5,R6);
and and16906(N28185,R6,N28189);
and and16914(N28197,N28200,N28201);
and and16922(N28209,N28213,R7);
and and16930(N28221,R6,N28225);
and and16938(N28233,R6,R7);
and and16946(N28245,N28248,N28249);
and and16954(N28257,N28260,N28261);
and and16962(N28269,N28272,N28273);
and and16970(N28281,R5,N28285);
and and16978(N28293,R6,R7);
and and16986(N28305,N28308,N28309);
and and16994(N28317,R6,N28321);
and and17002(N28329,R5,R7);
and and17010(N28341,R6,R7);
and and17018(N28353,N28357,R7);
and and17026(N28365,R6,N28369);
and and17034(N28377,R6,R7);
and and17042(N28389,N28393,R7);
and and17050(N28401,N28405,R7);
and and17058(N28413,R5,R6);
and and17066(N28425,N28428,N28429);
and and17074(N28437,R4,R7);
and and17082(N28449,N28453,R7);
and and17090(N28461,N28464,R7);
and and17098(N28472,R6,N28475);
and and17106(N28483,N28486,R7);
and and17114(N28494,R6,R7);
and and17122(N28505,R6,N28508);
and and17130(N28516,N28518,N28519);
and and17138(N28527,R4,N28530);
and and17146(N28538,N28540,N28541);
and and17154(N28549,N28552,R7);
and and17162(N28560,R6,N28563);
and and17170(N28571,N28574,R7);
and and17178(N28582,R6,R7);
and and17186(N28593,N28596,R7);
and and17194(N28604,N28607,R7);
and and17202(N28615,R6,N28618);
and and17210(N28626,R6,N28629);
and and17218(N28637,R6,N28640);
and and17226(N28648,R6,N28651);
and and17234(N28659,R5,N28662);
and and17242(N28670,R6,R7);
and and17250(N28681,N28684,R7);
and and17258(N28692,R5,R6);
and and17266(N28702,R6,R7);
and and17274(N28712,R6,R7);
and and17282(N28722,R5,R7);
and and17290(N28732,R6,R7);
and and17298(N28742,R6,R7);
and and17306(N28752,R6,R7);
and and17314(N28762,N28764,R7);
and and17322(N28772,R6,R7);
and and17330(N28782,R6,R7);
and and17338(N28792,R6,R7);
and and17346(N28802,R5,R6);
and and17354(N28812,R5,R6);
and and17362(N28822,R6,N28824);
and and17370(N28832,R4,N28834);
and and17378(N28842,R6,R7);
and and17386(N28851,R6,R7);
and and17394(N28859,R6,R7);
and and17521(N29216,N29217,N29218);
and and17531(N29234,N29235,N29236);
and and17541(N29252,N29253,N29254);
and and17551(N29267,N29268,N29269);
and and17560(N29285,N29286,N29287);
and and17569(N29303,N29304,N29305);
and and17578(N29321,N29322,N29323);
and and17587(N29339,N29340,N29341);
and and17596(N29357,N29358,N29359);
and and17605(N29374,N29375,N29376);
and and17614(N29391,N29392,N29393);
and and17623(N29408,N29409,N29410);
and and17632(N29425,N29426,N29427);
and and17641(N29442,N29443,N29444);
and and17650(N29459,N29460,N29461);
and and17659(N29476,N29477,N29478);
and and17668(N29493,N29494,N29495);
and and17677(N29510,N29511,N29512);
and and17686(N29527,N29528,N29529);
and and17695(N29543,N29544,N29545);
and and17704(N29559,N29560,N29561);
and and17713(N29575,N29576,N29577);
and and17722(N29591,N29592,N29593);
and and17731(N29607,N29608,N29609);
and and17740(N29623,N29624,N29625);
and and17749(N29639,N29640,N29641);
and and17758(N29655,N29656,N29657);
and and17767(N29671,N29672,N29673);
and and17776(N29687,N29688,N29689);
and and17785(N29703,N29704,N29705);
and and17794(N29719,N29720,N29721);
and and17803(N29735,N29736,N29737);
and and17812(N29751,N29752,N29753);
and and17821(N29766,N29767,N29768);
and and17830(N29781,N29782,N29783);
and and17839(N29796,N29797,N29798);
and and17848(N29811,N29812,N29813);
and and17857(N29826,N29827,N29828);
and and17866(N29841,N29842,N29843);
and and17875(N29856,N29857,N29858);
and and17884(N29871,N29872,N29873);
and and17893(N29886,N29887,N29888);
and and17902(N29901,N29902,N29903);
and and17911(N29916,N29917,N29918);
and and17920(N29931,N29932,N29933);
and and17929(N29946,N29947,N29948);
and and17938(N29961,N29962,N29963);
and and17947(N29976,N29977,N29978);
and and17956(N29991,N29992,N29993);
and and17965(N30006,N30007,N30008);
and and17974(N30021,N30022,N30023);
and and17983(N30036,N30037,N30038);
and and17992(N30051,N30052,N30053);
and and18001(N30066,N30067,N30068);
and and18010(N30080,N30081,N30082);
and and18019(N30094,N30095,N30096);
and and18028(N30108,N30109,N30110);
and and18037(N30122,N30123,N30124);
and and18046(N30136,N30137,N30138);
and and18055(N30150,N30151,N30152);
and and18064(N30164,N30165,N30166);
and and18073(N30178,N30179,N30180);
and and18082(N30192,N30193,N30194);
and and18091(N30206,N30207,N30208);
and and18100(N30220,N30221,N30222);
and and18109(N30234,N30235,N30236);
and and18118(N30248,N30249,N30250);
and and18127(N30262,N30263,N30264);
and and18136(N30276,N30277,N30278);
and and18145(N30290,N30291,N30292);
and and18154(N30304,N30305,N30306);
and and18163(N30318,N30319,N30320);
and and18172(N30332,N30333,N30334);
and and18181(N30346,N30347,N30348);
and and18190(N30360,N30361,N30362);
and and18199(N30374,N30375,N30376);
and and18208(N30388,N30389,N30390);
and and18217(N30402,N30403,N30404);
and and18226(N30416,N30417,N30418);
and and18235(N30430,N30431,N30432);
and and18244(N30444,N30445,N30446);
and and18253(N30458,N30459,N30460);
and and18262(N30472,N30473,N30474);
and and18271(N30486,N30487,N30488);
and and18280(N30500,N30501,N30502);
and and18289(N30514,N30515,N30516);
and and18298(N30528,N30529,N30530);
and and18307(N30542,N30543,N30544);
and and18316(N30556,N30557,N30558);
and and18325(N30570,N30571,N30572);
and and18334(N30584,N30585,N30586);
and and18343(N30598,N30599,N30600);
and and18352(N30612,N30613,N30614);
and and18361(N30626,N30627,N30628);
and and18370(N30640,N30641,N30642);
and and18379(N30654,N30655,N30656);
and and18388(N30668,N30669,N30670);
and and18397(N30682,N30683,N30684);
and and18406(N30696,N30697,N30698);
and and18415(N30710,N30711,N30712);
and and18424(N30723,N30724,N30725);
and and18433(N30736,N30737,N30738);
and and18442(N30749,N30750,N30751);
and and18451(N30762,N30763,N30764);
and and18460(N30775,N30776,N30777);
and and18469(N30788,N30789,N30790);
and and18478(N30801,N30802,N30803);
and and18487(N30814,N30815,N30816);
and and18496(N30827,N30828,N30829);
and and18505(N30840,N30841,N30842);
and and18514(N30853,N30854,N30855);
and and18523(N30866,N30867,N30868);
and and18532(N30879,N30880,N30881);
and and18541(N30892,N30893,N30894);
and and18550(N30905,N30906,N30907);
and and18559(N30918,N30919,N30920);
and and18568(N30931,N30932,N30933);
and and18577(N30944,N30945,N30946);
and and18586(N30957,N30958,N30959);
and and18595(N30970,N30971,N30972);
and and18604(N30983,N30984,N30985);
and and18613(N30996,N30997,N30998);
and and18622(N31009,N31010,N31011);
and and18631(N31022,N31023,N31024);
and and18640(N31034,N31035,N31036);
and and18649(N31046,N31047,N31048);
and and18658(N31058,N31059,N31060);
and and18667(N31070,N31071,N31072);
and and18676(N31082,N31083,N31084);
and and18685(N31094,N31095,N31096);
and and18694(N31106,N31107,N31108);
and and18703(N31118,N31119,N31120);
and and18712(N31130,N31131,N31132);
and and18721(N31142,N31143,N31144);
and and18730(N31154,N31155,N31156);
and and18739(N31166,N31167,N31168);
and and18748(N31178,N31179,N31180);
and and18757(N31190,N31191,N31192);
and and18766(N31202,N31203,N31204);
and and18775(N31213,N31214,N31215);
and and18784(N31224,N31225,N31226);
and and18793(N31235,N31236,N31237);
and and18801(N31250,N31251,N31252);
and and18809(N31265,N31266,N31267);
and and18817(N31280,N31281,N31282);
and and18825(N31295,N31296,N31297);
and and18833(N31309,N31310,N31311);
and and18841(N31323,N31324,N31325);
and and18849(N31337,N31338,N31339);
and and18857(N31351,N31352,N31353);
and and18865(N31365,N31366,N31367);
and and18873(N31379,N31380,N31381);
and and18881(N31393,N31394,N31395);
and and18889(N31406,N31407,N31408);
and and18897(N31419,N31420,N31421);
and and18905(N31432,N31433,N31434);
and and18913(N31445,N31446,N31447);
and and18921(N31458,N31459,N31460);
and and18929(N31471,N31472,N31473);
and and18937(N31484,N31485,N31486);
and and18945(N31496,N31497,N31498);
and and18953(N31508,N31509,N31510);
and and18961(N31520,N31521,N31522);
and and18969(N31532,N31533,N31534);
and and18977(N31543,N31544,N31545);
and and18985(N31554,N31555,N31556);
and and17522(N29217,N29219,N29220);
and and17523(N29218,N29221,N29222);
and and17532(N29235,N29237,N29238);
and and17533(N29236,N29239,N29240);
and and17542(N29253,N29255,N29256);
and and17543(N29254,N29257,N29258);
and and17552(N29268,N29270,N29271);
and and17553(N29269,N29272,N29273);
and and17561(N29286,N29288,N29289);
and and17562(N29287,N29290,N29291);
and and17570(N29304,N29306,N29307);
and and17571(N29305,N29308,N29309);
and and17579(N29322,N29324,N29325);
and and17580(N29323,N29326,N29327);
and and17588(N29340,N29342,N29343);
and and17589(N29341,N29344,N29345);
and and17597(N29358,N29360,N29361);
and and17598(N29359,N29362,N29363);
and and17606(N29375,N29377,N29378);
and and17607(N29376,N29379,N29380);
and and17615(N29392,N29394,N29395);
and and17616(N29393,N29396,N29397);
and and17624(N29409,N29411,N29412);
and and17625(N29410,N29413,N29414);
and and17633(N29426,N29428,N29429);
and and17634(N29427,N29430,N29431);
and and17642(N29443,N29445,N29446);
and and17643(N29444,N29447,N29448);
and and17651(N29460,N29462,N29463);
and and17652(N29461,N29464,N29465);
and and17660(N29477,N29479,N29480);
and and17661(N29478,N29481,N29482);
and and17669(N29494,N29496,N29497);
and and17670(N29495,N29498,N29499);
and and17678(N29511,N29513,N29514);
and and17679(N29512,N29515,N29516);
and and17687(N29528,N29530,N29531);
and and17688(N29529,N29532,N29533);
and and17696(N29544,N29546,N29547);
and and17697(N29545,N29548,N29549);
and and17705(N29560,N29562,N29563);
and and17706(N29561,N29564,N29565);
and and17714(N29576,N29578,N29579);
and and17715(N29577,N29580,N29581);
and and17723(N29592,N29594,N29595);
and and17724(N29593,N29596,N29597);
and and17732(N29608,N29610,N29611);
and and17733(N29609,N29612,N29613);
and and17741(N29624,N29626,N29627);
and and17742(N29625,N29628,N29629);
and and17750(N29640,N29642,N29643);
and and17751(N29641,N29644,N29645);
and and17759(N29656,N29658,N29659);
and and17760(N29657,N29660,N29661);
and and17768(N29672,N29674,N29675);
and and17769(N29673,N29676,N29677);
and and17777(N29688,N29690,N29691);
and and17778(N29689,N29692,N29693);
and and17786(N29704,N29706,N29707);
and and17787(N29705,N29708,N29709);
and and17795(N29720,N29722,N29723);
and and17796(N29721,N29724,N29725);
and and17804(N29736,N29738,N29739);
and and17805(N29737,N29740,N29741);
and and17813(N29752,N29754,N29755);
and and17814(N29753,N29756,N29757);
and and17822(N29767,N29769,N29770);
and and17823(N29768,N29771,N29772);
and and17831(N29782,N29784,N29785);
and and17832(N29783,N29786,N29787);
and and17840(N29797,N29799,N29800);
and and17841(N29798,N29801,N29802);
and and17849(N29812,N29814,N29815);
and and17850(N29813,N29816,N29817);
and and17858(N29827,N29829,N29830);
and and17859(N29828,N29831,N29832);
and and17867(N29842,N29844,N29845);
and and17868(N29843,N29846,N29847);
and and17876(N29857,N29859,N29860);
and and17877(N29858,N29861,N29862);
and and17885(N29872,N29874,N29875);
and and17886(N29873,N29876,N29877);
and and17894(N29887,N29889,N29890);
and and17895(N29888,N29891,N29892);
and and17903(N29902,N29904,N29905);
and and17904(N29903,N29906,N29907);
and and17912(N29917,N29919,N29920);
and and17913(N29918,N29921,N29922);
and and17921(N29932,N29934,N29935);
and and17922(N29933,N29936,N29937);
and and17930(N29947,N29949,N29950);
and and17931(N29948,N29951,N29952);
and and17939(N29962,N29964,N29965);
and and17940(N29963,N29966,N29967);
and and17948(N29977,N29979,N29980);
and and17949(N29978,N29981,N29982);
and and17957(N29992,N29994,N29995);
and and17958(N29993,N29996,N29997);
and and17966(N30007,N30009,N30010);
and and17967(N30008,N30011,N30012);
and and17975(N30022,N30024,N30025);
and and17976(N30023,N30026,N30027);
and and17984(N30037,N30039,N30040);
and and17985(N30038,N30041,N30042);
and and17993(N30052,N30054,N30055);
and and17994(N30053,N30056,N30057);
and and18002(N30067,N30069,N30070);
and and18003(N30068,N30071,N30072);
and and18011(N30081,N30083,N30084);
and and18012(N30082,N30085,N30086);
and and18020(N30095,N30097,N30098);
and and18021(N30096,N30099,N30100);
and and18029(N30109,N30111,N30112);
and and18030(N30110,N30113,N30114);
and and18038(N30123,N30125,N30126);
and and18039(N30124,N30127,N30128);
and and18047(N30137,N30139,N30140);
and and18048(N30138,N30141,N30142);
and and18056(N30151,N30153,N30154);
and and18057(N30152,N30155,N30156);
and and18065(N30165,N30167,N30168);
and and18066(N30166,N30169,N30170);
and and18074(N30179,N30181,N30182);
and and18075(N30180,N30183,N30184);
and and18083(N30193,N30195,N30196);
and and18084(N30194,N30197,N30198);
and and18092(N30207,N30209,N30210);
and and18093(N30208,N30211,N30212);
and and18101(N30221,N30223,N30224);
and and18102(N30222,N30225,N30226);
and and18110(N30235,N30237,N30238);
and and18111(N30236,N30239,N30240);
and and18119(N30249,N30251,N30252);
and and18120(N30250,N30253,N30254);
and and18128(N30263,N30265,N30266);
and and18129(N30264,N30267,N30268);
and and18137(N30277,N30279,N30280);
and and18138(N30278,N30281,N30282);
and and18146(N30291,N30293,N30294);
and and18147(N30292,N30295,N30296);
and and18155(N30305,N30307,N30308);
and and18156(N30306,N30309,N30310);
and and18164(N30319,N30321,N30322);
and and18165(N30320,N30323,N30324);
and and18173(N30333,N30335,N30336);
and and18174(N30334,N30337,N30338);
and and18182(N30347,N30349,N30350);
and and18183(N30348,N30351,N30352);
and and18191(N30361,N30363,N30364);
and and18192(N30362,N30365,N30366);
and and18200(N30375,N30377,N30378);
and and18201(N30376,N30379,N30380);
and and18209(N30389,N30391,N30392);
and and18210(N30390,N30393,N30394);
and and18218(N30403,N30405,N30406);
and and18219(N30404,N30407,N30408);
and and18227(N30417,N30419,N30420);
and and18228(N30418,N30421,N30422);
and and18236(N30431,N30433,N30434);
and and18237(N30432,N30435,N30436);
and and18245(N30445,N30447,N30448);
and and18246(N30446,N30449,N30450);
and and18254(N30459,N30461,N30462);
and and18255(N30460,N30463,N30464);
and and18263(N30473,N30475,N30476);
and and18264(N30474,N30477,N30478);
and and18272(N30487,N30489,N30490);
and and18273(N30488,N30491,N30492);
and and18281(N30501,N30503,N30504);
and and18282(N30502,N30505,N30506);
and and18290(N30515,N30517,N30518);
and and18291(N30516,N30519,N30520);
and and18299(N30529,N30531,N30532);
and and18300(N30530,N30533,N30534);
and and18308(N30543,N30545,N30546);
and and18309(N30544,N30547,N30548);
and and18317(N30557,N30559,N30560);
and and18318(N30558,N30561,N30562);
and and18326(N30571,N30573,N30574);
and and18327(N30572,N30575,N30576);
and and18335(N30585,N30587,N30588);
and and18336(N30586,N30589,N30590);
and and18344(N30599,N30601,N30602);
and and18345(N30600,N30603,N30604);
and and18353(N30613,N30615,N30616);
and and18354(N30614,N30617,N30618);
and and18362(N30627,N30629,N30630);
and and18363(N30628,N30631,N30632);
and and18371(N30641,N30643,N30644);
and and18372(N30642,N30645,N30646);
and and18380(N30655,N30657,N30658);
and and18381(N30656,N30659,N30660);
and and18389(N30669,N30671,N30672);
and and18390(N30670,N30673,N30674);
and and18398(N30683,N30685,N30686);
and and18399(N30684,N30687,N30688);
and and18407(N30697,N30699,N30700);
and and18408(N30698,N30701,N30702);
and and18416(N30711,N30713,N30714);
and and18417(N30712,N30715,N30716);
and and18425(N30724,N30726,N30727);
and and18426(N30725,N30728,N30729);
and and18434(N30737,N30739,N30740);
and and18435(N30738,N30741,N30742);
and and18443(N30750,N30752,N30753);
and and18444(N30751,N30754,N30755);
and and18452(N30763,N30765,N30766);
and and18453(N30764,N30767,N30768);
and and18461(N30776,N30778,N30779);
and and18462(N30777,N30780,N30781);
and and18470(N30789,N30791,N30792);
and and18471(N30790,N30793,N30794);
and and18479(N30802,N30804,N30805);
and and18480(N30803,N30806,N30807);
and and18488(N30815,N30817,N30818);
and and18489(N30816,N30819,N30820);
and and18497(N30828,N30830,N30831);
and and18498(N30829,N30832,N30833);
and and18506(N30841,N30843,N30844);
and and18507(N30842,N30845,N30846);
and and18515(N30854,N30856,N30857);
and and18516(N30855,N30858,N30859);
and and18524(N30867,N30869,N30870);
and and18525(N30868,N30871,N30872);
and and18533(N30880,N30882,N30883);
and and18534(N30881,N30884,N30885);
and and18542(N30893,N30895,N30896);
and and18543(N30894,N30897,N30898);
and and18551(N30906,N30908,N30909);
and and18552(N30907,N30910,N30911);
and and18560(N30919,N30921,N30922);
and and18561(N30920,N30923,N30924);
and and18569(N30932,N30934,N30935);
and and18570(N30933,N30936,N30937);
and and18578(N30945,N30947,N30948);
and and18579(N30946,N30949,N30950);
and and18587(N30958,N30960,N30961);
and and18588(N30959,N30962,N30963);
and and18596(N30971,N30973,N30974);
and and18597(N30972,N30975,N30976);
and and18605(N30984,N30986,N30987);
and and18606(N30985,N30988,N30989);
and and18614(N30997,N30999,N31000);
and and18615(N30998,N31001,N31002);
and and18623(N31010,N31012,N31013);
and and18624(N31011,N31014,N31015);
and and18632(N31023,N31025,N31026);
and and18633(N31024,N31027,N31028);
and and18641(N31035,N31037,N31038);
and and18642(N31036,N31039,N31040);
and and18650(N31047,N31049,N31050);
and and18651(N31048,N31051,N31052);
and and18659(N31059,N31061,N31062);
and and18660(N31060,N31063,N31064);
and and18668(N31071,N31073,N31074);
and and18669(N31072,N31075,N31076);
and and18677(N31083,N31085,N31086);
and and18678(N31084,N31087,N31088);
and and18686(N31095,N31097,N31098);
and and18687(N31096,N31099,N31100);
and and18695(N31107,N31109,N31110);
and and18696(N31108,N31111,N31112);
and and18704(N31119,N31121,N31122);
and and18705(N31120,N31123,N31124);
and and18713(N31131,N31133,N31134);
and and18714(N31132,N31135,N31136);
and and18722(N31143,N31145,N31146);
and and18723(N31144,N31147,N31148);
and and18731(N31155,N31157,N31158);
and and18732(N31156,N31159,N31160);
and and18740(N31167,N31169,N31170);
and and18741(N31168,N31171,N31172);
and and18749(N31179,N31181,N31182);
and and18750(N31180,N31183,N31184);
and and18758(N31191,N31193,N31194);
and and18759(N31192,N31195,N31196);
and and18767(N31203,N31205,N31206);
and and18768(N31204,N31207,N31208);
and and18776(N31214,N31216,N31217);
and and18777(N31215,N31218,N31219);
and and18785(N31225,N31227,N31228);
and and18786(N31226,N31229,N31230);
and and18794(N31236,N31238,N31239);
and and18795(N31237,N31240,N31241);
and and18802(N31251,N31253,N31254);
and and18803(N31252,N31255,N31256);
and and18810(N31266,N31268,N31269);
and and18811(N31267,N31270,N31271);
and and18818(N31281,N31283,N31284);
and and18819(N31282,N31285,N31286);
and and18826(N31296,N31298,N31299);
and and18827(N31297,N31300,N31301);
and and18834(N31310,N31312,N31313);
and and18835(N31311,N31314,N31315);
and and18842(N31324,N31326,N31327);
and and18843(N31325,N31328,N31329);
and and18850(N31338,N31340,N31341);
and and18851(N31339,N31342,N31343);
and and18858(N31352,N31354,N31355);
and and18859(N31353,N31356,N31357);
and and18866(N31366,N31368,N31369);
and and18867(N31367,N31370,N31371);
and and18874(N31380,N31382,N31383);
and and18875(N31381,N31384,N31385);
and and18882(N31394,N31396,N31397);
and and18883(N31395,N31398,N31399);
and and18890(N31407,N31409,N31410);
and and18891(N31408,N31411,N31412);
and and18898(N31420,N31422,N31423);
and and18899(N31421,N31424,N31425);
and and18906(N31433,N31435,N31436);
and and18907(N31434,N31437,N31438);
and and18914(N31446,N31448,N31449);
and and18915(N31447,N31450,N31451);
and and18922(N31459,N31461,N31462);
and and18923(N31460,N31463,N31464);
and and18930(N31472,N31474,N31475);
and and18931(N31473,N31476,N31477);
and and18938(N31485,N31487,N31488);
and and18939(N31486,N31489,N31490);
and and18946(N31497,N31499,N31500);
and and18947(N31498,N31501,N31502);
and and18954(N31509,N31511,N31512);
and and18955(N31510,N31513,N31514);
and and18962(N31521,N31523,N31524);
and and18963(N31522,N31525,N31526);
and and18970(N31533,N31535,N31536);
and and18971(N31534,N31537,N31538);
and and18978(N31544,N31546,N31547);
and and18979(N31545,N31548,N31549);
and and18986(N31555,N31557,N31558);
and and18987(N31556,N31559,N31560);
and and17524(N29219,N29223,N29224);
and and17525(N29220,N29225,N29226);
and and17526(N29221,in1,N29227);
and and17527(N29222,N29228,R1);
and and17534(N29237,N29241,N29242);
and and17535(N29238,N29243,N29244);
and and17536(N29239,N29245,N29246);
and and17537(N29240,N29247,N29248);
and and17544(N29255,N29259,N29260);
and and17545(N29256,N29261,N29262);
and and17546(N29257,N29263,in2);
and and17547(N29258,R0,R1);
and and17554(N29270,N29274,N29275);
and and17555(N29271,N29276,N29277);
and and17556(N29272,in2,N29278);
and and17557(N29273,N29279,N29280);
and and17563(N29288,N29292,N29293);
and and17564(N29289,N29294,in1);
and and17565(N29290,N29295,N29296);
and and17566(N29291,N29297,N29298);
and and17572(N29306,N29310,N29311);
and and17573(N29307,N29312,N29313);
and and17574(N29308,N29314,N29315);
and and17575(N29309,R2,N29316);
and and17581(N29324,N29328,N29329);
and and17582(N29325,N29330,N29331);
and and17583(N29326,N29332,N29333);
and and17584(N29327,N29334,N29335);
and and17590(N29342,N29346,N29347);
and and17591(N29343,N29348,N29349);
and and17592(N29344,in2,N29350);
and and17593(N29345,N29351,N29352);
and and17599(N29360,N29364,N29365);
and and17600(N29361,N29366,N29367);
and and17601(N29362,N29368,R1);
and and17602(N29363,N29369,N29370);
and and17608(N29377,N29381,N29382);
and and17609(N29378,N29383,in2);
and and17610(N29379,N29384,N29385);
and and17611(N29380,N29386,N29387);
and and17617(N29394,N29398,N29399);
and and17618(N29395,N29400,N29401);
and and17619(N29396,N29402,R0);
and and17620(N29397,N29403,N29404);
and and17626(N29411,N29415,N29416);
and and17627(N29412,N29417,N29418);
and and17628(N29413,in2,N29419);
and and17629(N29414,N29420,R3);
and and17635(N29428,N29432,N29433);
and and17636(N29429,N29434,N29435);
and and17637(N29430,N29436,N29437);
and and17638(N29431,R2,R3);
and and17644(N29445,N29449,N29450);
and and17645(N29446,N29451,N29452);
and and17646(N29447,N29453,N29454);
and and17647(N29448,N29455,R2);
and and17653(N29462,N29466,N29467);
and and17654(N29463,N29468,N29469);
and and17655(N29464,in2,N29470);
and and17656(N29465,N29471,N29472);
and and17662(N29479,N29483,N29484);
and and17663(N29480,N29485,N29486);
and and17664(N29481,N29487,N29488);
and and17665(N29482,N29489,R3);
and and17671(N29496,N29500,N29501);
and and17672(N29497,N29502,N29503);
and and17673(N29498,N29504,N29505);
and and17674(N29499,N29506,N29507);
and and17680(N29513,N29517,N29518);
and and17681(N29514,N29519,N29520);
and and17682(N29515,N29521,N29522);
and and17683(N29516,N29523,R3);
and and17689(N29530,N29534,N29535);
and and17690(N29531,N29536,in1);
and and17691(N29532,in2,R0);
and and17692(N29533,N29537,N29538);
and and17698(N29546,N29550,N29551);
and and17699(N29547,N29552,in1);
and and17700(N29548,in2,N29553);
and and17701(N29549,N29554,N29555);
and and17707(N29562,N29566,N29567);
and and17708(N29563,N29568,N29569);
and and17709(N29564,in2,R0);
and and17710(N29565,R1,N29570);
and and17716(N29578,N29582,N29583);
and and17717(N29579,N29584,in1);
and and17718(N29580,N29585,R0);
and and17719(N29581,R1,N29586);
and and17725(N29594,N29598,N29599);
and and17726(N29595,N29600,N29601);
and and17727(N29596,R0,R1);
and and17728(N29597,N29602,N29603);
and and17734(N29610,N29614,N29615);
and and17735(N29611,N29616,N29617);
and and17736(N29612,in2,N29618);
and and17737(N29613,N29619,R2);
and and17743(N29626,N29630,N29631);
and and17744(N29627,N29632,N29633);
and and17745(N29628,N29634,R1);
and and17746(N29629,N29635,R3);
and and17752(N29642,N29646,N29647);
and and17753(N29643,N29648,N29649);
and and17754(N29644,N29650,R0);
and and17755(N29645,N29651,N29652);
and and17761(N29658,N29662,N29663);
and and17762(N29659,N29664,N29665);
and and17763(N29660,N29666,N29667);
and and17764(N29661,R2,R3);
and and17770(N29674,N29678,N29679);
and and17771(N29675,N29680,N29681);
and and17772(N29676,N29682,N29683);
and and17773(N29677,N29684,R3);
and and17779(N29690,N29694,N29695);
and and17780(N29691,N29696,in2);
and and17781(N29692,N29697,R1);
and and17782(N29693,N29698,N29699);
and and17788(N29706,N29710,N29711);
and and17789(N29707,N29712,N29713);
and and17790(N29708,in2,N29714);
and and17791(N29709,N29715,R3);
and and17797(N29722,N29726,N29727);
and and17798(N29723,N29728,in1);
and and17799(N29724,N29729,N29730);
and and17800(N29725,N29731,R2);
and and17806(N29738,N29742,N29743);
and and17807(N29739,N29744,N29745);
and and17808(N29740,N29746,R0);
and and17809(N29741,N29747,N29748);
and and17815(N29754,N29758,N29759);
and and17816(N29755,N29760,N29761);
and and17817(N29756,N29762,N29763);
and and17818(N29757,N29764,R2);
and and17824(N29769,N29773,N29774);
and and17825(N29770,N29775,N29776);
and and17826(N29771,N29777,N29778);
and and17827(N29772,R2,N29779);
and and17833(N29784,N29788,N29789);
and and17834(N29785,N29790,N29791);
and and17835(N29786,in2,N29792);
and and17836(N29787,N29793,R3);
and and17842(N29799,N29803,N29804);
and and17843(N29800,N29805,in1);
and and17844(N29801,in2,R1);
and and17845(N29802,R2,N29806);
and and17851(N29814,N29818,N29819);
and and17852(N29815,N29820,in1);
and and17853(N29816,N29821,N29822);
and and17854(N29817,N29823,R2);
and and17860(N29829,N29833,N29834);
and and17861(N29830,N29835,N29836);
and and17862(N29831,R0,N29837);
and and17863(N29832,N29838,R3);
and and17869(N29844,N29848,N29849);
and and17870(N29845,N29850,N29851);
and and17871(N29846,N29852,N29853);
and and17872(N29847,N29854,N29855);
and and17878(N29859,N29863,N29864);
and and17879(N29860,N29865,N29866);
and and17880(N29861,N29867,N29868);
and and17881(N29862,R1,R2);
and and17887(N29874,N29878,N29879);
and and17888(N29875,N29880,in1);
and and17889(N29876,N29881,N29882);
and and17890(N29877,R1,R2);
and and17896(N29889,N29893,N29894);
and and17897(N29890,N29895,in1);
and and17898(N29891,N29896,R0);
and and17899(N29892,N29897,R2);
and and17905(N29904,N29908,N29909);
and and17906(N29905,N29910,in2);
and and17907(N29906,R0,N29911);
and and17908(N29907,N29912,N29913);
and and17914(N29919,N29923,N29924);
and and17915(N29920,N29925,N29926);
and and17916(N29921,in2,R0);
and and17917(N29922,N29927,R3);
and and17923(N29934,N29938,N29939);
and and17924(N29935,N29940,N29941);
and and17925(N29936,in2,R0);
and and17926(N29937,N29942,R2);
and and17932(N29949,N29953,N29954);
and and17933(N29950,N29955,N29956);
and and17934(N29951,in2,R0);
and and17935(N29952,R1,N29957);
and and17941(N29964,N29968,N29969);
and and17942(N29965,N29970,in1);
and and17943(N29966,in2,N29971);
and and17944(N29967,N29972,N29973);
and and17950(N29979,N29983,N29984);
and and17951(N29980,N29985,N29986);
and and17952(N29981,in2,R0);
and and17953(N29982,R2,N29987);
and and17959(N29994,N29998,N29999);
and and17960(N29995,N30000,N30001);
and and17961(N29996,N30002,R0);
and and17962(N29997,R1,R3);
and and17968(N30009,N30013,N30014);
and and17969(N30010,N30015,N30016);
and and17970(N30011,R0,N30017);
and and17971(N30012,N30018,R3);
and and17977(N30024,N30028,N30029);
and and17978(N30025,N30030,N30031);
and and17979(N30026,R0,R1);
and and17980(N30027,N30032,R3);
and and17986(N30039,N30043,N30044);
and and17987(N30040,N30045,N30046);
and and17988(N30041,R0,R1);
and and17989(N30042,N30047,R3);
and and17995(N30054,N30058,N30059);
and and17996(N30055,N30060,N30061);
and and17997(N30056,in2,N30062);
and and17998(N30057,N30063,R3);
and and18004(N30069,N30073,N30074);
and and18005(N30070,N30075,in1);
and and18006(N30071,in2,N30076);
and and18007(N30072,N30077,R2);
and and18013(N30083,N30087,N30088);
and and18014(N30084,N30089,N30090);
and and18015(N30085,R0,R1);
and and18016(N30086,R2,N30091);
and and18022(N30097,N30101,N30102);
and and18023(N30098,N30103,N30104);
and and18024(N30099,in2,N30105);
and and18025(N30100,R1,R2);
and and18031(N30111,N30115,N30116);
and and18032(N30112,N30117,in1);
and and18033(N30113,N30118,N30119);
and and18034(N30114,R1,R2);
and and18040(N30125,N30129,N30130);
and and18041(N30126,N30131,in1);
and and18042(N30127,R0,R1);
and and18043(N30128,R2,N30132);
and and18049(N30139,N30143,N30144);
and and18050(N30140,N30145,N30146);
and and18051(N30141,N30147,R0);
and and18052(N30142,N30148,R2);
and and18058(N30153,N30157,N30158);
and and18059(N30154,N30159,in1);
and and18060(N30155,N30160,R0);
and and18061(N30156,R1,R2);
and and18067(N30167,N30171,N30172);
and and18068(N30168,N30173,in1);
and and18069(N30169,N30174,N30175);
and and18070(N30170,R1,R2);
and and18076(N30181,N30185,N30186);
and and18077(N30182,N30187,in1);
and and18078(N30183,in2,N30188);
and and18079(N30184,R1,R3);
and and18085(N30195,N30199,N30200);
and and18086(N30196,N30201,in1);
and and18087(N30197,in2,N30202);
and and18088(N30198,R2,R3);
and and18094(N30209,N30213,N30214);
and and18095(N30210,N30215,in1);
and and18096(N30211,R0,N30216);
and and18097(N30212,N30217,R3);
and and18103(N30223,N30227,N30228);
and and18104(N30224,N30229,in1);
and and18105(N30225,R0,N30230);
and and18106(N30226,R2,N30231);
and and18112(N30237,N30241,N30242);
and and18113(N30238,N30243,N30244);
and and18114(N30239,N30245,R0);
and and18115(N30240,N30246,R2);
and and18121(N30251,N30255,N30256);
and and18122(N30252,N30257,N30258);
and and18123(N30253,in2,N30259);
and and18124(N30254,R1,R2);
and and18130(N30265,N30269,N30270);
and and18131(N30266,N30271,N30272);
and and18132(N30267,R0,R1);
and and18133(N30268,N30273,R3);
and and18139(N30279,N30283,N30284);
and and18140(N30280,N30285,N30286);
and and18141(N30281,N30287,R0);
and and18142(N30282,N30288,R3);
and and18148(N30293,N30297,N30298);
and and18149(N30294,N30299,N30300);
and and18150(N30295,in2,N30301);
and and18151(N30296,R1,R2);
and and18157(N30307,N30311,N30312);
and and18158(N30308,N30313,in1);
and and18159(N30309,in2,R0);
and and18160(N30310,R1,N30314);
and and18166(N30321,N30325,N30326);
and and18167(N30322,N30327,in1);
and and18168(N30323,N30328,N30329);
and and18169(N30324,R1,R2);
and and18175(N30335,N30339,N30340);
and and18176(N30336,N30341,in1);
and and18177(N30337,N30342,N30343);
and and18178(N30338,R1,R3);
and and18184(N30349,N30353,N30354);
and and18185(N30350,N30355,in1);
and and18186(N30351,N30356,R0);
and and18187(N30352,N30357,R2);
and and18193(N30363,N30367,N30368);
and and18194(N30364,N30369,N30370);
and and18195(N30365,N30371,N30372);
and and18196(N30366,R1,R2);
and and18202(N30377,N30381,N30382);
and and18203(N30378,N30383,N30384);
and and18204(N30379,R0,R1);
and and18205(N30380,R2,R3);
and and18211(N30391,N30395,N30396);
and and18212(N30392,N30397,N30398);
and and18213(N30393,R0,N30399);
and and18214(N30394,R2,N30400);
and and18220(N30405,N30409,N30410);
and and18221(N30406,N30411,N30412);
and and18222(N30407,N30413,R0);
and and18223(N30408,R1,R2);
and and18229(N30419,N30423,N30424);
and and18230(N30420,N30425,in1);
and and18231(N30421,N30426,R0);
and and18232(N30422,N30427,N30428);
and and18238(N30433,N30437,N30438);
and and18239(N30434,N30439,N30440);
and and18240(N30435,N30441,R0);
and and18241(N30436,N30442,N30443);
and and18247(N30447,N30451,N30452);
and and18248(N30448,N30453,N30454);
and and18249(N30449,N30455,N30456);
and and18250(N30450,R1,N30457);
and and18256(N30461,N30465,N30466);
and and18257(N30462,N30467,in1);
and and18258(N30463,in2,N30468);
and and18259(N30464,R1,R2);
and and18265(N30475,N30479,N30480);
and and18266(N30476,N30481,in1);
and and18267(N30477,in2,N30482);
and and18268(N30478,N30483,R2);
and and18274(N30489,N30493,N30494);
and and18275(N30490,N30495,N30496);
and and18276(N30491,in2,R0);
and and18277(N30492,N30497,R3);
and and18283(N30503,N30507,N30508);
and and18284(N30504,N30509,N30510);
and and18285(N30505,in2,N30511);
and and18286(N30506,N30512,R2);
and and18292(N30517,N30521,N30522);
and and18293(N30518,N30523,in1);
and and18294(N30519,in2,R0);
and and18295(N30520,N30524,N30525);
and and18301(N30531,N30535,N30536);
and and18302(N30532,N30537,in1);
and and18303(N30533,N30538,N30539);
and and18304(N30534,R1,R2);
and and18310(N30545,N30549,N30550);
and and18311(N30546,N30551,in1);
and and18312(N30547,N30552,N30553);
and and18313(N30548,N30554,N30555);
and and18319(N30559,N30563,N30564);
and and18320(N30560,N30565,N30566);
and and18321(N30561,in2,N30567);
and and18322(N30562,N30568,R3);
and and18328(N30573,N30577,N30578);
and and18329(N30574,N30579,N30580);
and and18330(N30575,R0,R1);
and and18331(N30576,R2,N30581);
and and18337(N30587,N30591,N30592);
and and18338(N30588,N30593,in1);
and and18339(N30589,N30594,R0);
and and18340(N30590,N30595,R3);
and and18346(N30601,N30605,N30606);
and and18347(N30602,N30607,N30608);
and and18348(N30603,in2,R0);
and and18349(N30604,R2,N30609);
and and18355(N30615,N30619,N30620);
and and18356(N30616,N30621,in1);
and and18357(N30617,N30622,R0);
and and18358(N30618,N30623,R2);
and and18364(N30629,N30633,N30634);
and and18365(N30630,N30635,in1);
and and18366(N30631,N30636,N30637);
and and18367(N30632,R1,R3);
and and18373(N30643,N30647,N30648);
and and18374(N30644,N30649,in1);
and and18375(N30645,in2,N30650);
and and18376(N30646,N30651,R2);
and and18382(N30657,N30661,N30662);
and and18383(N30658,N30663,N30664);
and and18384(N30659,R0,R1);
and and18385(N30660,R2,R3);
and and18391(N30671,N30675,N30676);
and and18392(N30672,N30677,N30678);
and and18393(N30673,N30679,R0);
and and18394(N30674,R1,N30680);
and and18400(N30685,N30689,N30690);
and and18401(N30686,N30691,N30692);
and and18402(N30687,in2,R0);
and and18403(N30688,R1,R2);
and and18409(N30699,N30703,N30704);
and and18410(N30700,N30705,in1);
and and18411(N30701,in2,R0);
and and18412(N30702,R1,N30706);
and and18418(N30713,N30717,N30718);
and and18419(N30714,N30719,in1);
and and18420(N30715,N30720,R0);
and and18421(N30716,R1,R2);
and and18427(N30726,N30730,N30731);
and and18428(N30727,N30732,in1);
and and18429(N30728,N30733,N30734);
and and18430(N30729,R2,R3);
and and18436(N30739,N30743,N30744);
and and18437(N30740,N30745,in2);
and and18438(N30741,N30746,R1);
and and18439(N30742,R2,R3);
and and18445(N30752,N30756,N30757);
and and18446(N30753,N30758,N30759);
and and18447(N30754,N30760,R0);
and and18448(N30755,R1,R2);
and and18454(N30765,N30769,N30770);
and and18455(N30766,N30771,in1);
and and18456(N30767,R0,N30772);
and and18457(N30768,R2,R3);
and and18463(N30778,N30782,N30783);
and and18464(N30779,N30784,N30785);
and and18465(N30780,R0,N30786);
and and18466(N30781,R2,R3);
and and18472(N30791,N30795,N30796);
and and18473(N30792,N30797,N30798);
and and18474(N30793,in2,N30799);
and and18475(N30794,R1,N30800);
and and18481(N30804,N30808,N30809);
and and18482(N30805,N30810,N30811);
and and18483(N30806,in2,R0);
and and18484(N30807,N30812,R2);
and and18490(N30817,N30821,N30822);
and and18491(N30818,N30823,in1);
and and18492(N30819,in2,R0);
and and18493(N30820,R1,R2);
and and18499(N30830,N30834,N30835);
and and18500(N30831,N30836,in1);
and and18501(N30832,N30837,R0);
and and18502(N30833,N30838,R3);
and and18508(N30843,N30847,N30848);
and and18509(N30844,N30849,in1);
and and18510(N30845,in2,R0);
and and18511(N30846,N30850,N30851);
and and18517(N30856,N30860,N30861);
and and18518(N30857,N30862,in1);
and and18519(N30858,R0,R1);
and and18520(N30859,N30863,R3);
and and18526(N30869,N30873,N30874);
and and18527(N30870,N30875,N30876);
and and18528(N30871,in2,R0);
and and18529(N30872,R1,R2);
and and18535(N30882,N30886,N30887);
and and18536(N30883,N30888,in1);
and and18537(N30884,in2,N30889);
and and18538(N30885,R2,R3);
and and18544(N30895,N30899,N30900);
and and18545(N30896,N30901,N30902);
and and18546(N30897,in2,R0);
and and18547(N30898,R1,R2);
and and18553(N30908,N30912,N30913);
and and18554(N30909,N30914,in1);
and and18555(N30910,in2,R0);
and and18556(N30911,R1,N30915);
and and18562(N30921,N30925,N30926);
and and18563(N30922,N30927,in1);
and and18564(N30923,in2,R0);
and and18565(N30924,R1,R2);
and and18571(N30934,N30938,N30939);
and and18572(N30935,N30940,in2);
and and18573(N30936,R0,R1);
and and18574(N30937,R2,R3);
and and18580(N30947,N30951,N30952);
and and18581(N30948,N30953,in1);
and and18582(N30949,R0,N30954);
and and18583(N30950,R2,N30955);
and and18589(N30960,N30964,N30965);
and and18590(N30961,N30966,in1);
and and18591(N30962,N30967,R0);
and and18592(N30963,R2,R3);
and and18598(N30973,N30977,N30978);
and and18599(N30974,N30979,N30980);
and and18600(N30975,N30981,R0);
and and18601(N30976,R1,R2);
and and18607(N30986,N30990,N30991);
and and18608(N30987,N30992,in1);
and and18609(N30988,N30993,R0);
and and18610(N30989,R1,R2);
and and18616(N30999,N31003,N31004);
and and18617(N31000,N31005,N31006);
and and18618(N31001,in2,R0);
and and18619(N31002,R1,R2);
and and18625(N31012,N31016,N31017);
and and18626(N31013,N31018,in1);
and and18627(N31014,in2,R0);
and and18628(N31015,R1,N31019);
and and18634(N31025,N31029,N31030);
and and18635(N31026,N31031,in1);
and and18636(N31027,N31032,R1);
and and18637(N31028,R2,R3);
and and18643(N31037,N31041,N31042);
and and18644(N31038,N31043,in1);
and and18645(N31039,in2,N31044);
and and18646(N31040,R1,R2);
and and18652(N31049,N31053,N31054);
and and18653(N31050,N31055,N31056);
and and18654(N31051,in2,R0);
and and18655(N31052,N31057,R2);
and and18661(N31061,N31065,N31066);
and and18662(N31062,N31067,N31068);
and and18663(N31063,in2,R0);
and and18664(N31064,N31069,R2);
and and18670(N31073,N31077,N31078);
and and18671(N31074,N31079,in2);
and and18672(N31075,R0,N31080);
and and18673(N31076,R2,R3);
and and18679(N31085,N31089,N31090);
and and18680(N31086,N31091,in1);
and and18681(N31087,N31092,R0);
and and18682(N31088,R1,R2);
and and18688(N31097,N31101,N31102);
and and18689(N31098,N31103,N31104);
and and18690(N31099,in2,R0);
and and18691(N31100,N31105,R3);
and and18697(N31109,N31113,N31114);
and and18698(N31110,N31115,N31116);
and and18699(N31111,in2,R1);
and and18700(N31112,R2,R3);
and and18706(N31121,N31125,N31126);
and and18707(N31122,N31127,in1);
and and18708(N31123,in2,R0);
and and18709(N31124,N31128,R2);
and and18715(N31133,N31137,N31138);
and and18716(N31134,N31139,in1);
and and18717(N31135,in2,N31140);
and and18718(N31136,N31141,R3);
and and18724(N31145,N31149,N31150);
and and18725(N31146,N31151,in1);
and and18726(N31147,in2,R0);
and and18727(N31148,N31152,R2);
and and18733(N31157,N31161,N31162);
and and18734(N31158,N31163,N31164);
and and18735(N31159,R0,R1);
and and18736(N31160,R2,R3);
and and18742(N31169,N31173,N31174);
and and18743(N31170,N31175,N31176);
and and18744(N31171,in2,R0);
and and18745(N31172,R1,R2);
and and18751(N31181,N31185,N31186);
and and18752(N31182,N31187,in1);
and and18753(N31183,in2,N31188);
and and18754(N31184,N31189,R2);
and and18760(N31193,N31197,N31198);
and and18761(N31194,N31199,N31200);
and and18762(N31195,R0,N31201);
and and18763(N31196,R2,R3);
and and18769(N31205,N31209,N31210);
and and18770(N31206,N31211,in1);
and and18771(N31207,in2,N31212);
and and18772(N31208,R1,R2);
and and18778(N31216,N31220,N31221);
and and18779(N31217,N31222,in1);
and and18780(N31218,in2,R1);
and and18781(N31219,R2,R3);
and and18787(N31227,N31231,N31232);
and and18788(N31228,N31233,N31234);
and and18789(N31229,in2,R0);
and and18790(N31230,R1,R2);
and and18796(N31238,N31242,N31243);
and and18797(N31239,R0,N31244);
and and18798(N31240,R2,N31245);
and and18799(N31241,N31246,N31247);
and and18804(N31253,N31257,N31258);
and and18805(N31254,N31259,R0);
and and18806(N31255,N31260,N31261);
and and18807(N31256,R3,N31262);
and and18812(N31268,N31272,N31273);
and and18813(N31269,N31274,N31275);
and and18814(N31270,N31276,N31277);
and and18815(N31271,N31278,R5);
and and18820(N31283,N31287,N31288);
and and18821(N31284,N31289,R0);
and and18822(N31285,N31290,R2);
and and18823(N31286,N31291,N31292);
and and18828(N31298,N31302,N31303);
and and18829(N31299,in2,N31304);
and and18830(N31300,R2,N31305);
and and18831(N31301,N31306,N31307);
and and18836(N31312,N31316,N31317);
and and18837(N31313,N31318,in2);
and and18838(N31314,R0,N31319);
and and18839(N31315,N31320,N31321);
and and18844(N31326,N31330,N31331);
and and18845(N31327,N31332,in2);
and and18846(N31328,N31333,N31334);
and and18847(N31329,N31335,R5);
and and18852(N31340,N31344,N31345);
and and18853(N31341,N31346,R0);
and and18854(N31342,N31347,N31348);
and and18855(N31343,N31349,N31350);
and and18860(N31354,N31358,N31359);
and and18861(N31355,in1,N31360);
and and18862(N31356,N31361,N31362);
and and18863(N31357,N31363,R4);
and and18868(N31368,N31372,N31373);
and and18869(N31369,N31374,R0);
and and18870(N31370,N31375,N31376);
and and18871(N31371,N31377,N31378);
and and18876(N31382,N31386,N31387);
and and18877(N31383,N31388,R0);
and and18878(N31384,R1,N31389);
and and18879(N31385,N31390,R5);
and and18884(N31396,N31400,N31401);
and and18885(N31397,N31402,R1);
and and18886(N31398,R2,N31403);
and and18887(N31399,R4,R5);
and and18892(N31409,N31413,N31414);
and and18893(N31410,in2,R0);
and and18894(N31411,N31415,N31416);
and and18895(N31412,R3,N31417);
and and18900(N31422,N31426,N31427);
and and18901(N31423,N31428,R1);
and and18902(N31424,R2,R3);
and and18903(N31425,N31429,R5);
and and18908(N31435,N31439,N31440);
and and18909(N31436,N31441,N31442);
and and18910(N31437,N31443,R2);
and and18911(N31438,R3,R4);
and and18916(N31448,N31452,N31453);
and and18917(N31449,N31454,N31455);
and and18918(N31450,N31456,R2);
and and18919(N31451,N31457,R5);
and and18924(N31461,N31465,N31466);
and and18925(N31462,N31467,R1);
and and18926(N31463,R2,R3);
and and18927(N31464,N31468,R5);
and and18932(N31474,N31478,N31479);
and and18933(N31475,N31480,N31481);
and and18934(N31476,R1,R2);
and and18935(N31477,N31482,R4);
and and18940(N31487,N31491,N31492);
and and18941(N31488,in2,R0);
and and18942(N31489,N31493,R2);
and and18943(N31490,N31494,N31495);
and and18948(N31499,N31503,N31504);
and and18949(N31500,in1,in2);
and and18950(N31501,R0,N31505);
and and18951(N31502,N31506,N31507);
and and18956(N31511,N31515,N31516);
and and18957(N31512,N31517,R0);
and and18958(N31513,R1,N31518);
and and18959(N31514,R3,N31519);
and and18964(N31523,N31527,N31528);
and and18965(N31524,in1,in2);
and and18966(N31525,R0,R1);
and and18967(N31526,N31529,R3);
and and18972(N31535,N31539,N31540);
and and18973(N31536,in1,in2);
and and18974(N31537,R0,R2);
and and18975(N31538,N31541,N31542);
and and18980(N31546,N31550,N31551);
and and18981(N31547,in1,in2);
and and18982(N31548,N31552,R2);
and and18983(N31549,R3,R4);
and and18988(N31557,N31561,N31562);
and and18989(N31558,in2,R0);
and and18990(N31559,R1,R3);
and and18991(N31560,N31563,R5);
and and17528(N29223,N29229,R3);
and and17529(N29224,N29230,N29231);
and and17530(N29225,N29232,N29233);
and and17538(N29241,R2,N29249);
and and17539(N29242,R4,N29250);
and and17540(N29243,R6,N29251);
and and17548(N29259,N29264,R3);
and and17549(N29260,R4,N29265);
and and17550(N29261,N29266,R7);
and and17558(N29274,N29281,N29282);
and and17559(N29275,N29283,N29284);
and and17567(N29292,N29299,N29300);
and and17568(N29293,N29301,N29302);
and and17576(N29310,N29317,N29318);
and and17577(N29311,N29319,N29320);
and and17585(N29328,N29336,R5);
and and17586(N29329,N29337,N29338);
and and17594(N29346,N29353,N29354);
and and17595(N29347,N29355,N29356);
and and17603(N29364,N29371,N29372);
and and17604(N29365,N29373,R7);
and and17612(N29381,R4,N29388);
and and17613(N29382,N29389,N29390);
and and17621(N29398,R4,N29405);
and and17622(N29399,N29406,N29407);
and and17630(N29415,N29421,N29422);
and and17631(N29416,N29423,N29424);
and and17639(N29432,N29438,N29439);
and and17640(N29433,N29440,N29441);
and and17648(N29449,N29456,R5);
and and17649(N29450,N29457,N29458);
and and17657(N29466,N29473,N29474);
and and17658(N29467,N29475,R7);
and and17666(N29483,N29490,N29491);
and and17667(N29484,N29492,R7);
and and17675(N29500,R3,R5);
and and17676(N29501,N29508,N29509);
and and17684(N29517,N29524,N29525);
and and17685(N29518,N29526,R7);
and and17693(N29534,N29539,N29540);
and and17694(N29535,N29541,N29542);
and and17702(N29550,N29556,R5);
and and17703(N29551,N29557,N29558);
and and17711(N29566,N29571,N29572);
and and17712(N29567,N29573,N29574);
and and17720(N29582,N29587,N29588);
and and17721(N29583,N29589,N29590);
and and17729(N29598,N29604,N29605);
and and17730(N29599,N29606,R7);
and and17738(N29614,N29620,N29621);
and and17739(N29615,R5,N29622);
and and17747(N29630,R4,N29636);
and and17748(N29631,N29637,N29638);
and and17756(N29646,R3,N29653);
and and17757(N29647,N29654,R7);
and and17765(N29662,R4,N29668);
and and17766(N29663,N29669,N29670);
and and17774(N29678,R4,N29685);
and and17775(N29679,R6,N29686);
and and17783(N29694,N29700,R5);
and and17784(N29695,N29701,N29702);
and and17792(N29710,N29716,N29717);
and and17793(N29711,N29718,R7);
and and17801(N29726,R4,N29732);
and and17802(N29727,N29733,N29734);
and and17810(N29742,R3,N29749);
and and17811(N29743,N29750,R6);
and and17819(N29758,R3,N29765);
and and17820(N29759,R5,R7);
and and17828(N29773,R4,R5);
and and17829(N29774,N29780,R7);
and and17837(N29788,R4,R5);
and and17838(N29789,N29794,N29795);
and and17846(N29803,N29807,N29808);
and and17847(N29804,N29809,N29810);
and and17855(N29818,R3,N29824);
and and17856(N29819,R6,N29825);
and and17864(N29833,R4,R5);
and and17865(N29834,N29839,N29840);
and and17873(N29848,R3,R5);
and and17874(N29849,R6,R7);
and and17882(N29863,R3,N29869);
and and17883(N29864,N29870,R6);
and and17891(N29878,N29883,N29884);
and and17892(N29879,R5,N29885);
and and17900(N29893,N29898,R5);
and and17901(N29894,N29899,N29900);
and and17909(N29908,R4,N29914);
and and17910(N29909,R6,N29915);
and and17918(N29923,R4,N29928);
and and17919(N29924,N29929,N29930);
and and17927(N29938,N29943,R4);
and and17928(N29939,N29944,N29945);
and and17936(N29953,N29958,R5);
and and17937(N29954,N29959,N29960);
and and17945(N29968,R3,N29974);
and and17946(N29969,N29975,R6);
and and17954(N29983,N29988,N29989);
and and17955(N29984,R6,N29990);
and and17963(N29998,N30003,N30004);
and and17964(N29999,N30005,R7);
and and17972(N30013,N30019,R5);
and and17973(N30014,N30020,R7);
and and17981(N30028,N30033,R5);
and and17982(N30029,N30034,N30035);
and and17990(N30043,R4,N30048);
and and17991(N30044,N30049,N30050);
and and17999(N30058,R4,R5);
and and18000(N30059,N30064,N30065);
and and18008(N30073,N30078,R5);
and and18009(N30074,N30079,R7);
and and18017(N30087,N30092,R5);
and and18018(N30088,R6,N30093);
and and18026(N30101,N30106,N30107);
and and18027(N30102,R6,R7);
and and18035(N30115,N30120,N30121);
and and18036(N30116,R6,R7);
and and18044(N30129,N30133,N30134);
and and18045(N30130,R6,N30135);
and and18053(N30143,N30149,R4);
and and18054(N30144,R6,R7);
and and18062(N30157,N30161,N30162);
and and18063(N30158,N30163,R7);
and and18071(N30171,R3,R4);
and and18072(N30172,N30176,N30177);
and and18080(N30185,N30189,R5);
and and18081(N30186,N30190,N30191);
and and18089(N30199,N30203,N30204);
and and18090(N30200,N30205,R7);
and and18098(N30213,R4,N30218);
and and18099(N30214,R6,N30219);
and and18107(N30227,R4,N30232);
and and18108(N30228,R6,N30233);
and and18116(N30241,R3,N30247);
and and18117(N30242,R6,R7);
and and18125(N30255,N30260,R5);
and and18126(N30256,N30261,R7);
and and18134(N30269,R4,N30274);
and and18135(N30270,R6,N30275);
and and18143(N30283,R4,N30289);
and and18144(N30284,R6,R7);
and and18152(N30297,N30302,R5);
and and18153(N30298,R6,N30303);
and and18161(N30311,N30315,R4);
and and18162(N30312,N30316,N30317);
and and18170(N30325,R4,N30330);
and and18171(N30326,N30331,R7);
and and18179(N30339,N30344,R5);
and and18180(N30340,R6,N30345);
and and18188(N30353,N30358,R5);
and and18189(N30354,R6,N30359);
and and18197(N30367,R3,R4);
and and18198(N30368,R5,N30373);
and and18206(N30381,R4,N30385);
and and18207(N30382,N30386,N30387);
and and18215(N30395,R4,R5);
and and18216(N30396,N30401,R7);
and and18224(N30409,N30414,N30415);
and and18225(N30410,R6,R7);
and and18233(N30423,R4,R5);
and and18234(N30424,R6,N30429);
and and18242(N30437,R4,R5);
and and18243(N30438,R6,R7);
and and18251(N30451,R3,R4);
and and18252(N30452,R5,R7);
and and18260(N30465,N30469,R4);
and and18261(N30466,N30470,N30471);
and and18269(N30479,R3,R4);
and and18270(N30480,N30484,N30485);
and and18278(N30493,N30498,N30499);
and and18279(N30494,R6,R7);
and and18287(N30507,R3,R4);
and and18288(N30508,N30513,R7);
and and18296(N30521,R4,R5);
and and18297(N30522,N30526,N30527);
and and18305(N30535,R3,N30540);
and and18306(N30536,N30541,R7);
and and18314(N30549,R3,R4);
and and18315(N30550,R5,R7);
and and18323(N30563,R4,R5);
and and18324(N30564,N30569,R7);
and and18332(N30577,R4,N30582);
and and18333(N30578,N30583,R7);
and and18341(N30591,N30596,R5);
and and18342(N30592,R6,N30597);
and and18350(N30605,R4,N30610);
and and18351(N30606,N30611,R7);
and and18359(N30619,N30624,R4);
and and18360(N30620,N30625,R7);
and and18368(N30633,R4,N30638);
and and18369(N30634,N30639,R7);
and and18377(N30647,R4,N30652);
and and18378(N30648,N30653,R7);
and and18386(N30661,N30665,N30666);
and and18387(N30662,N30667,R7);
and and18395(N30675,R3,R4);
and and18396(N30676,R6,N30681);
and and18404(N30689,N30693,N30694);
and and18405(N30690,R6,N30695);
and and18413(N30703,N30707,R4);
and and18414(N30704,N30708,N30709);
and and18422(N30717,R4,R5);
and and18423(N30718,N30721,N30722);
and and18431(N30730,R4,N30735);
and and18432(N30731,R6,R7);
and and18440(N30743,R4,N30747);
and and18441(N30744,N30748,R7);
and and18449(N30756,R3,N30761);
and and18450(N30757,R5,R7);
and and18458(N30769,N30773,N30774);
and and18459(N30770,R6,R7);
and and18467(N30782,N30787,R5);
and and18468(N30783,R6,R7);
and and18476(N30795,R3,R5);
and and18477(N30796,R6,R7);
and and18485(N30808,R3,R4);
and and18486(N30809,R6,N30813);
and and18494(N30821,R3,N30824);
and and18495(N30822,N30825,N30826);
and and18503(N30834,R4,R5);
and and18504(N30835,N30839,R7);
and and18512(N30847,R3,N30852);
and and18513(N30848,R5,R7);
and and18521(N30860,N30864,R5);
and and18522(N30861,N30865,R7);
and and18530(N30873,R4,R5);
and and18531(N30874,N30877,N30878);
and and18539(N30886,N30890,R5);
and and18540(N30887,N30891,R7);
and and18548(N30899,N30903,R4);
and and18549(N30900,R5,N30904);
and and18557(N30912,R3,N30916);
and and18558(N30913,R6,N30917);
and and18566(N30925,N30928,N30929);
and and18567(N30926,R6,N30930);
and and18575(N30938,R4,N30941);
and and18576(N30939,N30942,N30943);
and and18584(N30951,R4,R5);
and and18585(N30952,N30956,R7);
and and18593(N30964,N30968,R5);
and and18594(N30965,R6,N30969);
and and18602(N30977,R3,R5);
and and18603(N30978,N30982,R7);
and and18611(N30990,N30994,R4);
and and18612(N30991,R5,N30995);
and and18620(N31003,N31007,R4);
and and18621(N31004,R5,N31008);
and and18629(N31016,R4,N31020);
and and18630(N31017,N31021,R7);
and and18638(N31029,R4,R5);
and and18639(N31030,R6,N31033);
and and18647(N31041,R3,R5);
and and18648(N31042,R6,N31045);
and and18656(N31053,R4,R5);
and and18657(N31054,R6,R7);
and and18665(N31065,R3,R4);
and and18666(N31066,R5,R7);
and and18674(N31077,R4,N31081);
and and18675(N31078,R6,R7);
and and18683(N31089,R3,R4);
and and18684(N31090,N31093,R6);
and and18692(N31101,R4,R5);
and and18693(N31102,R6,R7);
and and18701(N31113,N31117,R5);
and and18702(N31114,R6,R7);
and and18710(N31125,R3,R4);
and and18711(N31126,N31129,R7);
and and18719(N31137,R4,R5);
and and18720(N31138,R6,R7);
and and18728(N31149,R3,R4);
and and18729(N31150,N31153,R6);
and and18737(N31161,R4,N31165);
and and18738(N31162,R6,R7);
and and18746(N31173,N31177,R5);
and and18747(N31174,R6,R7);
and and18755(N31185,R3,R5);
and and18756(N31186,R6,R7);
and and18764(N31197,R4,R5);
and and18765(N31198,R6,R7);
and and18773(N31209,R3,R4);
and and18774(N31210,R6,R7);
and and18782(N31220,R4,N31223);
and and18783(N31221,R6,R7);
and and18791(N31231,R3,R5);
and and18792(N31232,R6,R7);
and and18800(N31242,N31248,N31249);
and and18808(N31257,N31263,N31264);
and and18816(N31272,N31279,R7);
and and18824(N31287,N31293,N31294);
and and18832(N31302,N31308,R7);
and and18840(N31316,N31322,R5);
and and18848(N31330,N31336,R7);
and and18856(N31344,R5,R6);
and and18864(N31358,R5,N31364);
and and18872(N31372,R6,R7);
and and18880(N31386,N31391,N31392);
and and18888(N31400,N31404,N31405);
and and18896(N31413,R5,N31418);
and and18904(N31426,N31430,N31431);
and and18912(N31439,N31444,R7);
and and18920(N31452,R6,R7);
and and18928(N31465,N31469,N31470);
and and18936(N31478,R5,N31483);
and and18944(N31491,R5,R6);
and and18952(N31503,R5,R6);
and and18960(N31515,R6,R7);
and and18968(N31527,N31530,N31531);
and and18976(N31539,R6,R7);
and and18984(N31550,R6,N31553);
and and18992(N31561,R6,R7);
and and18993(N31784,N31785,N31786);
and and19003(N31799,N31800,N31801);
and and19012(N31817,N31818,N31819);
and and19021(N31835,N31836,N31837);
and and19030(N31853,N31854,N31855);
and and19039(N31871,N31872,N31873);
and and19048(N31889,N31890,N31891);
and and19057(N31907,N31908,N31909);
and and19066(N31925,N31926,N31927);
and and19075(N31942,N31943,N31944);
and and19084(N31959,N31960,N31961);
and and19093(N31976,N31977,N31978);
and and19102(N31993,N31994,N31995);
and and19111(N32010,N32011,N32012);
and and19120(N32027,N32028,N32029);
and and19129(N32043,N32044,N32045);
and and19138(N32059,N32060,N32061);
and and19147(N32075,N32076,N32077);
and and19156(N32091,N32092,N32093);
and and19165(N32107,N32108,N32109);
and and19174(N32123,N32124,N32125);
and and19183(N32139,N32140,N32141);
and and19192(N32155,N32156,N32157);
and and19201(N32171,N32172,N32173);
and and19210(N32187,N32188,N32189);
and and19219(N32203,N32204,N32205);
and and19228(N32219,N32220,N32221);
and and19237(N32235,N32236,N32237);
and and19246(N32251,N32252,N32253);
and and19255(N32267,N32268,N32269);
and and19264(N32283,N32284,N32285);
and and19273(N32299,N32300,N32301);
and and19282(N32315,N32316,N32317);
and and19291(N32331,N32332,N32333);
and and19300(N32347,N32348,N32349);
and and19309(N32363,N32364,N32365);
and and19318(N32379,N32380,N32381);
and and19327(N32395,N32396,N32397);
and and19336(N32411,N32412,N32413);
and and19345(N32427,N32428,N32429);
and and19354(N32442,N32443,N32444);
and and19363(N32457,N32458,N32459);
and and19372(N32472,N32473,N32474);
and and19381(N32487,N32488,N32489);
and and19390(N32502,N32503,N32504);
and and19399(N32517,N32518,N32519);
and and19408(N32532,N32533,N32534);
and and19417(N32547,N32548,N32549);
and and19426(N32562,N32563,N32564);
and and19435(N32577,N32578,N32579);
and and19444(N32592,N32593,N32594);
and and19453(N32607,N32608,N32609);
and and19462(N32622,N32623,N32624);
and and19471(N32637,N32638,N32639);
and and19480(N32652,N32653,N32654);
and and19489(N32667,N32668,N32669);
and and19498(N32682,N32683,N32684);
and and19507(N32697,N32698,N32699);
and and19516(N32712,N32713,N32714);
and and19525(N32727,N32728,N32729);
and and19534(N32742,N32743,N32744);
and and19543(N32757,N32758,N32759);
and and19552(N32772,N32773,N32774);
and and19561(N32787,N32788,N32789);
and and19570(N32802,N32803,N32804);
and and19579(N32817,N32818,N32819);
and and19588(N32831,N32832,N32833);
and and19597(N32845,N32846,N32847);
and and19606(N32859,N32860,N32861);
and and19615(N32873,N32874,N32875);
and and19624(N32887,N32888,N32889);
and and19633(N32901,N32902,N32903);
and and19642(N32915,N32916,N32917);
and and19651(N32929,N32930,N32931);
and and19660(N32943,N32944,N32945);
and and19669(N32957,N32958,N32959);
and and19678(N32971,N32972,N32973);
and and19687(N32985,N32986,N32987);
and and19696(N32999,N33000,N33001);
and and19705(N33013,N33014,N33015);
and and19714(N33027,N33028,N33029);
and and19723(N33041,N33042,N33043);
and and19732(N33055,N33056,N33057);
and and19741(N33069,N33070,N33071);
and and19750(N33083,N33084,N33085);
and and19759(N33097,N33098,N33099);
and and19768(N33111,N33112,N33113);
and and19777(N33125,N33126,N33127);
and and19786(N33139,N33140,N33141);
and and19795(N33153,N33154,N33155);
and and19804(N33167,N33168,N33169);
and and19813(N33181,N33182,N33183);
and and19822(N33195,N33196,N33197);
and and19831(N33209,N33210,N33211);
and and19840(N33223,N33224,N33225);
and and19849(N33237,N33238,N33239);
and and19858(N33251,N33252,N33253);
and and19867(N33265,N33266,N33267);
and and19876(N33279,N33280,N33281);
and and19885(N33293,N33294,N33295);
and and19894(N33307,N33308,N33309);
and and19903(N33321,N33322,N33323);
and and19912(N33335,N33336,N33337);
and and19921(N33349,N33350,N33351);
and and19930(N33363,N33364,N33365);
and and19939(N33377,N33378,N33379);
and and19948(N33391,N33392,N33393);
and and19957(N33405,N33406,N33407);
and and19966(N33418,N33419,N33420);
and and19975(N33431,N33432,N33433);
and and19984(N33444,N33445,N33446);
and and19993(N33457,N33458,N33459);
and and20002(N33470,N33471,N33472);
and and20011(N33483,N33484,N33485);
and and20020(N33496,N33497,N33498);
and and20029(N33509,N33510,N33511);
and and20038(N33522,N33523,N33524);
and and20047(N33535,N33536,N33537);
and and20056(N33548,N33549,N33550);
and and20065(N33561,N33562,N33563);
and and20074(N33574,N33575,N33576);
and and20083(N33587,N33588,N33589);
and and20092(N33600,N33601,N33602);
and and20101(N33613,N33614,N33615);
and and20110(N33626,N33627,N33628);
and and20119(N33639,N33640,N33641);
and and20128(N33652,N33653,N33654);
and and20137(N33665,N33666,N33667);
and and20146(N33678,N33679,N33680);
and and20155(N33691,N33692,N33693);
and and20164(N33704,N33705,N33706);
and and20173(N33717,N33718,N33719);
and and20182(N33729,N33730,N33731);
and and20191(N33741,N33742,N33743);
and and20200(N33753,N33754,N33755);
and and20209(N33765,N33766,N33767);
and and20218(N33777,N33778,N33779);
and and20227(N33789,N33790,N33791);
and and20236(N33801,N33802,N33803);
and and20245(N33813,N33814,N33815);
and and20254(N33825,N33826,N33827);
and and20263(N33837,N33838,N33839);
and and20272(N33849,N33850,N33851);
and and20281(N33861,N33862,N33863);
and and20290(N33873,N33874,N33875);
and and20299(N33885,N33886,N33887);
and and20308(N33897,N33898,N33899);
and and20317(N33909,N33910,N33911);
and and20326(N33921,N33922,N33923);
and and20335(N33933,N33934,N33935);
and and20344(N33945,N33946,N33947);
and and20353(N33957,N33958,N33959);
and and20362(N33969,N33970,N33971);
and and20371(N33980,N33981,N33982);
and and20380(N33991,N33992,N33993);
and and20389(N34002,N34003,N34004);
and and20398(N34013,N34014,N34015);
and and20407(N34024,N34025,N34026);
and and20416(N34035,N34036,N34037);
and and20425(N34045,N34046,N34047);
and and20433(N34061,N34062,N34063);
and and20441(N34076,N34077,N34078);
and and20449(N34091,N34092,N34093);
and and20457(N34106,N34107,N34108);
and and20465(N34120,N34121,N34122);
and and20473(N34134,N34135,N34136);
and and20481(N34148,N34149,N34150);
and and20489(N34162,N34163,N34164);
and and20497(N34176,N34177,N34178);
and and20505(N34190,N34191,N34192);
and and20513(N34204,N34205,N34206);
and and20521(N34218,N34219,N34220);
and and20529(N34232,N34233,N34234);
and and20537(N34246,N34247,N34248);
and and20545(N34260,N34261,N34262);
and and20553(N34274,N34275,N34276);
and and20561(N34288,N34289,N34290);
and and20569(N34302,N34303,N34304);
and and20577(N34316,N34317,N34318);
and and20585(N34329,N34330,N34331);
and and20593(N34342,N34343,N34344);
and and20601(N34355,N34356,N34357);
and and20609(N34368,N34369,N34370);
and and20617(N34381,N34382,N34383);
and and20625(N34394,N34395,N34396);
and and20633(N34407,N34408,N34409);
and and20641(N34420,N34421,N34422);
and and20649(N34433,N34434,N34435);
and and20657(N34445,N34446,N34447);
and and20665(N34457,N34458,N34459);
and and20673(N34469,N34470,N34471);
and and20681(N34481,N34482,N34483);
and and20689(N34493,N34494,N34495);
and and20697(N34505,N34506,N34507);
and and20705(N34517,N34518,N34519);
and and20713(N34529,N34530,N34531);
and and20721(N34541,N34542,N34543);
and and20729(N34553,N34554,N34555);
and and20737(N34565,N34566,N34567);
and and20745(N34577,N34578,N34579);
and and20753(N34589,N34590,N34591);
and and20761(N34601,N34602,N34603);
and and20769(N34613,N34614,N34615);
and and20777(N34625,N34626,N34627);
and and20785(N34637,N34638,N34639);
and and20793(N34649,N34650,N34651);
and and20801(N34661,N34662,N34663);
and and20809(N34673,N34674,N34675);
and and20817(N34685,N34686,N34687);
and and20825(N34697,N34698,N34699);
and and20833(N34708,N34709,N34710);
and and20841(N34719,N34720,N34721);
and and20849(N34730,N34731,N34732);
and and20857(N34741,N34742,N34743);
and and20865(N34752,N34753,N34754);
and and20873(N34762,N34763,N34764);
and and20881(N34772,N34773,N34774);
and and20889(N34782,N34783,N34784);
and and20897(N34791,N34792,N34793);
and and20904(N34802,N34803,N34804);
and and20911(N34813,N34814,N34815);
and and18994(N31785,N31787,N31788);
and and18995(N31786,N31789,N31790);
and and19004(N31800,N31802,N31803);
and and19005(N31801,N31804,N31805);
and and19013(N31818,N31820,N31821);
and and19014(N31819,N31822,N31823);
and and19022(N31836,N31838,N31839);
and and19023(N31837,N31840,N31841);
and and19031(N31854,N31856,N31857);
and and19032(N31855,N31858,N31859);
and and19040(N31872,N31874,N31875);
and and19041(N31873,N31876,N31877);
and and19049(N31890,N31892,N31893);
and and19050(N31891,N31894,N31895);
and and19058(N31908,N31910,N31911);
and and19059(N31909,N31912,N31913);
and and19067(N31926,N31928,N31929);
and and19068(N31927,N31930,N31931);
and and19076(N31943,N31945,N31946);
and and19077(N31944,N31947,N31948);
and and19085(N31960,N31962,N31963);
and and19086(N31961,N31964,N31965);
and and19094(N31977,N31979,N31980);
and and19095(N31978,N31981,N31982);
and and19103(N31994,N31996,N31997);
and and19104(N31995,N31998,N31999);
and and19112(N32011,N32013,N32014);
and and19113(N32012,N32015,N32016);
and and19121(N32028,N32030,N32031);
and and19122(N32029,N32032,N32033);
and and19130(N32044,N32046,N32047);
and and19131(N32045,N32048,N32049);
and and19139(N32060,N32062,N32063);
and and19140(N32061,N32064,N32065);
and and19148(N32076,N32078,N32079);
and and19149(N32077,N32080,N32081);
and and19157(N32092,N32094,N32095);
and and19158(N32093,N32096,N32097);
and and19166(N32108,N32110,N32111);
and and19167(N32109,N32112,N32113);
and and19175(N32124,N32126,N32127);
and and19176(N32125,N32128,N32129);
and and19184(N32140,N32142,N32143);
and and19185(N32141,N32144,N32145);
and and19193(N32156,N32158,N32159);
and and19194(N32157,N32160,N32161);
and and19202(N32172,N32174,N32175);
and and19203(N32173,N32176,N32177);
and and19211(N32188,N32190,N32191);
and and19212(N32189,N32192,N32193);
and and19220(N32204,N32206,N32207);
and and19221(N32205,N32208,N32209);
and and19229(N32220,N32222,N32223);
and and19230(N32221,N32224,N32225);
and and19238(N32236,N32238,N32239);
and and19239(N32237,N32240,N32241);
and and19247(N32252,N32254,N32255);
and and19248(N32253,N32256,N32257);
and and19256(N32268,N32270,N32271);
and and19257(N32269,N32272,N32273);
and and19265(N32284,N32286,N32287);
and and19266(N32285,N32288,N32289);
and and19274(N32300,N32302,N32303);
and and19275(N32301,N32304,N32305);
and and19283(N32316,N32318,N32319);
and and19284(N32317,N32320,N32321);
and and19292(N32332,N32334,N32335);
and and19293(N32333,N32336,N32337);
and and19301(N32348,N32350,N32351);
and and19302(N32349,N32352,N32353);
and and19310(N32364,N32366,N32367);
and and19311(N32365,N32368,N32369);
and and19319(N32380,N32382,N32383);
and and19320(N32381,N32384,N32385);
and and19328(N32396,N32398,N32399);
and and19329(N32397,N32400,N32401);
and and19337(N32412,N32414,N32415);
and and19338(N32413,N32416,N32417);
and and19346(N32428,N32430,N32431);
and and19347(N32429,N32432,N32433);
and and19355(N32443,N32445,N32446);
and and19356(N32444,N32447,N32448);
and and19364(N32458,N32460,N32461);
and and19365(N32459,N32462,N32463);
and and19373(N32473,N32475,N32476);
and and19374(N32474,N32477,N32478);
and and19382(N32488,N32490,N32491);
and and19383(N32489,N32492,N32493);
and and19391(N32503,N32505,N32506);
and and19392(N32504,N32507,N32508);
and and19400(N32518,N32520,N32521);
and and19401(N32519,N32522,N32523);
and and19409(N32533,N32535,N32536);
and and19410(N32534,N32537,N32538);
and and19418(N32548,N32550,N32551);
and and19419(N32549,N32552,N32553);
and and19427(N32563,N32565,N32566);
and and19428(N32564,N32567,N32568);
and and19436(N32578,N32580,N32581);
and and19437(N32579,N32582,N32583);
and and19445(N32593,N32595,N32596);
and and19446(N32594,N32597,N32598);
and and19454(N32608,N32610,N32611);
and and19455(N32609,N32612,N32613);
and and19463(N32623,N32625,N32626);
and and19464(N32624,N32627,N32628);
and and19472(N32638,N32640,N32641);
and and19473(N32639,N32642,N32643);
and and19481(N32653,N32655,N32656);
and and19482(N32654,N32657,N32658);
and and19490(N32668,N32670,N32671);
and and19491(N32669,N32672,N32673);
and and19499(N32683,N32685,N32686);
and and19500(N32684,N32687,N32688);
and and19508(N32698,N32700,N32701);
and and19509(N32699,N32702,N32703);
and and19517(N32713,N32715,N32716);
and and19518(N32714,N32717,N32718);
and and19526(N32728,N32730,N32731);
and and19527(N32729,N32732,N32733);
and and19535(N32743,N32745,N32746);
and and19536(N32744,N32747,N32748);
and and19544(N32758,N32760,N32761);
and and19545(N32759,N32762,N32763);
and and19553(N32773,N32775,N32776);
and and19554(N32774,N32777,N32778);
and and19562(N32788,N32790,N32791);
and and19563(N32789,N32792,N32793);
and and19571(N32803,N32805,N32806);
and and19572(N32804,N32807,N32808);
and and19580(N32818,N32820,N32821);
and and19581(N32819,N32822,N32823);
and and19589(N32832,N32834,N32835);
and and19590(N32833,N32836,N32837);
and and19598(N32846,N32848,N32849);
and and19599(N32847,N32850,N32851);
and and19607(N32860,N32862,N32863);
and and19608(N32861,N32864,N32865);
and and19616(N32874,N32876,N32877);
and and19617(N32875,N32878,N32879);
and and19625(N32888,N32890,N32891);
and and19626(N32889,N32892,N32893);
and and19634(N32902,N32904,N32905);
and and19635(N32903,N32906,N32907);
and and19643(N32916,N32918,N32919);
and and19644(N32917,N32920,N32921);
and and19652(N32930,N32932,N32933);
and and19653(N32931,N32934,N32935);
and and19661(N32944,N32946,N32947);
and and19662(N32945,N32948,N32949);
and and19670(N32958,N32960,N32961);
and and19671(N32959,N32962,N32963);
and and19679(N32972,N32974,N32975);
and and19680(N32973,N32976,N32977);
and and19688(N32986,N32988,N32989);
and and19689(N32987,N32990,N32991);
and and19697(N33000,N33002,N33003);
and and19698(N33001,N33004,N33005);
and and19706(N33014,N33016,N33017);
and and19707(N33015,N33018,N33019);
and and19715(N33028,N33030,N33031);
and and19716(N33029,N33032,N33033);
and and19724(N33042,N33044,N33045);
and and19725(N33043,N33046,N33047);
and and19733(N33056,N33058,N33059);
and and19734(N33057,N33060,N33061);
and and19742(N33070,N33072,N33073);
and and19743(N33071,N33074,N33075);
and and19751(N33084,N33086,N33087);
and and19752(N33085,N33088,N33089);
and and19760(N33098,N33100,N33101);
and and19761(N33099,N33102,N33103);
and and19769(N33112,N33114,N33115);
and and19770(N33113,N33116,N33117);
and and19778(N33126,N33128,N33129);
and and19779(N33127,N33130,N33131);
and and19787(N33140,N33142,N33143);
and and19788(N33141,N33144,N33145);
and and19796(N33154,N33156,N33157);
and and19797(N33155,N33158,N33159);
and and19805(N33168,N33170,N33171);
and and19806(N33169,N33172,N33173);
and and19814(N33182,N33184,N33185);
and and19815(N33183,N33186,N33187);
and and19823(N33196,N33198,N33199);
and and19824(N33197,N33200,N33201);
and and19832(N33210,N33212,N33213);
and and19833(N33211,N33214,N33215);
and and19841(N33224,N33226,N33227);
and and19842(N33225,N33228,N33229);
and and19850(N33238,N33240,N33241);
and and19851(N33239,N33242,N33243);
and and19859(N33252,N33254,N33255);
and and19860(N33253,N33256,N33257);
and and19868(N33266,N33268,N33269);
and and19869(N33267,N33270,N33271);
and and19877(N33280,N33282,N33283);
and and19878(N33281,N33284,N33285);
and and19886(N33294,N33296,N33297);
and and19887(N33295,N33298,N33299);
and and19895(N33308,N33310,N33311);
and and19896(N33309,N33312,N33313);
and and19904(N33322,N33324,N33325);
and and19905(N33323,N33326,N33327);
and and19913(N33336,N33338,N33339);
and and19914(N33337,N33340,N33341);
and and19922(N33350,N33352,N33353);
and and19923(N33351,N33354,N33355);
and and19931(N33364,N33366,N33367);
and and19932(N33365,N33368,N33369);
and and19940(N33378,N33380,N33381);
and and19941(N33379,N33382,N33383);
and and19949(N33392,N33394,N33395);
and and19950(N33393,N33396,N33397);
and and19958(N33406,N33408,N33409);
and and19959(N33407,N33410,N33411);
and and19967(N33419,N33421,N33422);
and and19968(N33420,N33423,N33424);
and and19976(N33432,N33434,N33435);
and and19977(N33433,N33436,N33437);
and and19985(N33445,N33447,N33448);
and and19986(N33446,N33449,N33450);
and and19994(N33458,N33460,N33461);
and and19995(N33459,N33462,N33463);
and and20003(N33471,N33473,N33474);
and and20004(N33472,N33475,N33476);
and and20012(N33484,N33486,N33487);
and and20013(N33485,N33488,N33489);
and and20021(N33497,N33499,N33500);
and and20022(N33498,N33501,N33502);
and and20030(N33510,N33512,N33513);
and and20031(N33511,N33514,N33515);
and and20039(N33523,N33525,N33526);
and and20040(N33524,N33527,N33528);
and and20048(N33536,N33538,N33539);
and and20049(N33537,N33540,N33541);
and and20057(N33549,N33551,N33552);
and and20058(N33550,N33553,N33554);
and and20066(N33562,N33564,N33565);
and and20067(N33563,N33566,N33567);
and and20075(N33575,N33577,N33578);
and and20076(N33576,N33579,N33580);
and and20084(N33588,N33590,N33591);
and and20085(N33589,N33592,N33593);
and and20093(N33601,N33603,N33604);
and and20094(N33602,N33605,N33606);
and and20102(N33614,N33616,N33617);
and and20103(N33615,N33618,N33619);
and and20111(N33627,N33629,N33630);
and and20112(N33628,N33631,N33632);
and and20120(N33640,N33642,N33643);
and and20121(N33641,N33644,N33645);
and and20129(N33653,N33655,N33656);
and and20130(N33654,N33657,N33658);
and and20138(N33666,N33668,N33669);
and and20139(N33667,N33670,N33671);
and and20147(N33679,N33681,N33682);
and and20148(N33680,N33683,N33684);
and and20156(N33692,N33694,N33695);
and and20157(N33693,N33696,N33697);
and and20165(N33705,N33707,N33708);
and and20166(N33706,N33709,N33710);
and and20174(N33718,N33720,N33721);
and and20175(N33719,N33722,N33723);
and and20183(N33730,N33732,N33733);
and and20184(N33731,N33734,N33735);
and and20192(N33742,N33744,N33745);
and and20193(N33743,N33746,N33747);
and and20201(N33754,N33756,N33757);
and and20202(N33755,N33758,N33759);
and and20210(N33766,N33768,N33769);
and and20211(N33767,N33770,N33771);
and and20219(N33778,N33780,N33781);
and and20220(N33779,N33782,N33783);
and and20228(N33790,N33792,N33793);
and and20229(N33791,N33794,N33795);
and and20237(N33802,N33804,N33805);
and and20238(N33803,N33806,N33807);
and and20246(N33814,N33816,N33817);
and and20247(N33815,N33818,N33819);
and and20255(N33826,N33828,N33829);
and and20256(N33827,N33830,N33831);
and and20264(N33838,N33840,N33841);
and and20265(N33839,N33842,N33843);
and and20273(N33850,N33852,N33853);
and and20274(N33851,N33854,N33855);
and and20282(N33862,N33864,N33865);
and and20283(N33863,N33866,N33867);
and and20291(N33874,N33876,N33877);
and and20292(N33875,N33878,N33879);
and and20300(N33886,N33888,N33889);
and and20301(N33887,N33890,N33891);
and and20309(N33898,N33900,N33901);
and and20310(N33899,N33902,N33903);
and and20318(N33910,N33912,N33913);
and and20319(N33911,N33914,N33915);
and and20327(N33922,N33924,N33925);
and and20328(N33923,N33926,N33927);
and and20336(N33934,N33936,N33937);
and and20337(N33935,N33938,N33939);
and and20345(N33946,N33948,N33949);
and and20346(N33947,N33950,N33951);
and and20354(N33958,N33960,N33961);
and and20355(N33959,N33962,N33963);
and and20363(N33970,N33972,N33973);
and and20364(N33971,N33974,N33975);
and and20372(N33981,N33983,N33984);
and and20373(N33982,N33985,N33986);
and and20381(N33992,N33994,N33995);
and and20382(N33993,N33996,N33997);
and and20390(N34003,N34005,N34006);
and and20391(N34004,N34007,N34008);
and and20399(N34014,N34016,N34017);
and and20400(N34015,N34018,N34019);
and and20408(N34025,N34027,N34028);
and and20409(N34026,N34029,N34030);
and and20417(N34036,N34038,N34039);
and and20418(N34037,N34040,N34041);
and and20426(N34046,N34048,N34049);
and and20427(N34047,N34050,N34051);
and and20434(N34062,N34064,N34065);
and and20435(N34063,N34066,N34067);
and and20442(N34077,N34079,N34080);
and and20443(N34078,N34081,N34082);
and and20450(N34092,N34094,N34095);
and and20451(N34093,N34096,N34097);
and and20458(N34107,N34109,N34110);
and and20459(N34108,N34111,N34112);
and and20466(N34121,N34123,N34124);
and and20467(N34122,N34125,N34126);
and and20474(N34135,N34137,N34138);
and and20475(N34136,N34139,N34140);
and and20482(N34149,N34151,N34152);
and and20483(N34150,N34153,N34154);
and and20490(N34163,N34165,N34166);
and and20491(N34164,N34167,N34168);
and and20498(N34177,N34179,N34180);
and and20499(N34178,N34181,N34182);
and and20506(N34191,N34193,N34194);
and and20507(N34192,N34195,N34196);
and and20514(N34205,N34207,N34208);
and and20515(N34206,N34209,N34210);
and and20522(N34219,N34221,N34222);
and and20523(N34220,N34223,N34224);
and and20530(N34233,N34235,N34236);
and and20531(N34234,N34237,N34238);
and and20538(N34247,N34249,N34250);
and and20539(N34248,N34251,N34252);
and and20546(N34261,N34263,N34264);
and and20547(N34262,N34265,N34266);
and and20554(N34275,N34277,N34278);
and and20555(N34276,N34279,N34280);
and and20562(N34289,N34291,N34292);
and and20563(N34290,N34293,N34294);
and and20570(N34303,N34305,N34306);
and and20571(N34304,N34307,N34308);
and and20578(N34317,N34319,N34320);
and and20579(N34318,N34321,N34322);
and and20586(N34330,N34332,N34333);
and and20587(N34331,N34334,N34335);
and and20594(N34343,N34345,N34346);
and and20595(N34344,N34347,N34348);
and and20602(N34356,N34358,N34359);
and and20603(N34357,N34360,N34361);
and and20610(N34369,N34371,N34372);
and and20611(N34370,N34373,N34374);
and and20618(N34382,N34384,N34385);
and and20619(N34383,N34386,N34387);
and and20626(N34395,N34397,N34398);
and and20627(N34396,N34399,N34400);
and and20634(N34408,N34410,N34411);
and and20635(N34409,N34412,N34413);
and and20642(N34421,N34423,N34424);
and and20643(N34422,N34425,N34426);
and and20650(N34434,N34436,N34437);
and and20651(N34435,N34438,N34439);
and and20658(N34446,N34448,N34449);
and and20659(N34447,N34450,N34451);
and and20666(N34458,N34460,N34461);
and and20667(N34459,N34462,N34463);
and and20674(N34470,N34472,N34473);
and and20675(N34471,N34474,N34475);
and and20682(N34482,N34484,N34485);
and and20683(N34483,N34486,N34487);
and and20690(N34494,N34496,N34497);
and and20691(N34495,N34498,N34499);
and and20698(N34506,N34508,N34509);
and and20699(N34507,N34510,N34511);
and and20706(N34518,N34520,N34521);
and and20707(N34519,N34522,N34523);
and and20714(N34530,N34532,N34533);
and and20715(N34531,N34534,N34535);
and and20722(N34542,N34544,N34545);
and and20723(N34543,N34546,N34547);
and and20730(N34554,N34556,N34557);
and and20731(N34555,N34558,N34559);
and and20738(N34566,N34568,N34569);
and and20739(N34567,N34570,N34571);
and and20746(N34578,N34580,N34581);
and and20747(N34579,N34582,N34583);
and and20754(N34590,N34592,N34593);
and and20755(N34591,N34594,N34595);
and and20762(N34602,N34604,N34605);
and and20763(N34603,N34606,N34607);
and and20770(N34614,N34616,N34617);
and and20771(N34615,N34618,N34619);
and and20778(N34626,N34628,N34629);
and and20779(N34627,N34630,N34631);
and and20786(N34638,N34640,N34641);
and and20787(N34639,N34642,N34643);
and and20794(N34650,N34652,N34653);
and and20795(N34651,N34654,N34655);
and and20802(N34662,N34664,N34665);
and and20803(N34663,N34666,N34667);
and and20810(N34674,N34676,N34677);
and and20811(N34675,N34678,N34679);
and and20818(N34686,N34688,N34689);
and and20819(N34687,N34690,N34691);
and and20826(N34698,N34700,N34701);
and and20827(N34699,N34702,N34703);
and and20834(N34709,N34711,N34712);
and and20835(N34710,N34713,N34714);
and and20842(N34720,N34722,N34723);
and and20843(N34721,N34724,N34725);
and and20850(N34731,N34733,N34734);
and and20851(N34732,N34735,N34736);
and and20858(N34742,N34744,N34745);
and and20859(N34743,N34746,N34747);
and and20866(N34753,N34755,N34756);
and and20867(N34754,N34757,N34758);
and and20874(N34763,N34765,N34766);
and and20875(N34764,N34767,N34768);
and and20882(N34773,N34775,N34776);
and and20883(N34774,N34777,N34778);
and and20890(N34783,N34785,N34786);
and and20891(N34784,N34787,N34788);
and and20898(N34792,N34794,N34795);
and and20899(N34793,N34796,N34797);
and and20905(N34803,N34805,N34806);
and and20906(N34804,N34807,N34808);
and and20912(N34814,N34816,N34817);
and and20913(N34815,N34818,N34819);
and and18996(N31787,N31791,N31792);
and and18997(N31788,N31793,N31794);
and and18998(N31789,in1,in2);
and and18999(N31790,N31795,R1);
and and19006(N31802,N31806,N31807);
and and19007(N31803,N31808,N31809);
and and19008(N31804,N31810,N31811);
and and19009(N31805,R1,N31812);
and and19015(N31820,N31824,N31825);
and and19016(N31821,N31826,N31827);
and and19017(N31822,N31828,N31829);
and and19018(N31823,N31830,N31831);
and and19024(N31838,N31842,N31843);
and and19025(N31839,N31844,in1);
and and19026(N31840,N31845,N31846);
and and19027(N31841,N31847,N31848);
and and19033(N31856,N31860,N31861);
and and19034(N31857,N31862,N31863);
and and19035(N31858,N31864,N31865);
and and19036(N31859,N31866,R2);
and and19042(N31874,N31878,N31879);
and and19043(N31875,N31880,N31881);
and and19044(N31876,N31882,N31883);
and and19045(N31877,N31884,N31885);
and and19051(N31892,N31896,N31897);
and and19052(N31893,N31898,N31899);
and and19053(N31894,N31900,N31901);
and and19054(N31895,N31902,R3);
and and19060(N31910,N31914,N31915);
and and19061(N31911,N31916,N31917);
and and19062(N31912,N31918,N31919);
and and19063(N31913,N31920,N31921);
and and19069(N31928,N31932,N31933);
and and19070(N31929,N31934,in2);
and and19071(N31930,R0,N31935);
and and19072(N31931,N31936,N31937);
and and19078(N31945,N31949,N31950);
and and19079(N31946,N31951,N31952);
and and19080(N31947,in2,N31953);
and and19081(N31948,N31954,N31955);
and and19087(N31962,N31966,N31967);
and and19088(N31963,N31968,N31969);
and and19089(N31964,N31970,N31971);
and and19090(N31965,N31972,N31973);
and and19096(N31979,N31983,N31984);
and and19097(N31980,N31985,N31986);
and and19098(N31981,R0,N31987);
and and19099(N31982,N31988,N31989);
and and19105(N31996,N32000,N32001);
and and19106(N31997,N32002,N32003);
and and19107(N31998,N32004,N32005);
and and19108(N31999,N32006,N32007);
and and19114(N32013,N32017,N32018);
and and19115(N32014,N32019,N32020);
and and19116(N32015,N32021,N32022);
and and19117(N32016,N32023,N32024);
and and19123(N32030,N32034,N32035);
and and19124(N32031,N32036,in1);
and and19125(N32032,in2,R1);
and and19126(N32033,N32037,N32038);
and and19132(N32046,N32050,N32051);
and and19133(N32047,in0,in2);
and and19134(N32048,N32052,N32053);
and and19135(N32049,N32054,N32055);
and and19141(N32062,N32066,N32067);
and and19142(N32063,in0,in1);
and and19143(N32064,N32068,N32069);
and and19144(N32065,N32070,N32071);
and and19150(N32078,N32082,N32083);
and and19151(N32079,N32084,N32085);
and and19152(N32080,in2,R0);
and and19153(N32081,N32086,N32087);
and and19159(N32094,N32098,N32099);
and and19160(N32095,N32100,N32101);
and and19161(N32096,in2,R0);
and and19162(N32097,N32102,N32103);
and and19168(N32110,N32114,N32115);
and and19169(N32111,N32116,N32117);
and and19170(N32112,N32118,R1);
and and19171(N32113,N32119,R3);
and and19177(N32126,N32130,N32131);
and and19178(N32127,N32132,in1);
and and19179(N32128,N32133,N32134);
and and19180(N32129,R2,N32135);
and and19186(N32142,N32146,N32147);
and and19187(N32143,N32148,N32149);
and and19188(N32144,N32150,N32151);
and and19189(N32145,R1,R2);
and and19195(N32158,N32162,N32163);
and and19196(N32159,N32164,N32165);
and and19197(N32160,N32166,N32167);
and and19198(N32161,N32168,R3);
and and19204(N32174,N32178,N32179);
and and19205(N32175,N32180,N32181);
and and19206(N32176,R0,R1);
and and19207(N32177,N32182,N32183);
and and19213(N32190,N32194,N32195);
and and19214(N32191,N32196,in1);
and and19215(N32192,N32197,R0);
and and19216(N32193,N32198,N32199);
and and19222(N32206,N32210,N32211);
and and19223(N32207,N32212,N32213);
and and19224(N32208,N32214,R0);
and and19225(N32209,N32215,R2);
and and19231(N32222,N32226,N32227);
and and19232(N32223,N32228,in1);
and and19233(N32224,N32229,N32230);
and and19234(N32225,R2,R3);
and and19240(N32238,N32242,N32243);
and and19241(N32239,N32244,N32245);
and and19242(N32240,in2,N32246);
and and19243(N32241,N32247,R2);
and and19249(N32254,N32258,N32259);
and and19250(N32255,N32260,in1);
and and19251(N32256,N32261,N32262);
and and19252(N32257,N32263,R2);
and and19258(N32270,N32274,N32275);
and and19259(N32271,N32276,in1);
and and19260(N32272,in2,N32277);
and and19261(N32273,N32278,N32279);
and and19267(N32286,N32290,N32291);
and and19268(N32287,N32292,in1);
and and19269(N32288,N32293,N32294);
and and19270(N32289,N32295,N32296);
and and19276(N32302,N32306,N32307);
and and19277(N32303,N32308,N32309);
and and19278(N32304,N32310,N32311);
and and19279(N32305,N32312,R3);
and and19285(N32318,N32322,N32323);
and and19286(N32319,N32324,in1);
and and19287(N32320,N32325,R0);
and and19288(N32321,N32326,N32327);
and and19294(N32334,N32338,N32339);
and and19295(N32335,N32340,N32341);
and and19296(N32336,N32342,R0);
and and19297(N32337,N32343,N32344);
and and19303(N32350,N32354,N32355);
and and19304(N32351,N32356,N32357);
and and19305(N32352,in2,N32358);
and and19306(N32353,N32359,R3);
and and19312(N32366,N32370,N32371);
and and19313(N32367,N32372,in1);
and and19314(N32368,N32373,N32374);
and and19315(N32369,N32375,R3);
and and19321(N32382,N32386,N32387);
and and19322(N32383,N32388,N32389);
and and19323(N32384,N32390,R0);
and and19324(N32385,N32391,R2);
and and19330(N32398,N32402,N32403);
and and19331(N32399,N32404,N32405);
and and19332(N32400,N32406,R0);
and and19333(N32401,R1,N32407);
and and19339(N32414,N32418,N32419);
and and19340(N32415,N32420,in1);
and and19341(N32416,N32421,N32422);
and and19342(N32417,N32423,N32424);
and and19348(N32430,N32434,N32435);
and and19349(N32431,N32436,N32437);
and and19350(N32432,R0,N32438);
and and19351(N32433,N32439,N32440);
and and19357(N32445,N32449,N32450);
and and19358(N32446,N32451,N32452);
and and19359(N32447,in2,R0);
and and19360(N32448,R1,R2);
and and19366(N32460,N32464,N32465);
and and19367(N32461,N32466,in2);
and and19368(N32462,N32467,R1);
and and19369(N32463,R2,R3);
and and19375(N32475,N32479,N32480);
and and19376(N32476,N32481,in1);
and and19377(N32477,in2,R0);
and and19378(N32478,N32482,R2);
and and19384(N32490,N32494,N32495);
and and19385(N32491,N32496,in1);
and and19386(N32492,N32497,R0);
and and19387(N32493,R1,N32498);
and and19393(N32505,N32509,N32510);
and and19394(N32506,N32511,in1);
and and19395(N32507,in2,R0);
and and19396(N32508,N32512,N32513);
and and19402(N32520,N32524,N32525);
and and19403(N32521,N32526,in2);
and and19404(N32522,R0,N32527);
and and19405(N32523,N32528,N32529);
and and19411(N32535,N32539,N32540);
and and19412(N32536,N32541,N32542);
and and19413(N32537,N32543,R1);
and and19414(N32538,N32544,R3);
and and19420(N32550,N32554,N32555);
and and19421(N32551,N32556,N32557);
and and19422(N32552,in2,R0);
and and19423(N32553,N32558,R3);
and and19429(N32565,N32569,N32570);
and and19430(N32566,N32571,in1);
and and19431(N32567,in2,N32572);
and and19432(N32568,N32573,R3);
and and19438(N32580,N32584,N32585);
and and19439(N32581,N32586,in1);
and and19440(N32582,in2,N32587);
and and19441(N32583,N32588,N32589);
and and19447(N32595,N32599,N32600);
and and19448(N32596,N32601,in2);
and and19449(N32597,R0,R1);
and and19450(N32598,N32602,N32603);
and and19456(N32610,N32614,N32615);
and and19457(N32611,N32616,N32617);
and and19458(N32612,N32618,N32619);
and and19459(N32613,R1,R2);
and and19465(N32625,N32629,N32630);
and and19466(N32626,N32631,in1);
and and19467(N32627,N32632,N32633);
and and19468(N32628,R2,N32634);
and and19474(N32640,N32644,N32645);
and and19475(N32641,N32646,N32647);
and and19476(N32642,in2,N32648);
and and19477(N32643,N32649,R2);
and and19483(N32655,N32659,N32660);
and and19484(N32656,N32661,N32662);
and and19485(N32657,N32663,N32664);
and and19486(N32658,N32665,N32666);
and and19492(N32670,N32674,N32675);
and and19493(N32671,N32676,in1);
and and19494(N32672,N32677,R0);
and and19495(N32673,N32678,R2);
and and19501(N32685,N32689,N32690);
and and19502(N32686,N32691,N32692);
and and19503(N32687,in2,R0);
and and19504(N32688,N32693,N32694);
and and19510(N32700,N32704,N32705);
and and19511(N32701,N32706,in1);
and and19512(N32702,N32707,R0);
and and19513(N32703,R1,N32708);
and and19519(N32715,N32719,N32720);
and and19520(N32716,N32721,in2);
and and19521(N32717,R0,R1);
and and19522(N32718,N32722,R3);
and and19528(N32730,N32734,N32735);
and and19529(N32731,N32736,N32737);
and and19530(N32732,N32738,N32739);
and and19531(N32733,N32740,R2);
and and19537(N32745,N32749,N32750);
and and19538(N32746,N32751,N32752);
and and19539(N32747,N32753,R1);
and and19540(N32748,N32754,R3);
and and19546(N32760,N32764,N32765);
and and19547(N32761,N32766,in1);
and and19548(N32762,N32767,R1);
and and19549(N32763,N32768,R3);
and and19555(N32775,N32779,N32780);
and and19556(N32776,N32781,N32782);
and and19557(N32777,in2,N32783);
and and19558(N32778,N32784,R2);
and and19564(N32790,N32794,N32795);
and and19565(N32791,N32796,N32797);
and and19566(N32792,N32798,N32799);
and and19567(N32793,R2,R3);
and and19573(N32805,N32809,N32810);
and and19574(N32806,N32811,in1);
and and19575(N32807,N32812,R0);
and and19576(N32808,R1,R3);
and and19582(N32820,N32824,N32825);
and and19583(N32821,N32826,in1);
and and19584(N32822,N32827,N32828);
and and19585(N32823,N32829,R2);
and and19591(N32834,N32838,N32839);
and and19592(N32835,N32840,in1);
and and19593(N32836,N32841,N32842);
and and19594(N32837,R2,R3);
and and19600(N32848,N32852,N32853);
and and19601(N32849,N32854,N32855);
and and19602(N32850,in2,N32856);
and and19603(N32851,R1,R2);
and and19609(N32862,N32866,N32867);
and and19610(N32863,N32868,N32869);
and and19611(N32864,N32870,N32871);
and and19612(N32865,R1,R2);
and and19618(N32876,N32880,N32881);
and and19619(N32877,N32882,in1);
and and19620(N32878,in2,N32883);
and and19621(N32879,R2,R3);
and and19627(N32890,N32894,N32895);
and and19628(N32891,N32896,in1);
and and19629(N32892,R0,N32897);
and and19630(N32893,N32898,R3);
and and19636(N32904,N32908,N32909);
and and19637(N32905,N32910,in1);
and and19638(N32906,in2,N32911);
and and19639(N32907,N32912,R2);
and and19645(N32918,N32922,N32923);
and and19646(N32919,N32924,in1);
and and19647(N32920,N32925,N32926);
and and19648(N32921,N32927,N32928);
and and19654(N32932,N32936,N32937);
and and19655(N32933,N32938,in2);
and and19656(N32934,N32939,R1);
and and19657(N32935,R2,N32940);
and and19663(N32946,N32950,N32951);
and and19664(N32947,N32952,N32953);
and and19665(N32948,in2,N32954);
and and19666(N32949,R1,R2);
and and19672(N32960,N32964,N32965);
and and19673(N32961,N32966,N32967);
and and19674(N32962,R0,R1);
and and19675(N32963,N32968,R3);
and and19681(N32974,N32978,N32979);
and and19682(N32975,N32980,N32981);
and and19683(N32976,in2,R1);
and and19684(N32977,R2,N32982);
and and19690(N32988,N32992,N32993);
and and19691(N32989,N32994,in1);
and and19692(N32990,in2,R0);
and and19693(N32991,R1,N32995);
and and19699(N33002,N33006,N33007);
and and19700(N33003,N33008,N33009);
and and19701(N33004,N33010,N33011);
and and19702(N33005,R2,N33012);
and and19708(N33016,N33020,N33021);
and and19709(N33017,N33022,N33023);
and and19710(N33018,R0,R1);
and and19711(N33019,R2,R3);
and and19717(N33030,N33034,N33035);
and and19718(N33031,N33036,in1);
and and19719(N33032,N33037,R0);
and and19720(N33033,N33038,N33039);
and and19726(N33044,N33048,N33049);
and and19727(N33045,N33050,N33051);
and and19728(N33046,N33052,R1);
and and19729(N33047,R2,N33053);
and and19735(N33058,N33062,N33063);
and and19736(N33059,N33064,in1);
and and19737(N33060,in2,N33065);
and and19738(N33061,N33066,R2);
and and19744(N33072,N33076,N33077);
and and19745(N33073,N33078,N33079);
and and19746(N33074,N33080,R1);
and and19747(N33075,N33081,R3);
and and19753(N33086,N33090,N33091);
and and19754(N33087,N33092,in1);
and and19755(N33088,N33093,R1);
and and19756(N33089,N33094,R3);
and and19762(N33100,N33104,N33105);
and and19763(N33101,N33106,N33107);
and and19764(N33102,R0,R1);
and and19765(N33103,R2,N33108);
and and19771(N33114,N33118,N33119);
and and19772(N33115,N33120,in1);
and and19773(N33116,in2,R0);
and and19774(N33117,N33121,N33122);
and and19780(N33128,N33132,N33133);
and and19781(N33129,N33134,in1);
and and19782(N33130,N33135,R0);
and and19783(N33131,R1,N33136);
and and19789(N33142,N33146,N33147);
and and19790(N33143,N33148,in1);
and and19791(N33144,R0,N33149);
and and19792(N33145,N33150,N33151);
and and19798(N33156,N33160,N33161);
and and19799(N33157,N33162,N33163);
and and19800(N33158,N33164,R0);
and and19801(N33159,N33165,N33166);
and and19807(N33170,N33174,N33175);
and and19808(N33171,N33176,in1);
and and19809(N33172,N33177,R0);
and and19810(N33173,N33178,R2);
and and19816(N33184,N33188,N33189);
and and19817(N33185,N33190,in1);
and and19818(N33186,N33191,N33192);
and and19819(N33187,R1,R2);
and and19825(N33198,N33202,N33203);
and and19826(N33199,N33204,in1);
and and19827(N33200,in2,R0);
and and19828(N33201,N33205,N33206);
and and19834(N33212,N33216,N33217);
and and19835(N33213,N33218,in1);
and and19836(N33214,N33219,R0);
and and19837(N33215,N33220,R3);
and and19843(N33226,N33230,N33231);
and and19844(N33227,N33232,in1);
and and19845(N33228,in2,N33233);
and and19846(N33229,N33234,R3);
and and19852(N33240,N33244,N33245);
and and19853(N33241,N33246,in1);
and and19854(N33242,N33247,N33248);
and and19855(N33243,N33249,R2);
and and19861(N33254,N33258,N33259);
and and19862(N33255,N33260,in1);
and and19863(N33256,in2,R0);
and and19864(N33257,N33261,N33262);
and and19870(N33268,N33272,N33273);
and and19871(N33269,N33274,N33275);
and and19872(N33270,N33276,R0);
and and19873(N33271,N33277,R3);
and and19879(N33282,N33286,N33287);
and and19880(N33283,N33288,N33289);
and and19881(N33284,in2,N33290);
and and19882(N33285,N33291,R2);
and and19888(N33296,N33300,N33301);
and and19889(N33297,N33302,in1);
and and19890(N33298,N33303,N33304);
and and19891(N33299,N33305,R3);
and and19897(N33310,N33314,N33315);
and and19898(N33311,N33316,in1);
and and19899(N33312,N33317,R0);
and and19900(N33313,N33318,N33319);
and and19906(N33324,N33328,N33329);
and and19907(N33325,N33330,in1);
and and19908(N33326,N33331,N33332);
and and19909(N33327,N33333,R2);
and and19915(N33338,N33342,N33343);
and and19916(N33339,N33344,in1);
and and19917(N33340,N33345,N33346);
and and19918(N33341,N33347,R2);
and and19924(N33352,N33356,N33357);
and and19925(N33353,N33358,N33359);
and and19926(N33354,in2,N33360);
and and19927(N33355,N33361,R2);
and and19933(N33366,N33370,N33371);
and and19934(N33367,N33372,in1);
and and19935(N33368,N33373,R0);
and and19936(N33369,N33374,R2);
and and19942(N33380,N33384,N33385);
and and19943(N33381,N33386,in1);
and and19944(N33382,N33387,R0);
and and19945(N33383,R1,N33388);
and and19951(N33394,N33398,N33399);
and and19952(N33395,N33400,in1);
and and19953(N33396,in2,R0);
and and19954(N33397,N33401,N33402);
and and19960(N33408,N33412,N33413);
and and19961(N33409,N33414,N33415);
and and19962(N33410,R0,N33416);
and and19963(N33411,R2,R3);
and and19969(N33421,N33425,N33426);
and and19970(N33422,N33427,N33428);
and and19971(N33423,R0,N33429);
and and19972(N33424,R2,R3);
and and19978(N33434,N33438,N33439);
and and19979(N33435,N33440,N33441);
and and19980(N33436,in2,N33442);
and and19981(N33437,R1,R2);
and and19987(N33447,N33451,N33452);
and and19988(N33448,N33453,N33454);
and and19989(N33449,N33455,R0);
and and19990(N33450,R1,R2);
and and19996(N33460,N33464,N33465);
and and19997(N33461,N33466,in1);
and and19998(N33462,N33467,R0);
and and19999(N33463,R1,R3);
and and20005(N33473,N33477,N33478);
and and20006(N33474,N33479,in2);
and and20007(N33475,R0,N33480);
and and20008(N33476,N33481,R3);
and and20014(N33486,N33490,N33491);
and and20015(N33487,N33492,in1);
and and20016(N33488,in2,N33493);
and and20017(N33489,R1,R2);
and and20023(N33499,N33503,N33504);
and and20024(N33500,N33505,N33506);
and and20025(N33501,in2,R0);
and and20026(N33502,R1,R2);
and and20032(N33512,N33516,N33517);
and and20033(N33513,N33518,N33519);
and and20034(N33514,N33520,R0);
and and20035(N33515,R1,R3);
and and20041(N33525,N33529,N33530);
and and20042(N33526,N33531,in1);
and and20043(N33527,in2,N33532);
and and20044(N33528,R1,R3);
and and20050(N33538,N33542,N33543);
and and20051(N33539,N33544,N33545);
and and20052(N33540,in2,R0);
and and20053(N33541,R1,R2);
and and20059(N33551,N33555,N33556);
and and20060(N33552,N33557,in1);
and and20061(N33553,N33558,R0);
and and20062(N33554,N33559,R2);
and and20068(N33564,N33568,N33569);
and and20069(N33565,in0,N33570);
and and20070(N33566,R0,N33571);
and and20071(N33567,R2,R3);
and and20077(N33577,N33581,N33582);
and and20078(N33578,N33583,N33584);
and and20079(N33579,in2,R0);
and and20080(N33580,N33585,N33586);
and and20086(N33590,N33594,N33595);
and and20087(N33591,N33596,N33597);
and and20088(N33592,in2,N33598);
and and20089(N33593,R1,N33599);
and and20095(N33603,N33607,N33608);
and and20096(N33604,in1,in2);
and and20097(N33605,R0,R1);
and and20098(N33606,R2,N33609);
and and20104(N33616,N33620,N33621);
and and20105(N33617,N33622,in1);
and and20106(N33618,in2,N33623);
and and20107(N33619,R1,R2);
and and20113(N33629,N33633,N33634);
and and20114(N33630,N33635,N33636);
and and20115(N33631,R0,R1);
and and20116(N33632,R2,N33637);
and and20122(N33642,N33646,N33647);
and and20123(N33643,N33648,in2);
and and20124(N33644,R0,N33649);
and and20125(N33645,N33650,R3);
and and20131(N33655,N33659,N33660);
and and20132(N33656,N33661,in1);
and and20133(N33657,in2,N33662);
and and20134(N33658,N33663,R3);
and and20140(N33668,N33672,N33673);
and and20141(N33669,N33674,in1);
and and20142(N33670,N33675,R0);
and and20143(N33671,R2,N33676);
and and20149(N33681,N33685,N33686);
and and20150(N33682,N33687,in1);
and and20151(N33683,in2,R0);
and and20152(N33684,R1,N33688);
and and20158(N33694,N33698,N33699);
and and20159(N33695,N33700,N33701);
and and20160(N33696,in2,N33702);
and and20161(N33697,N33703,R2);
and and20167(N33707,N33711,N33712);
and and20168(N33708,N33713,N33714);
and and20169(N33709,in2,R0);
and and20170(N33710,R1,N33715);
and and20176(N33720,N33724,N33725);
and and20177(N33721,N33726,in1);
and and20178(N33722,in2,N33727);
and and20179(N33723,R1,R2);
and and20185(N33732,N33736,N33737);
and and20186(N33733,N33738,in1);
and and20187(N33734,in2,N33739);
and and20188(N33735,R2,R3);
and and20194(N33744,N33748,N33749);
and and20195(N33745,N33750,in1);
and and20196(N33746,N33751,R1);
and and20197(N33747,R2,R3);
and and20203(N33756,N33760,N33761);
and and20204(N33757,N33762,N33763);
and and20205(N33758,in2,R1);
and and20206(N33759,R2,R3);
and and20212(N33768,N33772,N33773);
and and20213(N33769,N33774,in1);
and and20214(N33770,in2,R0);
and and20215(N33771,R1,R2);
and and20221(N33780,N33784,N33785);
and and20222(N33781,N33786,in1);
and and20223(N33782,R0,R1);
and and20224(N33783,N33787,R3);
and and20230(N33792,N33796,N33797);
and and20231(N33793,N33798,in1);
and and20232(N33794,N33799,R1);
and and20233(N33795,R2,N33800);
and and20239(N33804,N33808,N33809);
and and20240(N33805,N33810,in1);
and and20241(N33806,in2,N33811);
and and20242(N33807,R1,N33812);
and and20248(N33816,N33820,N33821);
and and20249(N33817,N33822,in1);
and and20250(N33818,in2,R0);
and and20251(N33819,R1,R2);
and and20257(N33828,N33832,N33833);
and and20258(N33829,N33834,in1);
and and20259(N33830,in2,R0);
and and20260(N33831,R1,R2);
and and20266(N33840,N33844,N33845);
and and20267(N33841,in1,in2);
and and20268(N33842,R0,N33846);
and and20269(N33843,R2,R3);
and and20275(N33852,N33856,N33857);
and and20276(N33853,in0,in1);
and and20277(N33854,N33858,R0);
and and20278(N33855,N33859,R2);
and and20284(N33864,N33868,N33869);
and and20285(N33865,N33870,in1);
and and20286(N33866,in2,R0);
and and20287(N33867,R1,N33871);
and and20293(N33876,N33880,N33881);
and and20294(N33877,N33882,in1);
and and20295(N33878,in2,N33883);
and and20296(N33879,R2,R3);
and and20302(N33888,N33892,N33893);
and and20303(N33889,N33894,in1);
and and20304(N33890,in2,R0);
and and20305(N33891,R2,R3);
and and20311(N33900,N33904,N33905);
and and20312(N33901,N33906,in1);
and and20313(N33902,in2,R0);
and and20314(N33903,N33907,N33908);
and and20320(N33912,N33916,N33917);
and and20321(N33913,N33918,in1);
and and20322(N33914,N33919,R1);
and and20323(N33915,R2,R3);
and and20329(N33924,N33928,N33929);
and and20330(N33925,N33930,N33931);
and and20331(N33926,in2,R0);
and and20332(N33927,R1,R2);
and and20338(N33936,N33940,N33941);
and and20339(N33937,N33942,in1);
and and20340(N33938,N33943,R1);
and and20341(N33939,R2,R3);
and and20347(N33948,N33952,N33953);
and and20348(N33949,N33954,N33955);
and and20349(N33950,N33956,R0);
and and20350(N33951,R1,R2);
and and20356(N33960,N33964,N33965);
and and20357(N33961,N33966,in1);
and and20358(N33962,N33967,R0);
and and20359(N33963,N33968,R2);
and and20365(N33972,N33976,N33977);
and and20366(N33973,in1,in2);
and and20367(N33974,R0,N33978);
and and20368(N33975,R2,N33979);
and and20374(N33983,N33987,N33988);
and and20375(N33984,in0,in2);
and and20376(N33985,R0,N33989);
and and20377(N33986,R2,R3);
and and20383(N33994,N33998,N33999);
and and20384(N33995,N34000,in1);
and and20385(N33996,in2,R0);
and and20386(N33997,R1,R2);
and and20392(N34005,N34009,N34010);
and and20393(N34006,N34011,in1);
and and20394(N34007,in2,R0);
and and20395(N34008,R1,R2);
and and20401(N34016,N34020,N34021);
and and20402(N34017,in0,in2);
and and20403(N34018,R0,R1);
and and20404(N34019,R2,N34022);
and and20410(N34027,N34031,N34032);
and and20411(N34028,in0,in1);
and and20412(N34029,R0,R1);
and and20413(N34030,R2,N34033);
and and20419(N34038,N34042,N34043);
and and20420(N34039,N34044,in1);
and and20421(N34040,in2,R0);
and and20422(N34041,R1,R2);
and and20428(N34048,N34052,N34053);
and and20429(N34049,N34054,N34055);
and and20430(N34050,N34056,N34057);
and and20431(N34051,R4,N34058);
and and20436(N34064,N34068,N34069);
and and20437(N34065,N34070,N34071);
and and20438(N34066,R0,R1);
and and20439(N34067,N34072,N34073);
and and20444(N34079,N34083,N34084);
and and20445(N34080,N34085,R0);
and and20446(N34081,N34086,N34087);
and and20447(N34082,N34088,N34089);
and and20452(N34094,N34098,N34099);
and and20453(N34095,N34100,N34101);
and and20454(N34096,R0,N34102);
and and20455(N34097,N34103,N34104);
and and20460(N34109,N34113,in0);
and and20461(N34110,N34114,R1);
and and20462(N34111,N34115,N34116);
and and20463(N34112,N34117,N34118);
and and20468(N34123,N34127,N34128);
and and20469(N34124,in1,in2);
and and20470(N34125,N34129,N34130);
and and20471(N34126,R4,N34131);
and and20476(N34137,N34141,N34142);
and and20477(N34138,in1,N34143);
and and20478(N34139,R1,R2);
and and20479(N34140,N34144,N34145);
and and20484(N34151,N34155,N34156);
and and20485(N34152,N34157,N34158);
and and20486(N34153,N34159,R2);
and and20487(N34154,R4,R5);
and and20492(N34165,N34169,N34170);
and and20493(N34166,N34171,in2);
and and20494(N34167,N34172,R2);
and and20495(N34168,R3,N34173);
and and20500(N34179,N34183,N34184);
and and20501(N34180,N34185,N34186);
and and20502(N34181,R2,N34187);
and and20503(N34182,N34188,N34189);
and and20508(N34193,N34197,N34198);
and and20509(N34194,N34199,in2);
and and20510(N34195,N34200,N34201);
and and20511(N34196,R3,R4);
and and20516(N34207,N34211,in0);
and and20517(N34208,N34212,N34213);
and and20518(N34209,N34214,N34215);
and and20519(N34210,R4,R5);
and and20524(N34221,N34225,N34226);
and and20525(N34222,N34227,N34228);
and and20526(N34223,R0,N34229);
and and20527(N34224,R2,N34230);
and and20532(N34235,N34239,in0);
and and20533(N34236,N34240,R1);
and and20534(N34237,N34241,N34242);
and and20535(N34238,N34243,R5);
and and20540(N34249,N34253,N34254);
and and20541(N34250,in1,N34255);
and and20542(N34251,R1,N34256);
and and20543(N34252,N34257,R5);
and and20548(N34263,N34267,N34268);
and and20549(N34264,N34269,N34270);
and and20550(N34265,R1,N34271);
and and20551(N34266,R3,N34272);
and and20556(N34277,N34281,N34282);
and and20557(N34278,in2,N34283);
and and20558(N34279,N34284,R3);
and and20559(N34280,N34285,R5);
and and20564(N34291,N34295,N34296);
and and20565(N34292,N34297,N34298);
and and20566(N34293,N34299,N34300);
and and20567(N34294,R2,R4);
and and20572(N34305,N34309,N34310);
and and20573(N34306,N34311,N34312);
and and20574(N34307,N34313,R2);
and and20575(N34308,N34314,R4);
and and20580(N34319,N34323,in0);
and and20581(N34320,R0,N34324);
and and20582(N34321,N34325,N34326);
and and20583(N34322,R4,N34327);
and and20588(N34332,N34336,N34337);
and and20589(N34333,N34338,R0);
and and20590(N34334,R1,R2);
and and20591(N34335,N34339,R4);
and and20596(N34345,N34349,in0);
and and20597(N34346,N34350,R1);
and and20598(N34347,R2,N34351);
and and20599(N34348,R4,N34352);
and and20604(N34358,N34362,N34363);
and and20605(N34359,in1,N34364);
and and20606(N34360,R1,R2);
and and20607(N34361,N34365,R4);
and and20612(N34371,N34375,N34376);
and and20613(N34372,N34377,N34378);
and and20614(N34373,R1,R2);
and and20615(N34374,R3,N34379);
and and20620(N34384,N34388,N34389);
and and20621(N34385,N34390,N34391);
and and20622(N34386,R0,N34392);
and and20623(N34387,R3,N34393);
and and20628(N34397,N34401,in0);
and and20629(N34398,N34402,R1);
and and20630(N34399,N34403,R3);
and and20631(N34400,N34404,N34405);
and and20636(N34410,N34414,N34415);
and and20637(N34411,N34416,N34417);
and and20638(N34412,R0,R1);
and and20639(N34413,N34418,R5);
and and20644(N34423,N34427,N34428);
and and20645(N34424,N34429,R0);
and and20646(N34425,N34430,R2);
and and20647(N34426,N34431,R4);
and and20652(N34436,N34440,N34441);
and and20653(N34437,in2,R0);
and and20654(N34438,N34442,R2);
and and20655(N34439,R3,R5);
and and20660(N34448,N34452,N34453);
and and20661(N34449,in2,R0);
and and20662(N34450,N34454,R2);
and and20663(N34451,N34455,R5);
and and20668(N34460,N34464,N34465);
and and20669(N34461,in2,R1);
and and20670(N34462,R2,N34466);
and and20671(N34463,R4,R5);
and and20676(N34472,N34476,N34477);
and and20677(N34473,N34478,in2);
and and20678(N34474,R0,N34479);
and and20679(N34475,R2,N34480);
and and20684(N34484,N34488,N34489);
and and20685(N34485,in1,R0);
and and20686(N34486,R1,R2);
and and20687(N34487,N34490,N34491);
and and20692(N34496,N34500,N34501);
and and20693(N34497,in1,N34502);
and and20694(N34498,R1,R2);
and and20695(N34499,R3,R4);
and and20700(N34508,N34512,N34513);
and and20701(N34509,in1,in2);
and and20702(N34510,R2,N34514);
and and20703(N34511,N34515,R5);
and and20708(N34520,N34524,N34525);
and and20709(N34521,in1,N34526);
and and20710(N34522,N34527,R1);
and and20711(N34523,R2,R3);
and and20716(N34532,N34536,N34537);
and and20717(N34533,in2,R0);
and and20718(N34534,N34538,R2);
and and20719(N34535,N34539,R4);
and and20724(N34544,N34548,N34549);
and and20725(N34545,N34550,R0);
and and20726(N34546,N34551,R2);
and and20727(N34547,R3,R4);
and and20732(N34556,N34560,N34561);
and and20733(N34557,N34562,in2);
and and20734(N34558,R0,R1);
and and20735(N34559,N34563,R4);
and and20740(N34568,N34572,in0);
and and20741(N34569,R0,R1);
and and20742(N34570,R2,N34573);
and and20743(N34571,N34574,R5);
and and20748(N34580,N34584,in0);
and and20749(N34581,N34585,N34586);
and and20750(N34582,R2,N34587);
and and20751(N34583,R4,R5);
and and20756(N34592,N34596,in0);
and and20757(N34593,N34597,N34598);
and and20758(N34594,R2,N34599);
and and20759(N34595,R4,N34600);
and and20764(N34604,N34608,in0);
and and20765(N34605,R0,R1);
and and20766(N34606,N34609,N34610);
and and20767(N34607,R4,R5);
and and20772(N34616,N34620,N34621);
and and20773(N34617,in1,in2);
and and20774(N34618,R0,R2);
and and20775(N34619,N34622,N34623);
and and20780(N34628,N34632,N34633);
and and20781(N34629,in1,in2);
and and20782(N34630,R0,N34634);
and and20783(N34631,R3,N34635);
and and20788(N34640,N34644,N34645);
and and20789(N34641,in1,in2);
and and20790(N34642,N34646,R1);
and and20791(N34643,R3,N34647);
and and20796(N34652,N34656,N34657);
and and20797(N34653,in1,N34658);
and and20798(N34654,R0,R1);
and and20799(N34655,R2,N34659);
and and20804(N34664,N34668,N34669);
and and20805(N34665,N34670,R0);
and and20806(N34666,R1,N34671);
and and20807(N34667,R3,N34672);
and and20812(N34676,N34680,N34681);
and and20813(N34677,N34682,in2);
and and20814(N34678,R0,R1);
and and20815(N34679,R4,N34683);
and and20820(N34688,N34692,N34693);
and and20821(N34689,N34694,N34695);
and and20822(N34690,R0,R1);
and and20823(N34691,R3,N34696);
and and20828(N34700,N34704,N34705);
and and20829(N34701,in2,N34706);
and and20830(N34702,N34707,R3);
and and20831(N34703,R4,R5);
and and20836(N34711,N34715,in0);
and and20837(N34712,N34716,R1);
and and20838(N34713,N34717,R3);
and and20839(N34714,R4,R5);
and and20844(N34722,N34726,N34727);
and and20845(N34723,N34728,in2);
and and20846(N34724,R1,R2);
and and20847(N34725,N34729,R4);
and and20852(N34733,N34737,N34738);
and and20853(N34734,in1,N34739);
and and20854(N34735,N34740,R1);
and and20855(N34736,R2,R3);
and and20860(N34744,N34748,N34749);
and and20861(N34745,N34750,in2);
and and20862(N34746,R0,R2);
and and20863(N34747,R3,N34751);
and and20868(N34755,N34759,in0);
and and20869(N34756,R0,N34760);
and and20870(N34757,R2,N34761);
and and20871(N34758,R4,R5);
and and20876(N34765,N34769,in0);
and and20877(N34766,R0,R1);
and and20878(N34767,R2,N34770);
and and20879(N34768,R4,N34771);
and and20884(N34775,N34779,in0);
and and20885(N34776,R0,R1);
and and20886(N34777,R2,N34780);
and and20887(N34778,R4,R5);
and and20892(N34785,N34789,in0);
and and20893(N34786,R0,R1);
and and20894(N34787,N34790,R3);
and and20895(N34788,R4,R5);
and and20900(N34794,in0,R0);
and and20901(N34795,N34798,N34799);
and and20902(N34796,R3,N34800);
and and20903(N34797,N34801,R7);
and and20907(N34805,in0,R0);
and and20908(N34806,N34809,N34810);
and and20909(N34807,N34811,N34812);
and and20910(N34808,R6,R7);
and and20914(N34816,in0,N34820);
and and20915(N34817,N34821,N34822);
and and20916(N34818,R3,R4);
and and20917(N34819,R6,N34823);
and and19000(N31791,N31796,R3);
and and19001(N31792,R4,R5);
and and19002(N31793,N31797,N31798);
and and19010(N31806,N31813,N31814);
and and19011(N31807,N31815,N31816);
and and19019(N31824,N31832,N31833);
and and19020(N31825,R6,N31834);
and and19028(N31842,N31849,N31850);
and and19029(N31843,N31851,N31852);
and and19037(N31860,N31867,N31868);
and and19038(N31861,N31869,N31870);
and and19046(N31878,N31886,R5);
and and19047(N31879,N31887,N31888);
and and19055(N31896,N31903,N31904);
and and19056(N31897,N31905,N31906);
and and19064(N31914,N31922,N31923);
and and19065(N31915,N31924,R7);
and and19073(N31932,N31938,N31939);
and and19074(N31933,N31940,N31941);
and and19082(N31949,N31956,N31957);
and and19083(N31950,N31958,R7);
and and19091(N31966,N31974,R5);
and and19092(N31967,N31975,R7);
and and19100(N31983,N31990,N31991);
and and19101(N31984,R6,N31992);
and and19109(N32000,R3,N32008);
and and19110(N32001,N32009,R7);
and and19118(N32017,R3,R5);
and and19119(N32018,N32025,N32026);
and and19127(N32034,N32039,N32040);
and and19128(N32035,N32041,N32042);
and and19136(N32050,N32056,N32057);
and and19137(N32051,R6,N32058);
and and19145(N32066,N32072,N32073);
and and19146(N32067,R6,N32074);
and and19154(N32082,N32088,N32089);
and and19155(N32083,N32090,R7);
and and19163(N32098,N32104,N32105);
and and19164(N32099,R5,N32106);
and and19172(N32114,N32120,R5);
and and19173(N32115,N32121,N32122);
and and19181(N32130,N32136,N32137);
and and19182(N32131,R6,N32138);
and and19190(N32146,N32152,R5);
and and19191(N32147,N32153,N32154);
and and19199(N32162,N32169,R5);
and and19200(N32163,R6,N32170);
and and19208(N32178,N32184,N32185);
and and19209(N32179,N32186,R7);
and and19217(N32194,R3,N32200);
and and19218(N32195,N32201,N32202);
and and19226(N32210,N32216,N32217);
and and19227(N32211,N32218,R7);
and and19235(N32226,N32231,N32232);
and and19236(N32227,N32233,N32234);
and and19244(N32242,N32248,N32249);
and and19245(N32243,R5,N32250);
and and19253(N32258,N32264,N32265);
and and19254(N32259,R5,N32266);
and and19262(N32274,N32280,N32281);
and and19263(N32275,N32282,R7);
and and19271(N32290,N32297,R5);
and and19272(N32291,N32298,R7);
and and19280(N32306,N32313,R5);
and and19281(N32307,N32314,R7);
and and19289(N32322,N32328,N32329);
and and19290(N32323,R6,N32330);
and and19298(N32338,R3,R4);
and and19299(N32339,N32345,N32346);
and and19307(N32354,N32360,N32361);
and and19308(N32355,R6,N32362);
and and19316(N32370,N32376,N32377);
and and19317(N32371,R6,N32378);
and and19325(N32386,N32392,N32393);
and and19326(N32387,R6,N32394);
and and19334(N32402,R3,N32408);
and and19335(N32403,N32409,N32410);
and and19343(N32418,R3,N32425);
and and19344(N32419,R5,N32426);
and and19352(N32434,R4,R5);
and and19353(N32435,N32441,R7);
and and19361(N32449,N32453,N32454);
and and19362(N32450,N32455,N32456);
and and19370(N32464,N32468,N32469);
and and19371(N32465,N32470,N32471);
and and19379(N32479,N32483,N32484);
and and19380(N32480,N32485,N32486);
and and19388(N32494,R4,N32499);
and and19389(N32495,N32500,N32501);
and and19397(N32509,R3,N32514);
and and19398(N32510,N32515,N32516);
and and19406(N32524,R4,N32530);
and and19407(N32525,N32531,R7);
and and19415(N32539,R4,R5);
and and19416(N32540,N32545,N32546);
and and19424(N32554,N32559,N32560);
and and19425(N32555,N32561,R7);
and and19433(N32569,R4,N32574);
and and19434(N32570,N32575,N32576);
and and19442(N32584,N32590,R4);
and and19443(N32585,R5,N32591);
and and19451(N32599,N32604,R5);
and and19452(N32600,N32605,N32606);
and and19460(N32614,R3,N32620);
and and19461(N32615,N32621,R7);
and and19469(N32629,R4,N32635);
and and19470(N32630,R6,N32636);
and and19478(N32644,R4,N32650);
and and19479(N32645,R6,N32651);
and and19487(N32659,R3,R4);
and and19488(N32660,R5,R7);
and and19496(N32674,N32679,N32680);
and and19497(N32675,N32681,R6);
and and19505(N32689,R3,N32695);
and and19506(N32690,R6,N32696);
and and19514(N32704,R3,N32709);
and and19515(N32705,N32710,N32711);
and and19523(N32719,N32723,N32724);
and and19524(N32720,N32725,N32726);
and and19532(N32734,R3,N32741);
and and19533(N32735,R6,R7);
and and19541(N32749,R4,N32755);
and and19542(N32750,N32756,R7);
and and19550(N32764,N32769,N32770);
and and19551(N32765,N32771,R7);
and and19559(N32779,R4,N32785);
and and19560(N32780,N32786,R7);
and and19568(N32794,N32800,R5);
and and19569(N32795,R6,N32801);
and and19577(N32809,N32813,N32814);
and and19578(N32810,N32815,N32816);
and and19586(N32824,R3,R4);
and and19587(N32825,R5,N32830);
and and19595(N32838,N32843,R5);
and and19596(N32839,N32844,R7);
and and19604(N32852,N32857,N32858);
and and19605(N32853,R6,R7);
and and19613(N32866,R3,R5);
and and19614(N32867,N32872,R7);
and and19622(N32880,N32884,N32885);
and and19623(N32881,R6,N32886);
and and19631(N32894,R4,R5);
and and19632(N32895,N32899,N32900);
and and19640(N32908,R3,N32913);
and and19641(N32909,N32914,R7);
and and19649(N32922,R3,R5);
and and19650(N32923,R6,R7);
and and19658(N32936,N32941,R5);
and and19659(N32937,N32942,R7);
and and19667(N32950,R3,N32955);
and and19668(N32951,R6,N32956);
and and19676(N32964,R4,N32969);
and and19677(N32965,R6,N32970);
and and19685(N32978,N32983,R5);
and and19686(N32979,R6,N32984);
and and19694(N32992,N32996,N32997);
and and19695(N32993,N32998,R7);
and and19703(N33006,R4,R5);
and and19704(N33007,R6,R7);
and and19712(N33020,N33024,N33025);
and and19713(N33021,N33026,R7);
and and19721(N33034,R3,R4);
and and19722(N33035,N33040,R7);
and and19730(N33048,R4,N33054);
and and19731(N33049,R6,R7);
and and19739(N33062,N33067,N33068);
and and19740(N33063,R6,R7);
and and19748(N33076,N33082,R5);
and and19749(N33077,R6,R7);
and and19757(N33090,N33095,R5);
and and19758(N33091,R6,N33096);
and and19766(N33104,N33109,N33110);
and and19767(N33105,R6,R7);
and and19775(N33118,N33123,N33124);
and and19776(N33119,R5,R6);
and and19784(N33132,N33137,R4);
and and19785(N33133,N33138,R7);
and and19793(N33146,R4,R5);
and and19794(N33147,R6,N33152);
and and19802(N33160,R4,R5);
and and19803(N33161,R6,R7);
and and19811(N33174,R3,N33179);
and and19812(N33175,R6,N33180);
and and19820(N33188,R3,R5);
and and19821(N33189,N33193,N33194);
and and19829(N33202,N33207,N33208);
and and19830(N33203,R6,R7);
and and19838(N33216,N33221,N33222);
and and19839(N33217,R6,R7);
and and19847(N33230,R4,N33235);
and and19848(N33231,R6,N33236);
and and19856(N33244,R3,R4);
and and19857(N33245,N33250,R7);
and and19865(N33258,R4,R5);
and and19866(N33259,N33263,N33264);
and and19874(N33272,R4,R5);
and and19875(N33273,N33278,R7);
and and19883(N33286,N33292,R5);
and and19884(N33287,R6,R7);
and and19892(N33300,R4,R5);
and and19893(N33301,N33306,R7);
and and19901(N33314,R3,R5);
and and19902(N33315,N33320,R7);
and and19910(N33328,R3,N33334);
and and19911(N33329,R6,R7);
and and19919(N33342,R3,R5);
and and19920(N33343,R6,N33348);
and and19928(N33356,R3,N33362);
and and19929(N33357,R5,R6);
and and19937(N33370,N33375,N33376);
and and19938(N33371,R6,R7);
and and19946(N33384,R3,R4);
and and19947(N33385,N33389,N33390);
and and19955(N33398,R4,N33403);
and and19956(N33399,N33404,R7);
and and19964(N33412,R4,R5);
and and19965(N33413,R6,N33417);
and and19973(N33425,R4,N33430);
and and19974(N33426,R6,R7);
and and19982(N33438,R3,R4);
and and19983(N33439,N33443,R7);
and and19991(N33451,N33456,R4);
and and19992(N33452,R5,R6);
and and20000(N33464,R4,N33468);
and and20001(N33465,R6,N33469);
and and20009(N33477,N33482,R5);
and and20010(N33478,R6,R7);
and and20018(N33490,N33494,R4);
and and20019(N33491,N33495,R7);
and and20027(N33503,R4,N33507);
and and20028(N33504,R6,N33508);
and and20036(N33516,R4,R5);
and and20037(N33517,R6,N33521);
and and20045(N33529,N33533,R5);
and and20046(N33530,R6,N33534);
and and20054(N33542,R3,R4);
and and20055(N33543,N33546,N33547);
and and20063(N33555,R4,R5);
and and20064(N33556,N33560,R7);
and and20072(N33568,R4,N33572);
and and20073(N33569,R6,N33573);
and and20081(N33581,R4,R5);
and and20082(N33582,R6,R7);
and and20090(N33594,R3,R4);
and and20091(N33595,R5,R7);
and and20099(N33607,N33610,R5);
and and20100(N33608,N33611,N33612);
and and20108(N33620,R3,N33624);
and and20109(N33621,R5,N33625);
and and20117(N33633,N33638,R5);
and and20118(N33634,R6,R7);
and and20126(N33646,R4,R5);
and and20127(N33647,N33651,R7);
and and20135(N33659,R4,R5);
and and20136(N33660,N33664,R7);
and and20144(N33672,R4,R5);
and and20145(N33673,R6,N33677);
and and20153(N33685,R3,N33689);
and and20154(N33686,R5,N33690);
and and20162(N33698,R4,R5);
and and20163(N33699,R6,R7);
and and20171(N33711,R3,R4);
and and20172(N33712,R6,N33716);
and and20180(N33724,R3,N33728);
and and20181(N33725,R6,R7);
and and20189(N33736,R4,N33740);
and and20190(N33737,R6,R7);
and and20198(N33748,R4,R5);
and and20199(N33749,N33752,R7);
and and20207(N33760,N33764,R5);
and and20208(N33761,R6,R7);
and and20216(N33772,R3,N33775);
and and20217(N33773,N33776,R7);
and and20225(N33784,N33788,R5);
and and20226(N33785,R6,R7);
and and20234(N33796,R4,R5);
and and20235(N33797,R6,R7);
and and20243(N33808,R3,R5);
and and20244(N33809,R6,R7);
and and20252(N33820,R3,N33823);
and and20253(N33821,R6,N33824);
and and20261(N33832,N33835,N33836);
and and20262(N33833,R6,R7);
and and20270(N33844,R4,N33847);
and and20271(N33845,R6,N33848);
and and20279(N33856,R3,R4);
and and20280(N33857,R6,N33860);
and and20288(N33868,R3,N33872);
and and20289(N33869,R6,R7);
and and20297(N33880,N33884,R5);
and and20298(N33881,R6,R7);
and and20306(N33892,R4,R5);
and and20307(N33893,N33895,N33896);
and and20315(N33904,R3,R5);
and and20316(N33905,R6,R7);
and and20324(N33916,R4,R5);
and and20325(N33917,R6,N33920);
and and20333(N33928,R3,R4);
and and20334(N33929,R5,N33932);
and and20342(N33940,R4,N33944);
and and20343(N33941,R6,R7);
and and20351(N33952,R4,R5);
and and20352(N33953,R6,R7);
and and20360(N33964,R3,R4);
and and20361(N33965,R5,R7);
and and20369(N33976,R4,R5);
and and20370(N33977,R6,R7);
and and20378(N33987,R4,R5);
and and20379(N33988,R6,N33990);
and and20387(N33998,N34001,R4);
and and20388(N33999,R5,R6);
and and20396(N34009,R3,N34012);
and and20397(N34010,R5,R6);
and and20405(N34020,N34023,R5);
and and20406(N34021,R6,R7);
and and20414(N34031,N34034,R5);
and and20415(N34032,R6,R7);
and and20423(N34042,R3,R5);
and and20424(N34043,R6,R7);
and and20432(N34052,N34059,N34060);
and and20440(N34068,N34074,N34075);
and and20448(N34083,R5,N34090);
and and20456(N34098,R5,N34105);
and and20464(N34113,N34119,R7);
and and20472(N34127,N34132,N34133);
and and20480(N34141,N34146,N34147);
and and20488(N34155,N34160,N34161);
and and20496(N34169,N34174,N34175);
and and20504(N34183,R6,R7);
and and20512(N34197,N34202,N34203);
and and20520(N34211,N34216,N34217);
and and20528(N34225,R4,N34231);
and and20536(N34239,N34244,N34245);
and and20544(N34253,N34258,N34259);
and and20552(N34267,N34273,R7);
and and20560(N34281,N34286,N34287);
and and20568(N34295,N34301,R7);
and and20576(N34309,N34315,R7);
and and20584(N34323,R6,N34328);
and and20592(N34336,N34340,N34341);
and and20600(N34349,N34353,N34354);
and and20608(N34362,N34366,N34367);
and and20616(N34375,R5,N34380);
and and20624(N34388,R6,R7);
and and20632(N34401,R6,N34406);
and and20640(N34414,N34419,R7);
and and20648(N34427,N34432,R7);
and and20656(N34440,N34443,N34444);
and and20664(N34452,N34456,R7);
and and20672(N34464,N34467,N34468);
and and20680(N34476,R6,R7);
and and20688(N34488,N34492,R7);
and and20696(N34500,N34503,N34504);
and and20704(N34512,R6,N34516);
and and20712(N34524,R6,N34528);
and and20720(N34536,R5,N34540);
and and20728(N34548,N34552,R7);
and and20736(N34560,N34564,R7);
and and20744(N34572,N34575,N34576);
and and20752(N34584,R6,N34588);
and and20760(N34596,R6,R7);
and and20768(N34608,N34611,N34612);
and and20776(N34620,R6,N34624);
and and20784(N34632,R6,N34636);
and and20792(N34644,N34648,R7);
and and20800(N34656,R4,N34660);
and and20808(N34668,R6,R7);
and and20816(N34680,N34684,R7);
and and20824(N34692,R6,R7);
and and20832(N34704,R6,R7);
and and20840(N34715,N34718,R7);
and and20848(N34726,R5,R7);
and and20856(N34737,R4,R6);
and and20864(N34748,R6,R7);
and and20872(N34759,R6,R7);
and and20880(N34769,R6,R7);
and and20888(N34779,N34781,R7);
and and20896(N34789,R6,R7);
and and20918(N34877,N34878,N34879);
and and20925(N34889,N34890,N34891);
and and20931(N34901,N34902,N34903);
and and20937(N34913,N34914,N34915);
and and20943(N34925,N34926,N34927);
and and20949(N34937,N34938,N34939);
and and20955(N34948,N34949,N34950);
and and20961(N34959,N34960,N34961);
and and20967(N34970,N34971,N34972);
and and20973(N34981,N34982,N34983);
and and20979(N34992,N34993,N34994);
and and20985(N35002,N35003,N35004);
and and20991(N35012,N35013,N35014);
and and20997(N35022,N35023,N35024);
and and21003(N35032,N35033,N35034);
and and21009(N35042,N35043,N35044);
and and21015(N35052,N35053,N35054);
and and21021(N35062,N35063,N35064);
and and21027(N35072,N35073,N35074);
and and21033(N35082,N35083,N35084);
and and21039(N35092,N35093,N35094);
and and21045(N35102,N35103,N35104);
and and21051(N35112,N35113,N35114);
and and21057(N35122,N35123,N35124);
and and21063(N35131,N35132,N35133);
and and21069(N35140,N35141,N35142);
and and21075(N35149,N35150,N35151);
and and21081(N35158,N35159,N35160);
and and21087(N35167,N35168,N35169);
and and21093(N35176,N35177,N35178);
and and21099(N35185,N35186,N35187);
and and21105(N35194,N35195,N35196);
and and21111(N35203,N35204,N35205);
and and21117(N35212,N35213,N35214);
and and21123(N35221,N35222,N35223);
and and21129(N35230,N35231,N35232);
and and21135(N35238,N35239,N35240);
and and21141(N35246,N35247,N35248);
and and21147(N35254,N35255,N35256);
and and21153(N35262,N35263,N35264);
and and21159(N35270,N35271,N35272);
and and21165(N35278,N35279,N35280);
and and21171(N35285,N35286,N35287);
and and21177(N35292,N35293,N35294);
and and21183(N35299,N35300,N35301);
and and21189(N35306,N35307,N35308);
and and21195(N35313,N35314,N35315);
and and21201(N35320,N35321,N35322);
and and21207(N35327,N35328,N35329);
and and21212(N35337,N35338,N35339);
and and21217(N35345,N35346,N35347);
and and21222(N35353,N35354,N35355);
and and21227(N35361,N35362,N35363);
and and21232(N35369,N35370,N35371);
and and20919(N34878,N34880,N34881);
and and20920(N34879,N34882,N34883);
and and20926(N34890,N34892,N34893);
and and20927(N34891,N34894,N34895);
and and20932(N34902,N34904,N34905);
and and20933(N34903,N34906,R0);
and and20938(N34914,N34916,N34917);
and and20939(N34915,N34918,N34919);
and and20944(N34926,N34928,N34929);
and and20945(N34927,N34930,N34931);
and and20950(N34938,N34940,N34941);
and and20951(N34939,N34942,N34943);
and and20956(N34949,N34951,N34952);
and and20957(N34950,N34953,N34954);
and and20962(N34960,N34962,N34963);
and and20963(N34961,N34964,N34965);
and and20968(N34971,N34973,N34974);
and and20969(N34972,N34975,N34976);
and and20974(N34982,N34984,N34985);
and and20975(N34983,N34986,N34987);
and and20980(N34993,N34995,N34996);
and and20981(N34994,N34997,N34998);
and and20986(N35003,N35005,N35006);
and and20987(N35004,N35007,N35008);
and and20992(N35013,N35015,N35016);
and and20993(N35014,N35017,N35018);
and and20998(N35023,N35025,N35026);
and and20999(N35024,N35027,R0);
and and21004(N35033,N35035,N35036);
and and21005(N35034,N35037,N35038);
and and21010(N35043,N35045,N35046);
and and21011(N35044,N35047,R0);
and and21016(N35053,N35055,N35056);
and and21017(N35054,N35057,N35058);
and and21022(N35063,N35065,N35066);
and and21023(N35064,N35067,R0);
and and21028(N35073,N35075,N35076);
and and21029(N35074,N35077,R0);
and and21034(N35083,N35085,N35086);
and and21035(N35084,N35087,N35088);
and and21040(N35093,N35095,N35096);
and and21041(N35094,N35097,R0);
and and21046(N35103,N35105,N35106);
and and21047(N35104,N35107,R0);
and and21052(N35113,N35115,N35116);
and and21053(N35114,N35117,R0);
and and21058(N35123,N35125,N35126);
and and21059(N35124,N35127,R0);
and and21064(N35132,N35134,N35135);
and and21065(N35133,N35136,N35137);
and and21070(N35141,N35143,N35144);
and and21071(N35142,N35145,N35146);
and and21076(N35150,N35152,N35153);
and and21077(N35151,N35154,N35155);
and and21082(N35159,N35161,N35162);
and and21083(N35160,N35163,N35164);
and and21088(N35168,N35170,N35171);
and and21089(N35169,N35172,R0);
and and21094(N35177,N35179,N35180);
and and21095(N35178,N35181,N35182);
and and21100(N35186,N35188,N35189);
and and21101(N35187,N35190,N35191);
and and21106(N35195,N35197,N35198);
and and21107(N35196,N35199,R0);
and and21112(N35204,N35206,N35207);
and and21113(N35205,N35208,N35209);
and and21118(N35213,N35215,N35216);
and and21119(N35214,N35217,R0);
and and21124(N35222,N35224,N35225);
and and21125(N35223,N35226,R0);
and and21130(N35231,N35233,N35234);
and and21131(N35232,N35235,R0);
and and21136(N35239,N35241,N35242);
and and21137(N35240,N35243,R0);
and and21142(N35247,N35249,N35250);
and and21143(N35248,N35251,N35252);
and and21148(N35255,N35257,N35258);
and and21149(N35256,N35259,R0);
and and21154(N35263,N35265,N35266);
and and21155(N35264,N35267,N35268);
and and21160(N35271,N35273,N35274);
and and21161(N35272,N35275,R0);
and and21166(N35279,N35281,N35282);
and and21167(N35280,N35283,R0);
and and21172(N35286,N35288,N35289);
and and21173(N35287,N35290,N35291);
and and21178(N35293,N35295,N35296);
and and21179(N35294,N35297,R0);
and and21184(N35300,N35302,N35303);
and and21185(N35301,N35304,R1);
and and21190(N35307,N35309,N35310);
and and21191(N35308,N35311,R0);
and and21196(N35314,N35316,N35317);
and and21197(N35315,N35318,N35319);
and and21202(N35321,N35323,N35324);
and and21203(N35322,N35325,N35326);
and and21208(N35328,N35330,N35331);
and and21209(N35329,N35332,N35333);
and and21213(N35338,N35340,N35341);
and and21214(N35339,R0,N35342);
and and21218(N35346,N35348,N35349);
and and21219(N35347,R0,N35350);
and and21223(N35354,N35356,N35357);
and and21224(N35355,N35358,R1);
and and21228(N35362,N35364,N35365);
and and21229(N35363,R1,R2);
and and21233(N35370,N35372,N35373);
and and21234(N35371,R0,R1);
and and20921(N34880,R0,N34884);
and and20922(N34881,N34885,R3);
and and20923(N34882,N34886,R5);
and and20924(N34883,N34887,N34888);
and and20928(N34892,R1,N34896);
and and20929(N34893,N34897,N34898);
and and20930(N34894,N34899,N34900);
and and20934(N34904,N34907,N34908);
and and20935(N34905,N34909,N34910);
and and20936(N34906,N34911,N34912);
and and20940(N34916,N34920,N34921);
and and20941(N34917,N34922,N34923);
and and20942(N34918,R6,N34924);
and and20946(N34928,N34932,N34933);
and and20947(N34929,N34934,N34935);
and and20948(N34930,N34936,R7);
and and20952(N34940,R2,R3);
and and20953(N34941,N34944,N34945);
and and20954(N34942,N34946,N34947);
and and20958(N34951,N34955,R2);
and and20959(N34952,N34956,N34957);
and and20960(N34953,R5,N34958);
and and20964(N34962,N34966,N34967);
and and20965(N34963,N34968,R5);
and and20966(N34964,N34969,R7);
and and20970(N34973,R1,N34977);
and and20971(N34974,N34978,N34979);
and and20972(N34975,R5,N34980);
and and20976(N34984,R1,N34988);
and and20977(N34985,R3,N34989);
and and20978(N34986,N34990,N34991);
and and20982(N34995,R1,R2);
and and20983(N34996,N34999,N35000);
and and20984(N34997,N35001,R7);
and and20988(N35005,N35009,R2);
and and20989(N35006,R3,N35010);
and and20990(N35007,N35011,R7);
and and20994(N35015,N35019,R3);
and and20995(N35016,R4,N35020);
and and20996(N35017,N35021,R7);
and and21000(N35025,N35028,N35029);
and and21001(N35026,N35030,R4);
and and21002(N35027,N35031,R7);
and and21006(N35035,R1,N35039);
and and21007(N35036,R3,R4);
and and21008(N35037,N35040,N35041);
and and21012(N35045,N35048,N35049);
and and21013(N35046,R3,N35050);
and and21014(N35047,N35051,R7);
and and21018(N35055,N35059,R2);
and and21019(N35056,R3,R4);
and and21020(N35057,N35060,N35061);
and and21024(N35065,N35068,N35069);
and and21025(N35066,R3,R4);
and and21026(N35067,N35070,N35071);
and and21030(N35075,N35078,N35079);
and and21031(N35076,N35080,N35081);
and and21032(N35077,R6,R7);
and and21036(N35085,N35089,N35090);
and and21037(N35086,R3,R4);
and and21038(N35087,R6,N35091);
and and21042(N35095,N35098,N35099);
and and21043(N35096,R4,R5);
and and21044(N35097,N35100,N35101);
and and21048(N35105,R1,N35108);
and and21049(N35106,N35109,R5);
and and21050(N35107,N35110,N35111);
and and21054(N35115,N35118,N35119);
and and21055(N35116,R4,N35120);
and and21056(N35117,N35121,R7);
and and21060(N35125,N35128,R2);
and and21061(N35126,N35129,R5);
and and21062(N35127,N35130,R7);
and and21066(N35134,N35138,R2);
and and21067(N35135,R4,R5);
and and21068(N35136,N35139,R7);
and and21072(N35143,R1,N35147);
and and21073(N35144,R3,R5);
and and21074(N35145,N35148,R7);
and and21078(N35152,N35156,N35157);
and and21079(N35153,R3,R5);
and and21080(N35154,R6,R7);
and and21084(N35161,R1,R2);
and and21085(N35162,N35165,R5);
and and21086(N35163,N35166,R7);
and and21090(N35170,N35173,R2);
and and21091(N35171,R3,N35174);
and and21092(N35172,N35175,R6);
and and21096(N35179,N35183,R2);
and and21097(N35180,N35184,R4);
and and21098(N35181,R5,R6);
and and21102(N35188,R1,R2);
and and21103(N35189,R3,N35192);
and and21104(N35190,R5,N35193);
and and21108(N35197,R1,R2);
and and21109(N35198,R3,N35200);
and and21110(N35199,N35201,N35202);
and and21114(N35206,N35210,R2);
and and21115(N35207,N35211,R4);
and and21116(N35208,R6,R7);
and and21120(N35215,R1,N35218);
and and21121(N35216,R4,R5);
and and21122(N35217,N35219,N35220);
and and21126(N35224,R1,R2);
and and21127(N35225,R3,N35227);
and and21128(N35226,N35228,N35229);
and and21132(N35233,R1,R2);
and and21133(N35234,N35236,N35237);
and and21134(N35235,R5,R6);
and and21138(N35241,N35244,R2);
and and21139(N35242,R3,R4);
and and21140(N35243,N35245,R7);
and and21144(N35249,R1,R2);
and and21145(N35250,R3,R4);
and and21146(N35251,R6,N35253);
and and21150(N35257,R1,R2);
and and21151(N35258,N35260,N35261);
and and21152(N35259,R6,R7);
and and21156(N35265,R2,N35269);
and and21157(N35266,R4,R5);
and and21158(N35267,R6,R7);
and and21162(N35273,R1,R2);
and and21163(N35274,N35276,R4);
and and21164(N35275,R5,N35277);
and and21168(N35281,R1,R2);
and and21169(N35282,R3,R4);
and and21170(N35283,R5,N35284);
and and21174(N35288,R1,R3);
and and21175(N35289,R4,R5);
and and21176(N35290,R6,R7);
and and21180(N35295,R2,R3);
and and21181(N35296,R4,R5);
and and21182(N35297,R6,N35298);
and and21186(N35302,R2,R3);
and and21187(N35303,R4,N35305);
and and21188(N35304,R6,R7);
and and21192(N35309,N35312,R3);
and and21193(N35310,R4,R5);
and and21194(N35311,R6,R7);
and and21198(N35316,R2,R3);
and and21199(N35317,R4,R5);
and and21200(N35318,R6,R7);
and and21204(N35323,R1,R2);
and and21205(N35324,R3,R4);
and and21206(N35325,R5,R7);
and and21210(N35330,N35334,R4);
and and21211(N35331,N35335,N35336);
and and21215(N35340,N35343,N35344);
and and21216(N35341,R5,R6);
and and21220(N35348,R4,N35351);
and and21221(N35349,R6,N35352);
and and21225(N35356,R2,N35359);
and and21226(N35357,R4,N35360);
and and21230(N35364,N35366,R4);
and and21231(N35365,N35367,N35368);
and and21235(N35372,N35374,R3);
and and21236(N35373,R6,R7);
and and21237(N35411,N35412,N35413);
and and21244(N35423,N35424,N35425);
and and21251(N35435,N35436,N35437);
and and21258(N35446,N35447,N35448);
and and21265(N35456,N35457,N35458);
and and21272(N35465,N35466,N35467);
and and21278(N35477,N35478,N35479);
and and21284(N35489,N35490,N35491);
and and21290(N35500,N35501,N35502);
and and21296(N35510,N35511,N35512);
and and21302(N35520,N35521,N35522);
and and21308(N35530,N35531,N35532);
and and21314(N35540,N35541,N35542);
and and21320(N35550,N35551,N35552);
and and21326(N35560,N35561,N35562);
and and21332(N35570,N35571,N35572);
and and21338(N35580,N35581,N35582);
and and21344(N35590,N35591,N35592);
and and21350(N35600,N35601,N35602);
and and21356(N35609,N35610,N35611);
and and21362(N35618,N35619,N35620);
and and21368(N35627,N35628,N35629);
and and21374(N35636,N35637,N35638);
and and21380(N35645,N35646,N35647);
and and21386(N35654,N35655,N35656);
and and21392(N35663,N35664,N35665);
and and21398(N35672,N35673,N35674);
and and21404(N35681,N35682,N35683);
and and21410(N35690,N35691,N35692);
and and21416(N35698,N35699,N35700);
and and21422(N35706,N35707,N35708);
and and21428(N35714,N35715,N35716);
and and21434(N35722,N35723,N35724);
and and21440(N35730,N35731,N35732);
and and21446(N35738,N35739,N35740);
and and21452(N35745,N35746,N35747);
and and21458(N35752,N35753,N35754);
and and21238(N35412,N35414,N35415);
and and21239(N35413,N35416,N35417);
and and21245(N35424,N35426,N35427);
and and21246(N35425,N35428,N35429);
and and21252(N35436,N35438,N35439);
and and21253(N35437,N35440,N35441);
and and21259(N35447,N35449,N35450);
and and21260(N35448,N35451,N35452);
and and21266(N35457,N35459,N35460);
and and21267(N35458,N35461,N35462);
and and21273(N35466,N35468,N35469);
and and21274(N35467,N35470,N35471);
and and21279(N35478,N35480,N35481);
and and21280(N35479,N35482,N35483);
and and21285(N35490,N35492,N35493);
and and21286(N35491,N35494,N35495);
and and21291(N35501,N35503,N35504);
and and21292(N35502,N35505,R0);
and and21297(N35511,N35513,N35514);
and and21298(N35512,N35515,N35516);
and and21303(N35521,N35523,N35524);
and and21304(N35522,N35525,N35526);
and and21309(N35531,N35533,N35534);
and and21310(N35532,N35535,R1);
and and21315(N35541,N35543,N35544);
and and21316(N35542,N35545,N35546);
and and21321(N35551,N35553,N35554);
and and21322(N35552,N35555,N35556);
and and21327(N35561,N35563,N35564);
and and21328(N35562,N35565,R0);
and and21333(N35571,N35573,N35574);
and and21334(N35572,N35575,R0);
and and21339(N35581,N35583,N35584);
and and21340(N35582,N35585,R0);
and and21345(N35591,N35593,N35594);
and and21346(N35592,N35595,R0);
and and21351(N35601,N35603,N35604);
and and21352(N35602,N35605,R0);
and and21357(N35610,N35612,N35613);
and and21358(N35611,N35614,R0);
and and21363(N35619,N35621,N35622);
and and21364(N35620,N35623,N35624);
and and21369(N35628,N35630,N35631);
and and21370(N35629,N35632,N35633);
and and21375(N35637,N35639,N35640);
and and21376(N35638,N35641,N35642);
and and21381(N35646,N35648,N35649);
and and21382(N35647,N35650,N35651);
and and21387(N35655,N35657,N35658);
and and21388(N35656,N35659,R0);
and and21393(N35664,N35666,N35667);
and and21394(N35665,N35668,R0);
and and21399(N35673,N35675,N35676);
and and21400(N35674,N35677,R0);
and and21405(N35682,N35684,N35685);
and and21406(N35683,N35686,R0);
and and21411(N35691,N35693,N35694);
and and21412(N35692,N35695,R0);
and and21417(N35699,N35701,N35702);
and and21418(N35700,N35703,R0);
and and21423(N35707,N35709,N35710);
and and21424(N35708,N35711,R0);
and and21429(N35715,N35717,N35718);
and and21430(N35716,N35719,R0);
and and21435(N35723,N35725,N35726);
and and21436(N35724,N35727,R0);
and and21441(N35731,N35733,N35734);
and and21442(N35732,N35735,N35736);
and and21447(N35739,N35741,N35742);
and and21448(N35740,N35743,R0);
and and21453(N35746,N35748,N35749);
and and21454(N35747,N35750,R0);
and and21459(N35753,N35755,N35756);
and and21460(N35754,N35757,R0);
and and21240(N35414,R0,R1);
and and21241(N35415,R2,N35418);
and and21242(N35416,N35419,N35420);
and and21243(N35417,N35421,N35422);
and and21247(N35426,N35430,N35431);
and and21248(N35427,R2,N35432);
and and21249(N35428,R4,R5);
and and21250(N35429,N35433,N35434);
and and21254(N35438,N35442,N35443);
and and21255(N35439,N35444,R3);
and and21256(N35440,R4,R5);
and and21257(N35441,N35445,R7);
and and21261(N35449,R0,R1);
and and21262(N35450,R2,N35453);
and and21263(N35451,N35454,R5);
and and21264(N35452,N35455,R7);
and and21268(N35459,R0,R1);
and and21269(N35460,R2,R3);
and and21270(N35461,N35463,N35464);
and and21271(N35462,R6,R7);
and and21275(N35468,N35472,R2);
and and21276(N35469,N35473,N35474);
and and21277(N35470,N35475,N35476);
and and21281(N35480,N35484,N35485);
and and21282(N35481,R3,N35486);
and and21283(N35482,N35487,N35488);
and and21287(N35492,N35496,R2);
and and21288(N35493,N35497,N35498);
and and21289(N35494,N35499,R7);
and and21293(N35503,N35506,N35507);
and and21294(N35504,N35508,R5);
and and21295(N35505,N35509,R7);
and and21299(N35513,R1,R2);
and and21300(N35514,R3,N35517);
and and21301(N35515,N35518,N35519);
and and21305(N35523,R2,R3);
and and21306(N35524,N35527,N35528);
and and21307(N35525,R6,N35529);
and and21311(N35533,N35536,R3);
and and21312(N35534,N35537,R5);
and and21313(N35535,N35538,N35539);
and and21317(N35543,R1,R2);
and and21318(N35544,N35547,N35548);
and and21319(N35545,R5,N35549);
and and21323(N35553,N35557,R3);
and and21324(N35554,N35558,R5);
and and21325(N35555,R6,N35559);
and and21329(N35563,R1,N35566);
and and21330(N35564,R4,N35567);
and and21331(N35565,N35568,N35569);
and and21335(N35573,R1,N35576);
and and21336(N35574,N35577,N35578);
and and21337(N35575,N35579,R7);
and and21341(N35583,N35586,R2);
and and21342(N35584,N35587,R5);
and and21343(N35585,N35588,N35589);
and and21347(N35593,N35596,R2);
and and21348(N35594,N35597,R4);
and and21349(N35595,N35598,N35599);
and and21353(N35603,R1,N35606);
and and21354(N35604,R3,N35607);
and and21355(N35605,R6,N35608);
and and21359(N35612,N35615,R2);
and and21360(N35613,N35616,R5);
and and21361(N35614,R6,N35617);
and and21365(N35621,N35625,R2);
and and21366(N35622,R3,R4);
and and21367(N35623,N35626,R6);
and and21371(N35630,N35634,R2);
and and21372(N35631,R3,N35635);
and and21373(N35632,R6,R7);
and and21377(N35639,N35643,R2);
and and21378(N35640,R3,N35644);
and and21379(N35641,R5,R6);
and and21383(N35648,R1,R2);
and and21384(N35649,R3,R4);
and and21385(N35650,N35652,N35653);
and and21389(N35657,N35660,N35661);
and and21390(N35658,R3,N35662);
and and21391(N35659,R5,R6);
and and21395(N35666,R1,R3);
and and21396(N35667,R4,N35669);
and and21397(N35668,N35670,N35671);
and and21401(N35675,N35678,R2);
and and21402(N35676,N35679,R4);
and and21403(N35677,N35680,R7);
and and21407(N35684,R2,N35687);
and and21408(N35685,R4,N35688);
and and21409(N35686,N35689,R7);
and and21413(N35693,R1,N35696);
and and21414(N35694,R3,R4);
and and21415(N35695,N35697,R7);
and and21419(N35701,R1,N35704);
and and21420(N35702,R4,R5);
and and21421(N35703,N35705,R7);
and and21425(N35709,R1,R3);
and and21426(N35710,N35712,R5);
and and21427(N35711,R6,N35713);
and and21431(N35717,N35720,R3);
and and21432(N35718,R4,N35721);
and and21433(N35719,R6,R7);
and and21437(N35725,R1,N35728);
and and21438(N35726,R3,R5);
and and21439(N35727,N35729,R7);
and and21443(N35733,R2,R3);
and and21444(N35734,N35737,R5);
and and21445(N35735,R6,R7);
and and21449(N35741,R1,R2);
and and21450(N35742,N35744,R4);
and and21451(N35743,R5,R6);
and and21455(N35748,R1,R3);
and and21456(N35749,R4,R5);
and and21457(N35750,N35751,R7);
and and21461(N35755,N35758,R2);
and and21462(N35756,R3,R4);
and and21463(N35757,R6,R7);
and and21464(N35772,N35773,N35774);
and and21471(N35785,N35786,N35787);
and and21478(N35798,N35799,N35800);
and and21485(N35810,N35811,N35812);
and and21492(N35822,N35823,N35824);
and and21499(N35834,N35835,N35836);
and and21506(N35846,N35847,N35848);
and and21513(N35857,N35858,N35859);
and and21520(N35868,N35869,N35870);
and and21527(N35878,N35879,N35880);
and and21534(N35887,N35888,N35889);
and and21541(N35896,N35897,N35898);
and and21548(N35905,N35906,N35907);
and and21554(N35914,N35915,N35916);
and and21465(N35773,N35775,N35776);
and and21466(N35774,N35777,N35778);
and and21472(N35786,N35788,N35789);
and and21473(N35787,N35790,N35791);
and and21479(N35799,N35801,N35802);
and and21480(N35800,N35803,N35804);
and and21486(N35811,N35813,N35814);
and and21487(N35812,N35815,N35816);
and and21493(N35823,N35825,N35826);
and and21494(N35824,N35827,N35828);
and and21500(N35835,N35837,N35838);
and and21501(N35836,N35839,N35840);
and and21507(N35847,N35849,N35850);
and and21508(N35848,N35851,N35852);
and and21514(N35858,N35860,N35861);
and and21515(N35859,N35862,N35863);
and and21521(N35869,N35871,N35872);
and and21522(N35870,N35873,N35874);
and and21528(N35879,N35881,N35882);
and and21529(N35880,N35883,N35884);
and and21535(N35888,N35890,N35891);
and and21536(N35889,N35892,N35893);
and and21542(N35897,N35899,N35900);
and and21543(N35898,N35901,N35902);
and and21549(N35906,N35908,N35909);
and and21550(N35907,N35910,N35911);
and and21555(N35915,N35917,N35918);
and and21556(N35916,N35919,N35920);
and and21467(N35775,R0,N35779);
and and21468(N35776,N35780,R3);
and and21469(N35777,N35781,N35782);
and and21470(N35778,N35783,N35784);
and and21474(N35788,R0,N35792);
and and21475(N35789,N35793,N35794);
and and21476(N35790,N35795,N35796);
and and21477(N35791,R6,N35797);
and and21481(N35801,R0,N35805);
and and21482(N35802,R2,N35806);
and and21483(N35803,N35807,N35808);
and and21484(N35804,N35809,R7);
and and21488(N35813,N35817,N35818);
and and21489(N35814,R2,R3);
and and21490(N35815,N35819,R5);
and and21491(N35816,N35820,N35821);
and and21495(N35825,N35829,N35830);
and and21496(N35826,N35831,R3);
and and21497(N35827,N35832,R5);
and and21498(N35828,N35833,R7);
and and21502(N35837,N35841,N35842);
and and21503(N35838,R2,N35843);
and and21504(N35839,N35844,N35845);
and and21505(N35840,R6,R7);
and and21509(N35849,R0,N35853);
and and21510(N35850,N35854,R3);
and and21511(N35851,R4,R5);
and and21512(N35852,N35855,N35856);
and and21516(N35860,R0,N35864);
and and21517(N35861,N35865,R3);
and and21518(N35862,R4,N35866);
and and21519(N35863,N35867,R7);
and and21523(N35871,R0,R1);
and and21524(N35872,R2,N35875);
and and21525(N35873,R4,N35876);
and and21526(N35874,R6,N35877);
and and21530(N35881,R0,N35885);
and and21531(N35882,R2,R3);
and and21532(N35883,N35886,R5);
and and21533(N35884,R6,R7);
and and21537(N35890,R0,R1);
and and21538(N35891,R2,R3);
and and21539(N35892,R4,N35894);
and and21540(N35893,N35895,R7);
and and21544(N35899,R0,R1);
and and21545(N35900,N35903,R3);
and and21546(N35901,R4,R5);
and and21547(N35902,R6,N35904);
and and21551(N35908,R1,N35912);
and and21552(N35909,R3,N35913);
and and21553(N35910,R5,R6);
and and21557(N35917,R1,R2);
and and21558(N35918,N35921,R4);
and and21559(N35919,R6,R7);
and and21560(N35966,N35967,N35968);
and and21567(N35979,N35980,N35981);
and and21574(N35991,N35992,N35993);
and and21581(N36003,N36004,N36005);
and and21588(N36014,N36015,N36016);
and and21595(N36024,N36025,N36026);
and and21602(N36033,N36034,N36035);
and and21608(N36045,N36046,N36047);
and and21614(N36057,N36058,N36059);
and and21620(N36068,N36069,N36070);
and and21626(N36079,N36080,N36081);
and and21632(N36089,N36090,N36091);
and and21638(N36099,N36100,N36101);
and and21644(N36109,N36110,N36111);
and and21650(N36119,N36120,N36121);
and and21656(N36129,N36130,N36131);
and and21662(N36139,N36140,N36141);
and and21668(N36149,N36150,N36151);
and and21674(N36159,N36160,N36161);
and and21680(N36169,N36170,N36171);
and and21686(N36179,N36180,N36181);
and and21692(N36189,N36190,N36191);
and and21698(N36199,N36200,N36201);
and and21704(N36209,N36210,N36211);
and and21710(N36218,N36219,N36220);
and and21716(N36227,N36228,N36229);
and and21722(N36236,N36237,N36238);
and and21728(N36245,N36246,N36247);
and and21734(N36254,N36255,N36256);
and and21740(N36262,N36263,N36264);
and and21746(N36270,N36271,N36272);
and and21752(N36278,N36279,N36280);
and and21758(N36286,N36287,N36288);
and and21764(N36294,N36295,N36296);
and and21770(N36302,N36303,N36304);
and and21776(N36310,N36311,N36312);
and and21782(N36318,N36319,N36320);
and and21788(N36326,N36327,N36328);
and and21794(N36334,N36335,N36336);
and and21800(N36342,N36343,N36344);
and and21806(N36350,N36351,N36352);
and and21812(N36358,N36359,N36360);
and and21818(N36365,N36366,N36367);
and and21824(N36372,N36373,N36374);
and and21830(N36379,N36380,N36381);
and and21561(N35967,N35969,N35970);
and and21562(N35968,N35971,N35972);
and and21568(N35980,N35982,N35983);
and and21569(N35981,N35984,N35985);
and and21575(N35992,N35994,N35995);
and and21576(N35993,N35996,N35997);
and and21582(N36004,N36006,N36007);
and and21583(N36005,N36008,N36009);
and and21589(N36015,N36017,N36018);
and and21590(N36016,N36019,N36020);
and and21596(N36025,N36027,N36028);
and and21597(N36026,N36029,N36030);
and and21603(N36034,N36036,N36037);
and and21604(N36035,N36038,N36039);
and and21609(N36046,N36048,N36049);
and and21610(N36047,N36050,N36051);
and and21615(N36058,N36060,N36061);
and and21616(N36059,N36062,N36063);
and and21621(N36069,N36071,N36072);
and and21622(N36070,N36073,N36074);
and and21627(N36080,N36082,N36083);
and and21628(N36081,N36084,R0);
and and21633(N36090,N36092,N36093);
and and21634(N36091,N36094,N36095);
and and21639(N36100,N36102,N36103);
and and21640(N36101,N36104,N36105);
and and21645(N36110,N36112,N36113);
and and21646(N36111,N36114,N36115);
and and21651(N36120,N36122,N36123);
and and21652(N36121,N36124,N36125);
and and21657(N36130,N36132,N36133);
and and21658(N36131,N36134,R0);
and and21663(N36140,N36142,N36143);
and and21664(N36141,N36144,R0);
and and21669(N36150,N36152,N36153);
and and21670(N36151,N36154,R0);
and and21675(N36160,N36162,N36163);
and and21676(N36161,N36164,N36165);
and and21681(N36170,N36172,N36173);
and and21682(N36171,N36174,N36175);
and and21687(N36180,N36182,N36183);
and and21688(N36181,N36184,R0);
and and21693(N36190,N36192,N36193);
and and21694(N36191,N36194,R0);
and and21699(N36200,N36202,N36203);
and and21700(N36201,N36204,N36205);
and and21705(N36210,N36212,N36213);
and and21706(N36211,N36214,R0);
and and21711(N36219,N36221,N36222);
and and21712(N36220,N36223,R0);
and and21717(N36228,N36230,N36231);
and and21718(N36229,N36232,N36233);
and and21723(N36237,N36239,N36240);
and and21724(N36238,N36241,N36242);
and and21729(N36246,N36248,N36249);
and and21730(N36247,N36250,R0);
and and21735(N36255,N36257,N36258);
and and21736(N36256,N36259,R1);
and and21741(N36263,N36265,N36266);
and and21742(N36264,N36267,R0);
and and21747(N36271,N36273,N36274);
and and21748(N36272,N36275,R0);
and and21753(N36279,N36281,N36282);
and and21754(N36280,N36283,R0);
and and21759(N36287,N36289,N36290);
and and21760(N36288,N36291,N36292);
and and21765(N36295,N36297,N36298);
and and21766(N36296,N36299,N36300);
and and21771(N36303,N36305,N36306);
and and21772(N36304,N36307,R0);
and and21777(N36311,N36313,N36314);
and and21778(N36312,N36315,R0);
and and21783(N36319,N36321,N36322);
and and21784(N36320,N36323,R0);
and and21789(N36327,N36329,N36330);
and and21790(N36328,N36331,R0);
and and21795(N36335,N36337,N36338);
and and21796(N36336,N36339,R0);
and and21801(N36343,N36345,N36346);
and and21802(N36344,N36347,R0);
and and21807(N36351,N36353,N36354);
and and21808(N36352,N36355,R0);
and and21813(N36359,N36361,N36362);
and and21814(N36360,N36363,R0);
and and21819(N36366,N36368,N36369);
and and21820(N36367,N36370,R0);
and and21825(N36373,N36375,N36376);
and and21826(N36374,N36377,R0);
and and21831(N36380,N36382,N36383);
and and21832(N36381,R1,N36384);
and and21563(N35969,R0,N35973);
and and21564(N35970,N35974,N35975);
and and21565(N35971,N35976,N35977);
and and21566(N35972,R6,N35978);
and and21570(N35982,R0,R1);
and and21571(N35983,R2,N35986);
and and21572(N35984,N35987,N35988);
and and21573(N35985,N35989,N35990);
and and21577(N35994,N35998,N35999);
and and21578(N35995,R2,N36000);
and and21579(N35996,R4,R5);
and and21580(N35997,N36001,N36002);
and and21584(N36006,R0,N36010);
and and21585(N36007,N36011,R3);
and and21586(N36008,R4,R5);
and and21587(N36009,N36012,N36013);
and and21591(N36017,R0,R1);
and and21592(N36018,R2,N36021);
and and21593(N36019,N36022,R5);
and and21594(N36020,N36023,R7);
and and21598(N36027,R0,R1);
and and21599(N36028,R2,R3);
and and21600(N36029,N36031,N36032);
and and21601(N36030,R6,R7);
and and21605(N36036,N36040,R2);
and and21606(N36037,N36041,N36042);
and and21607(N36038,N36043,N36044);
and and21611(N36048,N36052,R3);
and and21612(N36049,N36053,N36054);
and and21613(N36050,N36055,N36056);
and and21617(N36060,N36064,N36065);
and and21618(N36061,R3,N36066);
and and21619(N36062,N36067,R7);
and and21623(N36071,N36075,R2);
and and21624(N36072,N36076,N36077);
and and21625(N36073,N36078,R7);
and and21629(N36082,N36085,N36086);
and and21630(N36083,N36087,R5);
and and21631(N36084,N36088,R7);
and and21635(N36092,R1,R2);
and and21636(N36093,R3,N36096);
and and21637(N36094,N36097,N36098);
and and21641(N36102,R2,R3);
and and21642(N36103,N36106,N36107);
and and21643(N36104,R6,N36108);
and and21647(N36112,R1,R2);
and and21648(N36113,N36116,N36117);
and and21649(N36114,R5,N36118);
and and21653(N36122,N36126,R3);
and and21654(N36123,N36127,R5);
and and21655(N36124,R6,N36128);
and and21659(N36132,R1,N36135);
and and21660(N36133,R4,N36136);
and and21661(N36134,N36137,N36138);
and and21665(N36142,R1,N36145);
and and21666(N36143,N36146,N36147);
and and21667(N36144,N36148,R7);
and and21671(N36152,N36155,R2);
and and21672(N36153,N36156,N36157);
and and21673(N36154,N36158,R7);
and and21677(N36162,R2,R3);
and and21678(N36163,N36166,R5);
and and21679(N36164,N36167,N36168);
and and21683(N36172,N36176,R2);
and and21684(N36173,N36177,N36178);
and and21685(N36174,R6,R7);
and and21689(N36182,N36185,R2);
and and21690(N36183,N36186,N36187);
and and21691(N36184,R5,N36188);
and and21695(N36192,N36195,R2);
and and21696(N36193,N36196,R4);
and and21697(N36194,N36197,N36198);
and and21701(N36202,N36206,N36207);
and and21702(N36203,R3,R5);
and and21703(N36204,N36208,R7);
and and21707(N36212,R1,N36215);
and and21708(N36213,R3,N36216);
and and21709(N36214,R6,N36217);
and and21713(N36221,N36224,R3);
and and21714(N36222,R4,N36225);
and and21715(N36223,N36226,R7);
and and21719(N36230,N36234,R2);
and and21720(N36231,R3,R4);
and and21721(N36232,N36235,R6);
and and21725(N36239,N36243,R2);
and and21726(N36240,R3,N36244);
and and21727(N36241,R5,R6);
and and21731(N36248,N36251,R2);
and and21732(N36249,N36252,R4);
and and21733(N36250,N36253,R7);
and and21737(N36257,R2,R3);
and and21738(N36258,R4,N36260);
and and21739(N36259,N36261,R7);
and and21743(N36265,R1,N36268);
and and21744(N36266,R4,R5);
and and21745(N36267,N36269,R7);
and and21749(N36273,N36276,R3);
and and21750(N36274,R4,N36277);
and and21751(N36275,R6,R7);
and and21755(N36281,N36284,R3);
and and21756(N36282,N36285,R5);
and and21757(N36283,R6,R7);
and and21761(N36289,R1,R2);
and and21762(N36290,N36293,R4);
and and21763(N36291,R6,R7);
and and21767(N36297,R1,R3);
and and21768(N36298,N36301,R5);
and and21769(N36299,R6,R7);
and and21773(N36305,R1,R2);
and and21774(N36306,N36308,R4);
and and21775(N36307,R6,N36309);
and and21779(N36313,R1,R2);
and and21780(N36314,R3,R4);
and and21781(N36315,N36316,N36317);
and and21785(N36321,R1,R2);
and and21786(N36322,R4,N36324);
and and21787(N36323,N36325,R7);
and and21791(N36329,R2,N36332);
and and21792(N36330,R4,R5);
and and21793(N36331,R6,N36333);
and and21797(N36337,R1,N36340);
and and21798(N36338,R3,R5);
and and21799(N36339,N36341,R7);
and and21803(N36345,R1,N36348);
and and21804(N36346,R3,R4);
and and21805(N36347,R6,N36349);
and and21809(N36353,R1,R3);
and and21810(N36354,N36356,R5);
and and21811(N36355,R6,N36357);
and and21815(N36361,R1,R2);
and and21816(N36362,N36364,R4);
and and21817(N36363,R5,R6);
and and21821(N36368,R1,R3);
and and21822(N36369,R4,R5);
and and21823(N36370,N36371,R7);
and and21827(N36375,N36378,R2);
and and21828(N36376,R3,R4);
and and21829(N36377,R6,R7);
and and21833(N36382,R3,N36385);
and and21834(N36383,R5,N36386);
and and21835(N36408,N36409,N36410);
and and21842(N36422,N36423,N36424);
and and21849(N36435,N36436,N36437);
and and21856(N36448,N36449,N36450);
and and21863(N36461,N36462,N36463);
and and21870(N36473,N36474,N36475);
and and21877(N36485,N36486,N36487);
and and21884(N36496,N36497,N36498);
and and21891(N36507,N36508,N36509);
and and21898(N36518,N36519,N36520);
and and21905(N36529,N36530,N36531);
and and21912(N36540,N36541,N36542);
and and21919(N36551,N36552,N36553);
and and21926(N36561,N36562,N36563);
and and21933(N36569,N36570,N36571);
and and21939(N36580,N36581,N36582);
and and21945(N36591,N36592,N36593);
and and21951(N36601,N36602,N36603);
and and21957(N36611,N36612,N36613);
and and21963(N36620,N36621,N36622);
and and21969(N36629,N36630,N36631);
and and21975(N36638,N36639,N36640);
and and21836(N36409,N36411,N36412);
and and21837(N36410,N36413,N36414);
and and21843(N36423,N36425,N36426);
and and21844(N36424,N36427,N36428);
and and21850(N36436,N36438,N36439);
and and21851(N36437,N36440,N36441);
and and21857(N36449,N36451,N36452);
and and21858(N36450,N36453,N36454);
and and21864(N36462,N36464,N36465);
and and21865(N36463,N36466,N36467);
and and21871(N36474,N36476,N36477);
and and21872(N36475,N36478,N36479);
and and21878(N36486,N36488,N36489);
and and21879(N36487,N36490,N36491);
and and21885(N36497,N36499,N36500);
and and21886(N36498,N36501,N36502);
and and21892(N36508,N36510,N36511);
and and21893(N36509,N36512,N36513);
and and21899(N36519,N36521,N36522);
and and21900(N36520,N36523,N36524);
and and21906(N36530,N36532,N36533);
and and21907(N36531,N36534,N36535);
and and21913(N36541,N36543,N36544);
and and21914(N36542,N36545,N36546);
and and21920(N36552,N36554,N36555);
and and21921(N36553,N36556,N36557);
and and21927(N36562,N36564,N36565);
and and21928(N36563,N36566,N36567);
and and21934(N36570,N36572,N36573);
and and21935(N36571,N36574,N36575);
and and21940(N36581,N36583,N36584);
and and21941(N36582,N36585,N36586);
and and21946(N36592,N36594,N36595);
and and21947(N36593,N36596,R1);
and and21952(N36602,N36604,N36605);
and and21953(N36603,N36606,N36607);
and and21958(N36612,N36614,N36615);
and and21959(N36613,N36616,N36617);
and and21964(N36621,N36623,N36624);
and and21965(N36622,N36625,R0);
and and21970(N36630,N36632,N36633);
and and21971(N36631,N36634,R0);
and and21976(N36639,N36641,N36642);
and and21977(N36640,N36643,R0);
and and21838(N36411,N36415,N36416);
and and21839(N36412,N36417,N36418);
and and21840(N36413,N36419,N36420);
and and21841(N36414,R6,N36421);
and and21845(N36425,N36429,R1);
and and21846(N36426,N36430,N36431);
and and21847(N36427,N36432,N36433);
and and21848(N36428,N36434,R7);
and and21852(N36438,N36442,N36443);
and and21853(N36439,N36444,N36445);
and and21854(N36440,R4,R5);
and and21855(N36441,N36446,N36447);
and and21859(N36451,N36455,R1);
and and21860(N36452,N36456,N36457);
and and21861(N36453,N36458,R5);
and and21862(N36454,N36459,N36460);
and and21866(N36464,R0,N36468);
and and21867(N36465,N36469,R3);
and and21868(N36466,N36470,N36471);
and and21869(N36467,N36472,R7);
and and21873(N36476,N36480,R1);
and and21874(N36477,N36481,R3);
and and21875(N36478,N36482,N36483);
and and21876(N36479,R6,N36484);
and and21880(N36488,R0,R1);
and and21881(N36489,N36492,N36493);
and and21882(N36490,R4,N36494);
and and21883(N36491,N36495,R7);
and and21887(N36499,R0,R1);
and and21888(N36500,R2,N36503);
and and21889(N36501,N36504,R5);
and and21890(N36502,N36505,N36506);
and and21894(N36510,N36514,R1);
and and21895(N36511,R2,R3);
and and21896(N36512,N36515,R5);
and and21897(N36513,N36516,N36517);
and and21901(N36521,R0,R1);
and and21902(N36522,R2,R3);
and and21903(N36523,N36525,N36526);
and and21904(N36524,N36527,N36528);
and and21908(N36532,N36536,N36537);
and and21909(N36533,R2,N36538);
and and21910(N36534,R4,N36539);
and and21911(N36535,R6,R7);
and and21915(N36543,R0,R1);
and and21916(N36544,N36547,N36548);
and and21917(N36545,R4,R5);
and and21918(N36546,N36549,N36550);
and and21922(N36554,R0,N36558);
and and21923(N36555,R2,R3);
and and21924(N36556,N36559,R5);
and and21925(N36557,N36560,R7);
and and21929(N36564,R0,R1);
and and21930(N36565,N36568,R3);
and and21931(N36566,R4,R5);
and and21932(N36567,R6,R7);
and and21936(N36572,N36576,R3);
and and21937(N36573,R4,N36577);
and and21938(N36574,N36578,N36579);
and and21942(N36583,N36587,R3);
and and21943(N36584,R4,N36588);
and and21944(N36585,N36589,N36590);
and and21948(N36594,R2,N36597);
and and21949(N36595,R4,N36598);
and and21950(N36596,N36599,N36600);
and and21954(N36604,N36608,N36609);
and and21955(N36605,R3,R4);
and and21956(N36606,R6,N36610);
and and21960(N36614,R1,N36618);
and and21961(N36615,R3,R4);
and and21962(N36616,R5,N36619);
and and21966(N36623,N36626,N36627);
and and21967(N36624,N36628,R4);
and and21968(N36625,R5,R6);
and and21972(N36632,N36635,R2);
and and21973(N36633,R3,N36636);
and and21974(N36634,R6,N36637);
and and21978(N36641,N36644,R2);
and and21979(N36642,R3,R4);
and and21980(N36643,R6,N36645);
and and21981(N36693,N36694,N36695);
and and21988(N36707,N36708,N36709);
and and21995(N36719,N36720,N36721);
and and22002(N36731,N36732,N36733);
and and22009(N36742,N36743,N36744);
and and22016(N36752,N36753,N36754);
and and22022(N36764,N36765,N36766);
and and22028(N36776,N36777,N36778);
and and22034(N36788,N36789,N36790);
and and22040(N36799,N36800,N36801);
and and22046(N36810,N36811,N36812);
and and22052(N36821,N36822,N36823);
and and22058(N36832,N36833,N36834);
and and22064(N36842,N36843,N36844);
and and22070(N36852,N36853,N36854);
and and22076(N36862,N36863,N36864);
and and22082(N36872,N36873,N36874);
and and22088(N36882,N36883,N36884);
and and22094(N36892,N36893,N36894);
and and22100(N36902,N36903,N36904);
and and22106(N36912,N36913,N36914);
and and22112(N36922,N36923,N36924);
and and22118(N36932,N36933,N36934);
and and22124(N36942,N36943,N36944);
and and22130(N36952,N36953,N36954);
and and22136(N36961,N36962,N36963);
and and22142(N36970,N36971,N36972);
and and22148(N36979,N36980,N36981);
and and22154(N36988,N36989,N36990);
and and22160(N36997,N36998,N36999);
and and22166(N37006,N37007,N37008);
and and22172(N37015,N37016,N37017);
and and22178(N37023,N37024,N37025);
and and22184(N37031,N37032,N37033);
and and22190(N37039,N37040,N37041);
and and22196(N37047,N37048,N37049);
and and22202(N37055,N37056,N37057);
and and22208(N37063,N37064,N37065);
and and22214(N37071,N37072,N37073);
and and22220(N37079,N37080,N37081);
and and22226(N37087,N37088,N37089);
and and22232(N37095,N37096,N37097);
and and22238(N37103,N37104,N37105);
and and22244(N37111,N37112,N37113);
and and22250(N37118,N37119,N37120);
and and22256(N37125,N37126,N37127);
and and22262(N37132,N37133,N37134);
and and22268(N37139,N37140,N37141);
and and21982(N36694,N36696,N36697);
and and21983(N36695,N36698,N36699);
and and21989(N36708,N36710,N36711);
and and21990(N36709,N36712,N36713);
and and21996(N36720,N36722,N36723);
and and21997(N36721,N36724,N36725);
and and22003(N36732,N36734,N36735);
and and22004(N36733,N36736,N36737);
and and22010(N36743,N36745,N36746);
and and22011(N36744,N36747,N36748);
and and22017(N36753,N36755,N36756);
and and22018(N36754,N36757,N36758);
and and22023(N36765,N36767,N36768);
and and22024(N36766,N36769,R0);
and and22029(N36777,N36779,N36780);
and and22030(N36778,N36781,N36782);
and and22035(N36789,N36791,N36792);
and and22036(N36790,N36793,N36794);
and and22041(N36800,N36802,N36803);
and and22042(N36801,N36804,N36805);
and and22047(N36811,N36813,N36814);
and and22048(N36812,N36815,N36816);
and and22053(N36822,N36824,N36825);
and and22054(N36823,N36826,N36827);
and and22059(N36833,N36835,N36836);
and and22060(N36834,N36837,N36838);
and and22065(N36843,N36845,N36846);
and and22066(N36844,N36847,N36848);
and and22071(N36853,N36855,N36856);
and and22072(N36854,N36857,N36858);
and and22077(N36863,N36865,N36866);
and and22078(N36864,N36867,N36868);
and and22083(N36873,N36875,N36876);
and and22084(N36874,N36877,N36878);
and and22089(N36883,N36885,N36886);
and and22090(N36884,N36887,N36888);
and and22095(N36893,N36895,N36896);
and and22096(N36894,N36897,R0);
and and22101(N36903,N36905,N36906);
and and22102(N36904,N36907,R0);
and and22107(N36913,N36915,N36916);
and and22108(N36914,N36917,R0);
and and22113(N36923,N36925,N36926);
and and22114(N36924,N36927,R0);
and and22119(N36933,N36935,N36936);
and and22120(N36934,N36937,R0);
and and22125(N36943,N36945,N36946);
and and22126(N36944,N36947,R0);
and and22131(N36953,N36955,N36956);
and and22132(N36954,N36957,N36958);
and and22137(N36962,N36964,N36965);
and and22138(N36963,N36966,R1);
and and22143(N36971,N36973,N36974);
and and22144(N36972,N36975,N36976);
and and22149(N36980,N36982,N36983);
and and22150(N36981,N36984,N36985);
and and22155(N36989,N36991,N36992);
and and22156(N36990,N36993,N36994);
and and22161(N36998,N37000,N37001);
and and22162(N36999,N37002,N37003);
and and22167(N37007,N37009,N37010);
and and22168(N37008,N37011,R0);
and and22173(N37016,N37018,N37019);
and and22174(N37017,N37020,N37021);
and and22179(N37024,N37026,N37027);
and and22180(N37025,N37028,R0);
and and22185(N37032,N37034,N37035);
and and22186(N37033,N37036,R0);
and and22191(N37040,N37042,N37043);
and and22192(N37041,N37044,R0);
and and22197(N37048,N37050,N37051);
and and22198(N37049,N37052,R0);
and and22203(N37056,N37058,N37059);
and and22204(N37057,N37060,N37061);
and and22209(N37064,N37066,N37067);
and and22210(N37065,N37068,R0);
and and22215(N37072,N37074,N37075);
and and22216(N37073,N37076,R0);
and and22221(N37080,N37082,N37083);
and and22222(N37081,N37084,N37085);
and and22227(N37088,N37090,N37091);
and and22228(N37089,N37092,N37093);
and and22233(N37096,N37098,N37099);
and and22234(N37097,N37100,R0);
and and22239(N37104,N37106,N37107);
and and22240(N37105,N37108,R0);
and and22245(N37112,N37114,N37115);
and and22246(N37113,N37116,N37117);
and and22251(N37119,N37121,N37122);
and and22252(N37120,N37123,N37124);
and and22257(N37126,N37128,N37129);
and and22258(N37127,N37130,N37131);
and and22263(N37133,N37135,N37136);
and and22264(N37134,N37137,R0);
and and22269(N37140,N37142,N37143);
and and22270(N37141,N37144,R1);
and and21984(N36696,N36700,N36701);
and and21985(N36697,N36702,N36703);
and and21986(N36698,R4,N36704);
and and21987(N36699,N36705,N36706);
and and21991(N36710,R0,N36714);
and and21992(N36711,N36715,R3);
and and21993(N36712,N36716,R5);
and and21994(N36713,N36717,N36718);
and and21998(N36722,R0,R1);
and and21999(N36723,N36726,N36727);
and and22000(N36724,N36728,R5);
and and22001(N36725,N36729,N36730);
and and22005(N36734,R0,N36738);
and and22006(N36735,R2,N36739);
and and22007(N36736,N36740,R5);
and and22008(N36737,N36741,R7);
and and22012(N36745,R0,R1);
and and22013(N36746,R2,R3);
and and22014(N36747,N36749,N36750);
and and22015(N36748,N36751,R7);
and and22019(N36755,R1,N36759);
and and22020(N36756,N36760,N36761);
and and22021(N36757,N36762,N36763);
and and22025(N36767,N36770,N36771);
and and22026(N36768,N36772,N36773);
and and22027(N36769,N36774,N36775);
and and22031(N36779,N36783,N36784);
and and22032(N36780,N36785,N36786);
and and22033(N36781,N36787,R7);
and and22037(N36791,N36795,R2);
and and22038(N36792,N36796,N36797);
and and22039(N36793,R6,N36798);
and and22043(N36802,R2,R3);
and and22044(N36803,N36806,N36807);
and and22045(N36804,N36808,N36809);
and and22049(N36813,N36817,R2);
and and22050(N36814,N36818,N36819);
and and22051(N36815,R5,N36820);
and and22055(N36824,R1,N36828);
and and22056(N36825,R3,N36829);
and and22057(N36826,N36830,N36831);
and and22061(N36835,R1,R2);
and and22062(N36836,N36839,N36840);
and and22063(N36837,N36841,R7);
and and22067(N36845,N36849,R3);
and and22068(N36846,R4,R5);
and and22069(N36847,N36850,N36851);
and and22073(N36855,N36859,N36860);
and and22074(N36856,R4,R5);
and and22075(N36857,N36861,R7);
and and22079(N36865,N36869,R2);
and and22080(N36866,R3,N36870);
and and22081(N36867,N36871,R7);
and and22085(N36875,N36879,R3);
and and22086(N36876,R4,N36880);
and and22087(N36877,N36881,R7);
and and22091(N36885,R1,N36889);
and and22092(N36886,N36890,R5);
and and22093(N36887,N36891,R7);
and and22097(N36895,N36898,N36899);
and and22098(N36896,N36900,R4);
and and22099(N36897,N36901,R7);
and and22103(N36905,N36908,N36909);
and and22104(N36906,N36910,N36911);
and and22105(N36907,R5,R6);
and and22109(N36915,N36918,N36919);
and and22110(N36916,R4,N36920);
and and22111(N36917,R6,N36921);
and and22115(N36925,N36928,N36929);
and and22116(N36926,N36930,N36931);
and and22117(N36927,R6,R7);
and and22121(N36935,N36938,N36939);
and and22122(N36936,R4,R5);
and and22123(N36937,N36940,N36941);
and and22127(N36945,N36948,N36949);
and and22128(N36946,R4,N36950);
and and22129(N36947,R6,N36951);
and and22133(N36955,N36959,R2);
and and22134(N36956,R4,R5);
and and22135(N36957,N36960,R7);
and and22139(N36964,R2,N36967);
and and22140(N36965,R4,R5);
and and22141(N36966,N36968,N36969);
and and22145(N36973,N36977,N36978);
and and22146(N36974,R3,R5);
and and22147(N36975,R6,R7);
and and22151(N36982,R1,R2);
and and22152(N36983,N36986,R5);
and and22153(N36984,N36987,R7);
and and22157(N36991,R1,R2);
and and22158(N36992,N36995,R4);
and and22159(N36993,N36996,R7);
and and22163(N37000,N37004,R2);
and and22164(N37001,N37005,R4);
and and22165(N37002,R5,R6);
and and22169(N37009,N37012,R3);
and and22170(N37010,N37013,N37014);
and and22171(N37011,R6,R7);
and and22175(N37018,R1,R2);
and and22176(N37019,R3,R5);
and and22177(N37020,R6,N37022);
and and22181(N37026,R1,R2);
and and22182(N37027,N37029,N37030);
and and22183(N37028,R5,R6);
and and22187(N37034,R1,R2);
and and22188(N37035,R3,R5);
and and22189(N37036,N37037,N37038);
and and22193(N37042,N37045,R2);
and and22194(N37043,R3,R4);
and and22195(N37044,N37046,R7);
and and22199(N37050,R1,R3);
and and22200(N37051,R4,R5);
and and22201(N37052,N37053,N37054);
and and22205(N37058,R1,R2);
and and22206(N37059,R3,R4);
and and22207(N37060,N37062,R6);
and and22211(N37066,R1,R2);
and and22212(N37067,N37069,N37070);
and and22213(N37068,R6,R7);
and and22217(N37074,R1,N37077);
and and22218(N37075,R3,N37078);
and and22219(N37076,R6,R7);
and and22223(N37082,R2,N37086);
and and22224(N37083,R4,R5);
and and22225(N37084,R6,R7);
and and22229(N37090,N37094,R3);
and and22230(N37091,R4,R5);
and and22231(N37092,R6,R7);
and and22235(N37098,R1,N37101);
and and22236(N37099,R3,N37102);
and and22237(N37100,R6,R7);
and and22241(N37106,R1,R2);
and and22242(N37107,N37109,R4);
and and22243(N37108,R5,N37110);
and and22247(N37114,R1,R3);
and and22248(N37115,R4,R5);
and and22249(N37116,R6,R7);
and and22253(N37121,R2,R3);
and and22254(N37122,R4,R5);
and and22255(N37123,R6,R7);
and and22259(N37128,R1,R2);
and and22260(N37129,R3,R4);
and and22261(N37130,R5,R7);
and and22265(N37135,R1,R2);
and and22266(N37136,R3,R4);
and and22267(N37137,R5,N37138);
and and22271(N37142,R2,R3);
and and22272(N37143,R4,N37145);
and and22273(N37144,R6,R7);

or or0(N0,N1,N2);
or or1(N1,N3,N4);
or or2(N2,N5,N6);
or or3(N3,N7,N8);
or or4(N4,N9,N10);
or or5(N5,N11,N12);
or or6(N6,N13,N14);
or or7(N7,N15,N16);
or or8(N8,N17,N18);
or or9(N9,N19,N20);
or or10(N10,N21,N22);
or or11(N11,N23,N24);
or or12(N12,N25,N26);
or or13(N13,N27,N28);
or or14(N14,N29,N30);
or or15(N15,N31,N32);
or or16(N16,N33,N34);
or or17(N17,N35,N36);
or or18(N18,N37,N38);
or or19(N19,N39,N40);
or or20(N20,N41,N42);
or or21(N21,N43,N44);
or or22(N22,N45,N46);
or or23(N23,N47,N48);
or or24(N24,N49,N50);
or or25(N25,N51,N52);
or or26(N26,N53,N54);
or or27(N27,N55,N56);
or or28(N28,N57,N58);
or or29(N29,N59,N60);
or or30(N30,N61,N62);
or or31(N31,N63,N64);
or or32(N32,N65,N66);
or or33(N33,N67,N68);
or or34(N34,N69,N70);
or or35(N35,N71,N72);
or or36(N36,N73,N74);
or or37(N37,N75,N76);
or or38(N38,N77,N78);
or or39(N39,N79,N80);
or or40(N40,N81,N82);
or or41(N41,N83,N84);
or or42(N42,N85,N86);
or or43(N43,N87,N88);
or or44(N44,N89,N90);
or or45(N45,N91,N92);
or or46(N46,N93,N94);
or or47(N47,N95,N96);
or or48(N48,N97,N98);
or or49(N49,N99,N100);
or or50(N50,N101,N102);
or or51(N51,N103,N104);
or or52(N52,N105,N106);
or or53(N53,N107,N108);
or or54(N54,N109,N110);
or or55(N55,N111,N112);
or or56(N56,N113,N114);
or or57(N57,N115,N116);
or or58(N58,N117,N118);
or or59(N59,N119,N120);
or or60(N60,N121,N122);
or or61(N61,N123,N124);
or or62(N62,N125,N126);
or or63(N63,N127,N128);
or or64(N64,N129,N130);
or or65(N65,N131,N132);
or or66(N66,N133,N134);
or or67(N67,N135,N136);
or or68(N68,N137,N138);
or or69(N69,N139,N140);
or or70(N70,N141,N142);
or or71(N71,N143,N144);
or or72(N72,N145,N146);
or or73(N73,N147,N148);
or or74(N74,N149,N150);
or or75(N75,N151,N152);
or or76(N76,N153,N154);
or or77(N77,N155,N156);
or or78(N78,N157,N158);
or or79(N79,N159,N160);
or or80(N80,N161,N162);
or or81(N81,N163,N164);
or or82(N82,N165,N166);
or or83(N83,N167,N168);
or or84(N84,N169,N170);
or or85(N85,N171,N172);
or or86(N86,N173,N174);
or or87(N87,N175,N176);
or or88(N88,N177,N178);
or or89(N89,N179,N180);
or or90(N90,N181,N182);
or or91(N91,N183,N184);
or or92(N92,N185,N186);
or or93(N93,N187,N188);
or or94(N94,N189,N190);
or or95(N95,N191,N192);
or or96(N96,N193,N194);
or or97(N97,N195,N196);
or or98(N98,N197,N198);
or or99(N99,N199,N200);
or or100(N100,N201,N202);
or or101(N101,N203,N204);
or or102(N102,N205,N206);
or or103(N103,N207,N208);
or or104(N104,N209,N210);
or or105(N105,N211,N212);
or or106(N106,N213,N214);
or or107(N107,N215,N216);
or or108(N108,N217,N218);
or or109(N109,N219,N220);
or or110(N110,N221,N222);
or or111(N111,N223,N224);
or or112(N112,N225,N226);
or or113(N113,N227,N228);
or or114(N114,N229,N230);
or or115(N115,N231,N232);
or or116(N116,N233,N234);
or or117(N117,N235,N236);
or or118(N118,N237,N238);
or or119(N119,N239,N240);
or or120(N120,N241,N242);
or or121(N121,N243,N244);
or or122(N122,N245,N246);
or or123(N123,N247,N248);
or or124(N124,N249,N250);
or or125(N125,N251,N252);
or or126(N126,N253,N254);
or or127(N127,N255,N256);
or or128(N128,N257,N258);
or or129(N129,N259,N260);
or or130(N130,N261,N262);
or or131(N131,N263,N264);
or or132(N132,N265,N266);
or or133(N133,N267,N268);
or or134(N134,N269,N270);
or or135(N135,N271,N272);
or or136(N136,N273,N274);
or or137(N137,N275,N276);
or or138(N138,N277,N278);
or or139(N139,N279,N280);
or or140(N140,N281,N282);
or or141(N141,N283,N284);
or or142(N142,N285,N286);
or or143(N143,N287,N288);
or or144(N144,N289,N290);
or or145(N145,N291,N292);
or or146(N146,N293,N294);
or or147(N147,N295,N296);
or or148(N148,N297,N298);
or or149(N149,N299,N300);
or or150(N150,N301,N302);
or or151(N151,N303,N304);
or or152(N152,N305,N306);
or or153(N153,N307,N308);
or or154(N154,N309,N310);
or or155(N155,N311,N312);
or or156(N156,N313,N314);
or or157(N157,N315,N316);
or or158(N158,N317,N318);
or or159(N159,N319,N320);
or or160(N160,N321,N322);
or or161(N161,N323,N324);
or or162(N162,N325,N326);
or or163(N163,N327,N328);
or or164(N164,N329,N330);
or or165(N165,N331,N332);
or or166(N166,N333,N334);
or or167(N167,N335,N336);
or or168(N168,N337,N338);
or or169(N169,N339,N340);
or or170(N170,N341,N342);
or or171(N171,N343,N344);
or or172(N172,N345,N346);
or or173(N173,N347,N348);
or or174(N174,N349,N350);
or or175(N175,N351,N352);
or or176(N176,N353,N354);
or or177(N177,N355,N356);
or or178(N178,N357,N358);
or or179(N179,N359,N360);
or or180(N180,N361,N362);
or or181(N181,N363,N364);
or or182(N182,N365,N366);
or or183(N183,N367,N368);
or or184(N184,N369,N370);
or or185(N185,N371,N372);
or or186(N186,N373,N374);
or or187(N187,N375,N376);
or or188(N188,N377,N378);
or or189(N189,N379,N380);
or or190(N190,N381,N382);
or or191(N191,N383,N384);
or or192(N192,N385,N386);
or or193(N193,N387,N388);
or or194(N194,N389,N390);
or or195(N195,N391,N392);
or or196(N196,N393,N394);
or or197(N197,N395,N396);
or or198(N198,N397,N398);
or or199(N199,N399,N400);
or or200(N200,N401,N402);
or or201(N201,N403,N404);
or or202(N202,N405,N406);
or or203(N203,N407,N408);
or or204(N204,N409,N410);
or or205(N205,N411,N428);
or or206(N206,N445,N462);
or or207(N207,N479,N496);
or or208(N208,N513,N530);
or or209(N209,N547,N564);
or or210(N210,N581,N598);
or or211(N211,N615,N631);
or or212(N212,N647,N663);
or or213(N213,N679,N695);
or or214(N214,N711,N727);
or or215(N215,N743,N759);
or or216(N216,N775,N791);
or or217(N217,N807,N822);
or or218(N218,N837,N852);
or or219(N219,N867,N882);
or or220(N220,N897,N912);
or or221(N221,N927,N942);
or or222(N222,N957,N972);
or or223(N223,N987,N1002);
or or224(N224,N1017,N1032);
or or225(N225,N1047,N1062);
or or226(N226,N1077,N1092);
or or227(N227,N1107,N1122);
or or228(N228,N1137,N1152);
or or229(N229,N1167,N1182);
or or230(N230,N1197,N1212);
or or231(N231,N1227,N1242);
or or232(N232,N1257,N1272);
or or233(N233,N1287,N1302);
or or234(N234,N1317,N1332);
or or235(N235,N1347,N1361);
or or236(N236,N1375,N1389);
or or237(N237,N1403,N1417);
or or238(N238,N1431,N1445);
or or239(N239,N1459,N1473);
or or240(N240,N1487,N1501);
or or241(N241,N1515,N1529);
or or242(N242,N1543,N1557);
or or243(N243,N1571,N1585);
or or244(N244,N1599,N1613);
or or245(N245,N1627,N1641);
or or246(N246,N1655,N1669);
or or247(N247,N1683,N1697);
or or248(N248,N1711,N1725);
or or249(N249,N1738,N1751);
or or250(N250,N1764,N1777);
or or251(N251,N1790,N1803);
or or252(N252,N1816,N1829);
or or253(N253,N1842,N1855);
or or254(N254,N1868,N1881);
or or255(N255,N1894,N1907);
or or256(N256,N1920,N1933);
or or257(N257,N1946,N1959);
or or258(N258,N1972,N1985);
or or259(N259,N1998,N2011);
or or260(N260,N2024,N2037);
or or261(N261,N2050,N2063);
or or262(N262,N2076,N2089);
or or263(N263,N2102,N2115);
or or264(N264,N2128,N2141);
or or265(N265,N2154,N2167);
or or266(N266,N2180,N2193);
or or267(N267,N2206,N2219);
or or268(N268,N2232,N2245);
or or269(N269,N2258,N2271);
or or270(N270,N2284,N2297);
or or271(N271,N2310,N2323);
or or272(N272,N2336,N2348);
or or273(N273,N2360,N2372);
or or274(N274,N2384,N2396);
or or275(N275,N2408,N2420);
or or276(N276,N2432,N2444);
or or277(N277,N2456,N2468);
or or278(N278,N2480,N2492);
or or279(N279,N2504,N2516);
or or280(N280,N2528,N2540);
or or281(N281,N2552,N2564);
or or282(N282,N2575,N2586);
or or283(N283,N2597,N2608);
or or284(N284,N2619,N2630);
or or285(N285,N2641,N2652);
or or286(N286,N2663,N2674);
or or287(N287,N2685,N2696);
or or288(N288,N2707,N2718);
or or289(N289,N2729,N2740);
or or290(N290,N2751,N2762);
or or291(N291,N2773,N2784);
or or292(N292,N2793,N2802);
or or293(N293,N2818,N2834);
or or294(N294,N2850,N2866);
or or295(N295,N2881,N2896);
or or296(N296,N2911,N2926);
or or297(N297,N2941,N2956);
or or298(N298,N2971,N2985);
or or299(N299,N2999,N3013);
or or300(N300,N3027,N3041);
or or301(N301,N3055,N3069);
or or302(N302,N3083,N3097);
or or303(N303,N3111,N3125);
or or304(N304,N3139,N3153);
or or305(N305,N3167,N3181);
or or306(N306,N3195,N3209);
or or307(N307,N3223,N3237);
or or308(N308,N3251,N3265);
or or309(N309,N3279,N3293);
or or310(N310,N3307,N3321);
or or311(N311,N3335,N3349);
or or312(N312,N3363,N3377);
or or313(N313,N3391,N3405);
or or314(N314,N3419,N3433);
or or315(N315,N3447,N3461);
or or316(N316,N3475,N3488);
or or317(N317,N3501,N3514);
or or318(N318,N3527,N3540);
or or319(N319,N3553,N3566);
or or320(N320,N3579,N3592);
or or321(N321,N3605,N3618);
or or322(N322,N3631,N3644);
or or323(N323,N3657,N3670);
or or324(N324,N3683,N3696);
or or325(N325,N3709,N3722);
or or326(N326,N3735,N3748);
or or327(N327,N3761,N3774);
or or328(N328,N3787,N3800);
or or329(N329,N3813,N3826);
or or330(N330,N3839,N3852);
or or331(N331,N3865,N3878);
or or332(N332,N3891,N3904);
or or333(N333,N3917,N3930);
or or334(N334,N3943,N3956);
or or335(N335,N3969,N3981);
or or336(N336,N3993,N4005);
or or337(N337,N4017,N4029);
or or338(N338,N4041,N4053);
or or339(N339,N4065,N4077);
or or340(N340,N4089,N4101);
or or341(N341,N4113,N4125);
or or342(N342,N4137,N4149);
or or343(N343,N4161,N4173);
or or344(N344,N4185,N4197);
or or345(N345,N4209,N4221);
or or346(N346,N4233,N4245);
or or347(N347,N4257,N4269);
or or348(N348,N4281,N4293);
or or349(N349,N4305,N4317);
or or350(N350,N4329,N4341);
or or351(N351,N4353,N4365);
or or352(N352,N4377,N4389);
or or353(N353,N4401,N4413);
or or354(N354,N4425,N4437);
or or355(N355,N4449,N4461);
or or356(N356,N4473,N4485);
or or357(N357,N4497,N4509);
or or358(N358,N4521,N4533);
or or359(N359,N4545,N4557);
or or360(N360,N4569,N4581);
or or361(N361,N4593,N4604);
or or362(N362,N4615,N4626);
or or363(N363,N4637,N4648);
or or364(N364,N4659,N4670);
or or365(N365,N4681,N4692);
or or366(N366,N4703,N4714);
or or367(N367,N4725,N4736);
or or368(N368,N4747,N4758);
or or369(N369,N4769,N4780);
or or370(N370,N4791,N4802);
or or371(N371,N4813,N4824);
or or372(N372,N4835,N4846);
or or373(N373,N4857,N4868);
or or374(N374,N4879,N4890);
or or375(N375,N4900,N4910);
or or376(N376,N4920,N4930);
or or377(N377,N4940,N4950);
or or378(N378,N4960,N4970);
or or379(N379,N4980,N4990);
or or380(N380,N5000,N5010);
or or381(N381,N5020,N5030);
or or382(N382,N5040,N5050);
or or383(N383,N5060,N5070);
or or384(N384,N5079,N5088);
or or385(N385,N5097,N5106);
or or386(N386,N5115,N5124);
or or387(N387,N5138,N5152);
or or388(N388,N5166,N5179);
or or389(N389,N5192,N5205);
or or390(N390,N5218,N5231);
or or391(N391,N5243,N5255);
or or392(N392,N5267,N5279);
or or393(N393,N5291,N5303);
or or394(N394,N5315,N5327);
or or395(N395,N5338,N5349);
or or396(N396,N5360,N5371);
or or397(N397,N5382,N5393);
or or398(N398,N5404,N5415);
or or399(N399,N5426,N5437);
or or400(N400,N5448,N5459);
or or401(N401,N5470,N5481);
or or402(N402,N5491,N5501);
or or403(N403,N5511,N5521);
or or404(N404,N5531,N5541);
or or405(N405,N5551,N5561);
or or406(N406,N5571,N5581);
or or407(N407,N5591,N5601);
or or408(N408,N5610,N5619);
or or409(N409,N5628,N5637);
or or410(N410,N5646,N5654);
or or411(N5661,N5662,N5663);
or or412(N5662,N5664,N5665);
or or413(N5663,N5666,N5667);
or or414(N5664,N5668,N5669);
or or415(N5665,N5670,N5671);
or or416(N5666,N5672,N5673);
or or417(N5667,N5674,N5675);
or or418(N5668,N5676,N5677);
or or419(N5669,N5678,N5679);
or or420(N5670,N5680,N5681);
or or421(N5671,N5682,N5683);
or or422(N5672,N5684,N5685);
or or423(N5673,N5686,N5687);
or or424(N5674,N5688,N5689);
or or425(N5675,N5690,N5691);
or or426(N5676,N5692,N5693);
or or427(N5677,N5694,N5695);
or or428(N5678,N5696,N5697);
or or429(N5679,N5698,N5699);
or or430(N5680,N5700,N5701);
or or431(N5681,N5702,N5703);
or or432(N5682,N5704,N5705);
or or433(N5683,N5706,N5707);
or or434(N5684,N5708,N5709);
or or435(N5685,N5710,N5711);
or or436(N5686,N5712,N5713);
or or437(N5687,N5714,N5715);
or or438(N5688,N5716,N5717);
or or439(N5689,N5718,N5719);
or or440(N5690,N5720,N5721);
or or441(N5691,N5722,N5723);
or or442(N5692,N5724,N5725);
or or443(N5693,N5726,N5727);
or or444(N5694,N5728,N5729);
or or445(N5695,N5730,N5731);
or or446(N5696,N5732,N5733);
or or447(N5697,N5734,N5735);
or or448(N5698,N5736,N5737);
or or449(N5699,N5738,N5739);
or or450(N5700,N5740,N5741);
or or451(N5701,N5742,N5743);
or or452(N5702,N5744,N5745);
or or453(N5703,N5746,N5747);
or or454(N5704,N5748,N5749);
or or455(N5705,N5750,N5751);
or or456(N5706,N5752,N5753);
or or457(N5707,N5754,N5755);
or or458(N5708,N5756,N5757);
or or459(N5709,N5758,N5759);
or or460(N5710,N5760,N5761);
or or461(N5711,N5762,N5763);
or or462(N5712,N5764,N5765);
or or463(N5713,N5766,N5767);
or or464(N5714,N5768,N5769);
or or465(N5715,N5770,N5771);
or or466(N5716,N5772,N5773);
or or467(N5717,N5774,N5775);
or or468(N5718,N5776,N5777);
or or469(N5719,N5778,N5779);
or or470(N5720,N5780,N5781);
or or471(N5721,N5782,N5783);
or or472(N5722,N5784,N5785);
or or473(N5723,N5786,N5787);
or or474(N5724,N5788,N5789);
or or475(N5725,N5790,N5791);
or or476(N5726,N5792,N5793);
or or477(N5727,N5794,N5795);
or or478(N5728,N5796,N5797);
or or479(N5729,N5798,N5799);
or or480(N5730,N5800,N5801);
or or481(N5731,N5802,N5803);
or or482(N5732,N5804,N5805);
or or483(N5733,N5806,N5807);
or or484(N5734,N5808,N5809);
or or485(N5735,N5810,N5811);
or or486(N5736,N5812,N5813);
or or487(N5737,N5814,N5815);
or or488(N5738,N5816,N5817);
or or489(N5739,N5818,N5819);
or or490(N5740,N5820,N5821);
or or491(N5741,N5822,N5823);
or or492(N5742,N5824,N5825);
or or493(N5743,N5826,N5827);
or or494(N5744,N5828,N5829);
or or495(N5745,N5830,N5831);
or or496(N5746,N5832,N5833);
or or497(N5747,N5834,N5835);
or or498(N5748,N5836,N5837);
or or499(N5749,N5838,N5839);
or or500(N5750,N5840,N5841);
or or501(N5751,N5842,N5843);
or or502(N5752,N5844,N5860);
or or503(N5753,N5875,N5892);
or or504(N5754,N5909,N5926);
or or505(N5755,N5943,N5960);
or or506(N5756,N5977,N5994);
or or507(N5757,N6011,N6028);
or or508(N5758,N6045,N6062);
or or509(N5759,N6078,N6094);
or or510(N5760,N6110,N6126);
or or511(N5761,N6142,N6158);
or or512(N5762,N6174,N6190);
or or513(N5763,N6206,N6222);
or or514(N5764,N6238,N6254);
or or515(N5765,N6270,N6286);
or or516(N5766,N6301,N6316);
or or517(N5767,N6331,N6346);
or or518(N5768,N6361,N6376);
or or519(N5769,N6391,N6406);
or or520(N5770,N6421,N6436);
or or521(N5771,N6451,N6466);
or or522(N5772,N6481,N6496);
or or523(N5773,N6511,N6526);
or or524(N5774,N6541,N6556);
or or525(N5775,N6571,N6586);
or or526(N5776,N6601,N6616);
or or527(N5777,N6631,N6646);
or or528(N5778,N6661,N6676);
or or529(N5779,N6691,N6706);
or or530(N5780,N6721,N6736);
or or531(N5781,N6751,N6766);
or or532(N5782,N6781,N6796);
or or533(N5783,N6811,N6826);
or or534(N5784,N6841,N6856);
or or535(N5785,N6871,N6886);
or or536(N5786,N6901,N6916);
or or537(N5787,N6931,N6946);
or or538(N5788,N6960,N6974);
or or539(N5789,N6988,N7002);
or or540(N5790,N7016,N7030);
or or541(N5791,N7044,N7058);
or or542(N5792,N7072,N7086);
or or543(N5793,N7100,N7114);
or or544(N5794,N7128,N7142);
or or545(N5795,N7156,N7170);
or or546(N5796,N7184,N7198);
or or547(N5797,N7212,N7226);
or or548(N5798,N7240,N7254);
or or549(N5799,N7268,N7281);
or or550(N5800,N7294,N7307);
or or551(N5801,N7320,N7333);
or or552(N5802,N7346,N7359);
or or553(N5803,N7372,N7385);
or or554(N5804,N7398,N7411);
or or555(N5805,N7424,N7437);
or or556(N5806,N7450,N7463);
or or557(N5807,N7476,N7489);
or or558(N5808,N7502,N7515);
or or559(N5809,N7528,N7541);
or or560(N5810,N7554,N7567);
or or561(N5811,N7580,N7593);
or or562(N5812,N7606,N7619);
or or563(N5813,N7632,N7645);
or or564(N5814,N7658,N7671);
or or565(N5815,N7684,N7697);
or or566(N5816,N7710,N7723);
or or567(N5817,N7736,N7749);
or or568(N5818,N7762,N7775);
or or569(N5819,N7788,N7801);
or or570(N5820,N7814,N7826);
or or571(N5821,N7838,N7850);
or or572(N5822,N7862,N7874);
or or573(N5823,N7886,N7898);
or or574(N5824,N7910,N7922);
or or575(N5825,N7934,N7946);
or or576(N5826,N7958,N7970);
or or577(N5827,N7981,N7992);
or or578(N5828,N8003,N8014);
or or579(N5829,N8025,N8036);
or or580(N5830,N8047,N8058);
or or581(N5831,N8068,N8084);
or or582(N5832,N8100,N8116);
or or583(N5833,N8132,N8147);
or or584(N5834,N8162,N8177);
or or585(N5835,N8192,N8206);
or or586(N5836,N8220,N8234);
or or587(N5837,N8248,N8262);
or or588(N5838,N8275,N8288);
or or589(N5839,N8301,N8314);
or or590(N5840,N8327,N8340);
or or591(N5841,N8353,N8365);
or or592(N5842,N8377,N8389);
or or593(N5843,N8401,N8413);
or or594(N8425,N8426,N8427);
or or595(N8426,N8428,N8429);
or or596(N8427,N8430,N8431);
or or597(N8428,N8432,N8433);
or or598(N8429,N8434,N8435);
or or599(N8430,N8436,N8437);
or or600(N8431,N8438,N8439);
or or601(N8432,N8440,N8441);
or or602(N8433,N8442,N8443);
or or603(N8434,N8444,N8445);
or or604(N8435,N8446,N8447);
or or605(N8436,N8448,N8449);
or or606(N8437,N8450,N8451);
or or607(N8438,N8452,N8453);
or or608(N8439,N8454,N8455);
or or609(N8440,N8456,N8457);
or or610(N8441,N8458,N8459);
or or611(N8442,N8460,N8461);
or or612(N8443,N8462,N8463);
or or613(N8444,N8464,N8465);
or or614(N8445,N8466,N8467);
or or615(N8446,N8468,N8469);
or or616(N8447,N8470,N8471);
or or617(N8448,N8472,N8473);
or or618(N8449,N8474,N8475);
or or619(N8450,N8476,N8477);
or or620(N8451,N8478,N8479);
or or621(N8452,N8480,N8481);
or or622(N8453,N8482,N8483);
or or623(N8454,N8484,N8485);
or or624(N8455,N8486,N8487);
or or625(N8456,N8488,N8489);
or or626(N8457,N8490,N8491);
or or627(N8458,N8492,N8493);
or or628(N8459,N8494,N8495);
or or629(N8460,N8496,N8497);
or or630(N8461,N8498,N8499);
or or631(N8462,N8500,N8501);
or or632(N8463,N8502,N8503);
or or633(N8464,N8504,N8505);
or or634(N8465,N8506,N8507);
or or635(N8466,N8508,N8509);
or or636(N8467,N8510,N8511);
or or637(N8468,N8512,N8513);
or or638(N8469,N8514,N8515);
or or639(N8470,N8516,N8517);
or or640(N8471,N8518,N8519);
or or641(N8472,N8520,N8521);
or or642(N8473,N8522,N8523);
or or643(N8474,N8524,N8525);
or or644(N8475,N8526,N8527);
or or645(N8476,N8528,N8529);
or or646(N8477,N8530,N8531);
or or647(N8478,N8532,N8533);
or or648(N8479,N8534,N8535);
or or649(N8480,N8536,N8537);
or or650(N8481,N8538,N8539);
or or651(N8482,N8540,N8541);
or or652(N8483,N8542,N8543);
or or653(N8484,N8544,N8545);
or or654(N8485,N8546,N8547);
or or655(N8486,N8548,N8549);
or or656(N8487,N8550,N8551);
or or657(N8488,N8552,N8553);
or or658(N8489,N8554,N8555);
or or659(N8490,N8556,N8557);
or or660(N8491,N8558,N8559);
or or661(N8492,N8560,N8561);
or or662(N8493,N8562,N8563);
or or663(N8494,N8564,N8565);
or or664(N8495,N8566,N8567);
or or665(N8496,N8568,N8569);
or or666(N8497,N8570,N8571);
or or667(N8498,N8572,N8573);
or or668(N8499,N8574,N8575);
or or669(N8500,N8576,N8577);
or or670(N8501,N8578,N8579);
or or671(N8502,N8580,N8581);
or or672(N8503,N8582,N8583);
or or673(N8504,N8584,N8585);
or or674(N8505,N8586,N8587);
or or675(N8506,N8588,N8589);
or or676(N8507,N8590,N8591);
or or677(N8508,N8592,N8593);
or or678(N8509,N8594,N8595);
or or679(N8510,N8596,N8597);
or or680(N8511,N8598,N8599);
or or681(N8512,N8600,N8601);
or or682(N8513,N8602,N8603);
or or683(N8514,N8604,N8605);
or or684(N8515,N8606,N8607);
or or685(N8516,N8608,N8609);
or or686(N8517,N8610,N8611);
or or687(N8518,N8612,N8613);
or or688(N8519,N8614,N8615);
or or689(N8520,N8616,N8617);
or or690(N8521,N8618,N8619);
or or691(N8522,N8620,N8621);
or or692(N8523,N8622,N8623);
or or693(N8524,N8624,N8625);
or or694(N8525,N8626,N8627);
or or695(N8526,N8628,N8629);
or or696(N8527,N8630,N8631);
or or697(N8528,N8632,N8633);
or or698(N8529,N8634,N8635);
or or699(N8530,N8636,N8637);
or or700(N8531,N8638,N8639);
or or701(N8532,N8640,N8641);
or or702(N8533,N8642,N8643);
or or703(N8534,N8644,N8645);
or or704(N8535,N8646,N8647);
or or705(N8536,N8648,N8649);
or or706(N8537,N8650,N8651);
or or707(N8538,N8652,N8653);
or or708(N8539,N8654,N8655);
or or709(N8540,N8656,N8657);
or or710(N8541,N8658,N8659);
or or711(N8542,N8660,N8661);
or or712(N8543,N8662,N8663);
or or713(N8544,N8664,N8665);
or or714(N8545,N8666,N8667);
or or715(N8546,N8668,N8669);
or or716(N8547,N8670,N8671);
or or717(N8548,N8672,N8673);
or or718(N8549,N8674,N8675);
or or719(N8550,N8676,N8677);
or or720(N8551,N8678,N8679);
or or721(N8552,N8680,N8681);
or or722(N8553,N8682,N8683);
or or723(N8554,N8684,N8685);
or or724(N8555,N8686,N8687);
or or725(N8556,N8688,N8689);
or or726(N8557,N8690,N8691);
or or727(N8558,N8692,N8693);
or or728(N8559,N8694,N8695);
or or729(N8560,N8696,N8697);
or or730(N8561,N8698,N8699);
or or731(N8562,N8700,N8701);
or or732(N8563,N8702,N8703);
or or733(N8564,N8704,N8705);
or or734(N8565,N8706,N8707);
or or735(N8566,N8708,N8709);
or or736(N8567,N8710,N8711);
or or737(N8568,N8712,N8713);
or or738(N8569,N8714,N8715);
or or739(N8570,N8716,N8717);
or or740(N8571,N8718,N8719);
or or741(N8572,N8720,N8721);
or or742(N8573,N8722,N8723);
or or743(N8574,N8724,N8725);
or or744(N8575,N8726,N8727);
or or745(N8576,N8728,N8729);
or or746(N8577,N8730,N8731);
or or747(N8578,N8732,N8733);
or or748(N8579,N8734,N8735);
or or749(N8580,N8736,N8737);
or or750(N8581,N8738,N8739);
or or751(N8582,N8740,N8741);
or or752(N8583,N8742,N8743);
or or753(N8584,N8744,N8745);
or or754(N8585,N8746,N8747);
or or755(N8586,N8748,N8749);
or or756(N8587,N8750,N8751);
or or757(N8588,N8752,N8753);
or or758(N8589,N8754,N8755);
or or759(N8590,N8756,N8757);
or or760(N8591,N8758,N8759);
or or761(N8592,N8760,N8761);
or or762(N8593,N8762,N8763);
or or763(N8594,N8764,N8765);
or or764(N8595,N8766,N8767);
or or765(N8596,N8768,N8769);
or or766(N8597,N8770,N8771);
or or767(N8598,N8772,N8773);
or or768(N8599,N8774,N8775);
or or769(N8600,N8776,N8777);
or or770(N8601,N8778,N8779);
or or771(N8602,N8780,N8781);
or or772(N8603,N8782,N8783);
or or773(N8604,N8784,N8785);
or or774(N8605,N8786,N8787);
or or775(N8606,N8788,N8789);
or or776(N8607,N8790,N8791);
or or777(N8608,N8792,N8793);
or or778(N8609,N8794,N8795);
or or779(N8610,N8796,N8797);
or or780(N8611,N8798,N8799);
or or781(N8612,N8800,N8801);
or or782(N8613,N8802,N8803);
or or783(N8614,N8804,N8805);
or or784(N8615,N8806,N8807);
or or785(N8616,N8808,N8809);
or or786(N8617,N8810,N8811);
or or787(N8618,N8812,N8813);
or or788(N8619,N8814,N8815);
or or789(N8620,N8816,N8817);
or or790(N8621,N8818,N8819);
or or791(N8622,N8820,N8821);
or or792(N8623,N8822,N8823);
or or793(N8624,N8824,N8825);
or or794(N8625,N8826,N8827);
or or795(N8626,N8828,N8829);
or or796(N8627,N8830,N8831);
or or797(N8628,N8832,N8833);
or or798(N8629,N8834,N8835);
or or799(N8630,N8836,N8837);
or or800(N8631,N8838,N8839);
or or801(N8632,N8840,N8841);
or or802(N8633,N8842,N8843);
or or803(N8634,N8844,N8845);
or or804(N8635,N8846,N8847);
or or805(N8636,N8848,N8849);
or or806(N8637,N8850,N8851);
or or807(N8638,N8852,N8853);
or or808(N8639,N8854,N8855);
or or809(N8640,N8856,N8857);
or or810(N8641,N8858,N8859);
or or811(N8642,N8860,N8861);
or or812(N8643,N8862,N8863);
or or813(N8644,N8864,N8865);
or or814(N8645,N8866,N8867);
or or815(N8646,N8868,N8869);
or or816(N8647,N8870,N8871);
or or817(N8648,N8872,N8873);
or or818(N8649,N8874,N8875);
or or819(N8650,N8876,N8877);
or or820(N8651,N8878,N8879);
or or821(N8652,N8880,N8881);
or or822(N8653,N8882,N8883);
or or823(N8654,N8884,N8885);
or or824(N8655,N8903,N8920);
or or825(N8656,N8937,N8954);
or or826(N8657,N8971,N8988);
or or827(N8658,N9004,N9020);
or or828(N8659,N9036,N9052);
or or829(N8660,N9068,N9084);
or or830(N8661,N9100,N9116);
or or831(N8662,N9132,N9148);
or or832(N8663,N9164,N9180);
or or833(N8664,N9196,N9212);
or or834(N8665,N9228,N9243);
or or835(N8666,N9258,N9273);
or or836(N8667,N9288,N9303);
or or837(N8668,N9318,N9333);
or or838(N8669,N9348,N9363);
or or839(N8670,N9378,N9393);
or or840(N8671,N9408,N9423);
or or841(N8672,N9438,N9453);
or or842(N8673,N9468,N9483);
or or843(N8674,N9498,N9513);
or or844(N8675,N9528,N9543);
or or845(N8676,N9558,N9573);
or or846(N8677,N9588,N9603);
or or847(N8678,N9618,N9633);
or or848(N8679,N9648,N9663);
or or849(N8680,N9678,N9693);
or or850(N8681,N9708,N9723);
or or851(N8682,N9738,N9752);
or or852(N8683,N9766,N9780);
or or853(N8684,N9794,N9808);
or or854(N8685,N9822,N9836);
or or855(N8686,N9850,N9864);
or or856(N8687,N9878,N9892);
or or857(N8688,N9906,N9920);
or or858(N8689,N9934,N9948);
or or859(N8690,N9962,N9976);
or or860(N8691,N9990,N10004);
or or861(N8692,N10018,N10032);
or or862(N8693,N10046,N10060);
or or863(N8694,N10074,N10088);
or or864(N8695,N10102,N10116);
or or865(N8696,N10130,N10144);
or or866(N8697,N10158,N10172);
or or867(N8698,N10186,N10200);
or or868(N8699,N10214,N10228);
or or869(N8700,N10242,N10256);
or or870(N8701,N10270,N10284);
or or871(N8702,N10298,N10311);
or or872(N8703,N10324,N10337);
or or873(N8704,N10350,N10363);
or or874(N8705,N10376,N10389);
or or875(N8706,N10402,N10415);
or or876(N8707,N10428,N10441);
or or877(N8708,N10454,N10467);
or or878(N8709,N10480,N10493);
or or879(N8710,N10506,N10519);
or or880(N8711,N10532,N10545);
or or881(N8712,N10558,N10571);
or or882(N8713,N10584,N10597);
or or883(N8714,N10610,N10623);
or or884(N8715,N10636,N10649);
or or885(N8716,N10662,N10675);
or or886(N8717,N10688,N10701);
or or887(N8718,N10714,N10727);
or or888(N8719,N10740,N10753);
or or889(N8720,N10766,N10779);
or or890(N8721,N10792,N10805);
or or891(N8722,N10818,N10830);
or or892(N8723,N10842,N10854);
or or893(N8724,N10866,N10878);
or or894(N8725,N10890,N10902);
or or895(N8726,N10914,N10926);
or or896(N8727,N10938,N10950);
or or897(N8728,N10962,N10974);
or or898(N8729,N10986,N10998);
or or899(N8730,N11010,N11022);
or or900(N8731,N11034,N11046);
or or901(N8732,N11058,N11070);
or or902(N8733,N11082,N11094);
or or903(N8734,N11106,N11118);
or or904(N8735,N11130,N11142);
or or905(N8736,N11153,N11164);
or or906(N8737,N11175,N11186);
or or907(N8738,N11197,N11208);
or or908(N8739,N11219,N11230);
or or909(N8740,N11241,N11252);
or or910(N8741,N11263,N11274);
or or911(N8742,N11285,N11296);
or or912(N8743,N11307,N11318);
or or913(N8744,N11328,N11338);
or or914(N8745,N11348,N11358);
or or915(N8746,N11368,N11384);
or or916(N8747,N11400,N11416);
or or917(N8748,N11432,N11448);
or or918(N8749,N11464,N11480);
or or919(N8750,N11495,N11510);
or or920(N8751,N11525,N11540);
or or921(N8752,N11555,N11570);
or or922(N8753,N11585,N11599);
or or923(N8754,N11613,N11627);
or or924(N8755,N11641,N11655);
or or925(N8756,N11669,N11683);
or or926(N8757,N11697,N11711);
or or927(N8758,N11725,N11739);
or or928(N8759,N11753,N11767);
or or929(N8760,N11781,N11795);
or or930(N8761,N11809,N11823);
or or931(N8762,N11837,N11851);
or or932(N8763,N11865,N11879);
or or933(N8764,N11893,N11907);
or or934(N8765,N11921,N11935);
or or935(N8766,N11949,N11963);
or or936(N8767,N11977,N11991);
or or937(N8768,N12005,N12019);
or or938(N8769,N12033,N12047);
or or939(N8770,N12061,N12075);
or or940(N8771,N12088,N12101);
or or941(N8772,N12114,N12127);
or or942(N8773,N12140,N12153);
or or943(N8774,N12166,N12179);
or or944(N8775,N12192,N12205);
or or945(N8776,N12218,N12231);
or or946(N8777,N12244,N12257);
or or947(N8778,N12270,N12283);
or or948(N8779,N12296,N12309);
or or949(N8780,N12322,N12335);
or or950(N8781,N12348,N12361);
or or951(N8782,N12374,N12387);
or or952(N8783,N12400,N12413);
or or953(N8784,N12426,N12439);
or or954(N8785,N12452,N12465);
or or955(N8786,N12478,N12491);
or or956(N8787,N12504,N12517);
or or957(N8788,N12530,N12543);
or or958(N8789,N12556,N12569);
or or959(N8790,N12582,N12595);
or or960(N8791,N12608,N12621);
or or961(N8792,N12634,N12647);
or or962(N8793,N12660,N12673);
or or963(N8794,N12685,N12697);
or or964(N8795,N12709,N12721);
or or965(N8796,N12733,N12745);
or or966(N8797,N12757,N12769);
or or967(N8798,N12781,N12793);
or or968(N8799,N12805,N12817);
or or969(N8800,N12829,N12841);
or or970(N8801,N12853,N12865);
or or971(N8802,N12877,N12889);
or or972(N8803,N12901,N12913);
or or973(N8804,N12925,N12937);
or or974(N8805,N12949,N12961);
or or975(N8806,N12973,N12985);
or or976(N8807,N12997,N13009);
or or977(N8808,N13021,N13033);
or or978(N8809,N13045,N13057);
or or979(N8810,N13069,N13081);
or or980(N8811,N13093,N13105);
or or981(N8812,N13117,N13129);
or or982(N8813,N13141,N13153);
or or983(N8814,N13165,N13177);
or or984(N8815,N13189,N13201);
or or985(N8816,N13213,N13225);
or or986(N8817,N13237,N13249);
or or987(N8818,N13261,N13273);
or or988(N8819,N13285,N13297);
or or989(N8820,N13309,N13321);
or or990(N8821,N13333,N13345);
or or991(N8822,N13357,N13369);
or or992(N8823,N13381,N13393);
or or993(N8824,N13404,N13415);
or or994(N8825,N13426,N13437);
or or995(N8826,N13448,N13459);
or or996(N8827,N13470,N13481);
or or997(N8828,N13492,N13503);
or or998(N8829,N13514,N13525);
or or999(N8830,N13536,N13547);
or or1000(N8831,N13558,N13569);
or or1001(N8832,N13580,N13591);
or or1002(N8833,N13602,N13613);
or or1003(N8834,N13624,N13635);
or or1004(N8835,N13646,N13657);
or or1005(N8836,N13668,N13679);
or or1006(N8837,N13690,N13701);
or or1007(N8838,N13712,N13723);
or or1008(N8839,N13734,N13745);
or or1009(N8840,N13756,N13767);
or or1010(N8841,N13778,N13789);
or or1011(N8842,N13800,N13811);
or or1012(N8843,N13822,N13833);
or or1013(N8844,N13844,N13855);
or or1014(N8845,N13866,N13877);
or or1015(N8846,N13888,N13899);
or or1016(N8847,N13910,N13921);
or or1017(N8848,N13932,N13943);
or or1018(N8849,N13954,N13964);
or or1019(N8850,N13974,N13984);
or or1020(N8851,N13994,N14004);
or or1021(N8852,N14014,N14024);
or or1022(N8853,N14034,N14044);
or or1023(N8854,N14054,N14064);
or or1024(N8855,N14074,N14084);
or or1025(N8856,N14094,N14104);
or or1026(N8857,N14114,N14123);
or or1027(N8858,N14132,N14141);
or or1028(N8859,N14150,N14159);
or or1029(N8860,N14168,N14177);
or or1030(N8861,N14186,N14195);
or or1031(N8862,N14204,N14218);
or or1032(N8863,N14232,N14246);
or or1033(N8864,N14260,N14273);
or or1034(N8865,N14286,N14299);
or or1035(N8866,N14312,N14325);
or or1036(N8867,N14338,N14351);
or or1037(N8868,N14363,N14375);
or or1038(N8869,N14387,N14399);
or or1039(N8870,N14411,N14423);
or or1040(N8871,N14435,N14447);
or or1041(N8872,N14459,N14471);
or or1042(N8873,N14483,N14495);
or or1043(N8874,N14507,N14518);
or or1044(N8875,N14529,N14540);
or or1045(N8876,N14551,N14562);
or or1046(N8877,N14573,N14584);
or or1047(N8878,N14595,N14606);
or or1048(N8879,N14616,N14626);
or or1049(N8880,N14636,N14646);
or or1050(N8881,N14656,N14665);
or or1051(N8882,N14674,N14683);
or or1052(N8883,N14692,N14701);
or or1053(N8884,N14708,N14718);
or or1054(N14726,N14727,N14728);
or or1055(N14727,N14729,N14730);
or or1056(N14728,N14731,N14732);
or or1057(N14729,N14733,N14734);
or or1058(N14730,N14735,N14736);
or or1059(N14731,N14737,N14738);
or or1060(N14732,N14739,N14740);
or or1061(N14733,N14741,N14742);
or or1062(N14734,N14743,N14744);
or or1063(N14735,N14745,N14746);
or or1064(N14736,N14747,N14748);
or or1065(N14737,N14749,N14750);
or or1066(N14738,N14751,N14752);
or or1067(N14739,N14753,N14754);
or or1068(N14740,N14755,N14756);
or or1069(N14741,N14757,N14758);
or or1070(N14742,N14759,N14760);
or or1071(N14743,N14761,N14762);
or or1072(N14744,N14763,N14764);
or or1073(N14745,N14765,N14766);
or or1074(N14746,N14767,N14768);
or or1075(N14747,N14769,N14770);
or or1076(N14748,N14771,N14772);
or or1077(N14749,N14773,N14774);
or or1078(N14750,N14775,N14776);
or or1079(N14751,N14777,N14778);
or or1080(N14752,N14779,N14780);
or or1081(N14753,N14781,N14782);
or or1082(N14754,N14783,N14784);
or or1083(N14755,N14785,N14786);
or or1084(N14756,N14787,N14788);
or or1085(N14757,N14789,N14790);
or or1086(N14758,N14791,N14792);
or or1087(N14759,N14793,N14794);
or or1088(N14760,N14795,N14796);
or or1089(N14761,N14797,N14798);
or or1090(N14762,N14799,N14800);
or or1091(N14763,N14801,N14802);
or or1092(N14764,N14803,N14804);
or or1093(N14765,N14805,N14806);
or or1094(N14766,N14807,N14808);
or or1095(N14767,N14809,N14810);
or or1096(N14768,N14811,N14812);
or or1097(N14769,N14813,N14814);
or or1098(N14770,N14815,N14816);
or or1099(N14771,N14817,N14818);
or or1100(N14772,N14819,N14820);
or or1101(N14773,N14821,N14822);
or or1102(N14774,N14823,N14824);
or or1103(N14775,N14825,N14826);
or or1104(N14776,N14827,N14828);
or or1105(N14777,N14829,N14830);
or or1106(N14778,N14831,N14832);
or or1107(N14779,N14833,N14834);
or or1108(N14780,N14835,N14836);
or or1109(N14781,N14837,N14838);
or or1110(N14782,N14839,N14840);
or or1111(N14783,N14841,N14842);
or or1112(N14784,N14843,N14844);
or or1113(N14785,N14845,N14846);
or or1114(N14786,N14847,N14848);
or or1115(N14787,N14849,N14850);
or or1116(N14788,N14851,N14852);
or or1117(N14789,N14853,N14854);
or or1118(N14790,N14855,N14856);
or or1119(N14791,N14857,N14858);
or or1120(N14792,N14859,N14860);
or or1121(N14793,N14861,N14862);
or or1122(N14794,N14863,N14864);
or or1123(N14795,N14865,N14866);
or or1124(N14796,N14867,N14868);
or or1125(N14797,N14869,N14870);
or or1126(N14798,N14871,N14872);
or or1127(N14799,N14873,N14874);
or or1128(N14800,N14875,N14876);
or or1129(N14801,N14877,N14878);
or or1130(N14802,N14879,N14880);
or or1131(N14803,N14881,N14882);
or or1132(N14804,N14883,N14884);
or or1133(N14805,N14885,N14886);
or or1134(N14806,N14887,N14888);
or or1135(N14807,N14889,N14890);
or or1136(N14808,N14891,N14892);
or or1137(N14809,N14893,N14894);
or or1138(N14810,N14895,N14896);
or or1139(N14811,N14897,N14898);
or or1140(N14812,N14899,N14900);
or or1141(N14813,N14901,N14902);
or or1142(N14814,N14903,N14904);
or or1143(N14815,N14905,N14906);
or or1144(N14816,N14907,N14908);
or or1145(N14817,N14909,N14910);
or or1146(N14818,N14911,N14912);
or or1147(N14819,N14913,N14914);
or or1148(N14820,N14915,N14916);
or or1149(N14821,N14917,N14918);
or or1150(N14822,N14919,N14920);
or or1151(N14823,N14921,N14922);
or or1152(N14824,N14923,N14924);
or or1153(N14825,N14925,N14926);
or or1154(N14826,N14927,N14928);
or or1155(N14827,N14929,N14930);
or or1156(N14828,N14931,N14932);
or or1157(N14829,N14933,N14934);
or or1158(N14830,N14935,N14936);
or or1159(N14831,N14937,N14938);
or or1160(N14832,N14939,N14940);
or or1161(N14833,N14941,N14942);
or or1162(N14834,N14943,N14944);
or or1163(N14835,N14945,N14946);
or or1164(N14836,N14947,N14948);
or or1165(N14837,N14949,N14950);
or or1166(N14838,N14951,N14952);
or or1167(N14839,N14953,N14954);
or or1168(N14840,N14955,N14956);
or or1169(N14841,N14957,N14958);
or or1170(N14842,N14959,N14960);
or or1171(N14843,N14961,N14962);
or or1172(N14844,N14963,N14964);
or or1173(N14845,N14965,N14966);
or or1174(N14846,N14967,N14968);
or or1175(N14847,N14969,N14970);
or or1176(N14848,N14971,N14972);
or or1177(N14849,N14973,N14974);
or or1178(N14850,N14975,N14976);
or or1179(N14851,N14977,N14978);
or or1180(N14852,N14979,N14980);
or or1181(N14853,N14981,N14982);
or or1182(N14854,N14983,N14984);
or or1183(N14855,N14985,N14986);
or or1184(N14856,N14987,N14988);
or or1185(N14857,N14989,N14990);
or or1186(N14858,N14991,N14992);
or or1187(N14859,N14993,N14994);
or or1188(N14860,N14995,N14996);
or or1189(N14861,N14997,N14998);
or or1190(N14862,N14999,N15000);
or or1191(N14863,N15001,N15002);
or or1192(N14864,N15003,N15004);
or or1193(N14865,N15005,N15006);
or or1194(N14866,N15007,N15008);
or or1195(N14867,N15009,N15010);
or or1196(N14868,N15011,N15012);
or or1197(N14869,N15013,N15014);
or or1198(N14870,N15015,N15016);
or or1199(N14871,N15017,N15018);
or or1200(N14872,N15019,N15020);
or or1201(N14873,N15021,N15022);
or or1202(N14874,N15023,N15024);
or or1203(N14875,N15025,N15026);
or or1204(N14876,N15027,N15028);
or or1205(N14877,N15029,N15030);
or or1206(N14878,N15031,N15032);
or or1207(N14879,N15033,N15034);
or or1208(N14880,N15035,N15036);
or or1209(N14881,N15037,N15038);
or or1210(N14882,N15039,N15040);
or or1211(N14883,N15041,N15042);
or or1212(N14884,N15043,N15044);
or or1213(N14885,N15045,N15046);
or or1214(N14886,N15047,N15048);
or or1215(N14887,N15049,N15050);
or or1216(N14888,N15051,N15052);
or or1217(N14889,N15053,N15054);
or or1218(N14890,N15055,N15056);
or or1219(N14891,N15057,N15058);
or or1220(N14892,N15059,N15060);
or or1221(N14893,N15061,N15062);
or or1222(N14894,N15063,N15064);
or or1223(N14895,N15065,N15066);
or or1224(N14896,N15067,N15068);
or or1225(N14897,N15069,N15070);
or or1226(N14898,N15071,N15072);
or or1227(N14899,N15073,N15074);
or or1228(N14900,N15075,N15076);
or or1229(N14901,N15077,N15078);
or or1230(N14902,N15079,N15080);
or or1231(N14903,N15081,N15082);
or or1232(N14904,N15083,N15084);
or or1233(N14905,N15085,N15086);
or or1234(N14906,N15087,N15088);
or or1235(N14907,N15089,N15090);
or or1236(N14908,N15091,N15092);
or or1237(N14909,N15093,N15094);
or or1238(N14910,N15095,N15096);
or or1239(N14911,N15097,N15098);
or or1240(N14912,N15099,N15100);
or or1241(N14913,N15101,N15102);
or or1242(N14914,N15103,N15104);
or or1243(N14915,N15105,N15106);
or or1244(N14916,N15107,N15108);
or or1245(N14917,N15109,N15110);
or or1246(N14918,N15111,N15112);
or or1247(N14919,N15113,N15114);
or or1248(N14920,N15115,N15116);
or or1249(N14921,N15117,N15118);
or or1250(N14922,N15119,N15120);
or or1251(N14923,N15121,N15122);
or or1252(N14924,N15123,N15124);
or or1253(N14925,N15125,N15126);
or or1254(N14926,N15127,N15128);
or or1255(N14927,N15129,N15130);
or or1256(N14928,N15131,N15132);
or or1257(N14929,N15133,N15134);
or or1258(N14930,N15135,N15136);
or or1259(N14931,N15137,N15138);
or or1260(N14932,N15139,N15140);
or or1261(N14933,N15141,N15142);
or or1262(N14934,N15143,N15144);
or or1263(N14935,N15145,N15146);
or or1264(N14936,N15164,N15181);
or or1265(N14937,N15198,N15214);
or or1266(N14938,N15230,N15246);
or or1267(N14939,N15262,N15278);
or or1268(N14940,N15294,N15310);
or or1269(N14941,N15326,N15342);
or or1270(N14942,N15357,N15372);
or or1271(N14943,N15387,N15402);
or or1272(N14944,N15417,N15432);
or or1273(N14945,N15447,N15462);
or or1274(N14946,N15477,N15492);
or or1275(N14947,N15507,N15522);
or or1276(N14948,N15537,N15552);
or or1277(N14949,N15566,N15580);
or or1278(N14950,N15594,N15608);
or or1279(N14951,N15622,N15636);
or or1280(N14952,N15650,N15664);
or or1281(N14953,N15678,N15692);
or or1282(N14954,N15706,N15720);
or or1283(N14955,N15734,N15748);
or or1284(N14956,N15762,N15776);
or or1285(N14957,N15790,N15804);
or or1286(N14958,N15818,N15832);
or or1287(N14959,N15846,N15860);
or or1288(N14960,N15874,N15888);
or or1289(N14961,N15902,N15916);
or or1290(N14962,N15930,N15944);
or or1291(N14963,N15958,N15972);
or or1292(N14964,N15986,N16000);
or or1293(N14965,N16014,N16028);
or or1294(N14966,N16042,N16056);
or or1295(N14967,N16070,N16084);
or or1296(N14968,N16098,N16111);
or or1297(N14969,N16124,N16137);
or or1298(N14970,N16150,N16163);
or or1299(N14971,N16176,N16189);
or or1300(N14972,N16202,N16215);
or or1301(N14973,N16228,N16241);
or or1302(N14974,N16254,N16267);
or or1303(N14975,N16280,N16293);
or or1304(N14976,N16306,N16319);
or or1305(N14977,N16332,N16345);
or or1306(N14978,N16358,N16371);
or or1307(N14979,N16384,N16397);
or or1308(N14980,N16410,N16422);
or or1309(N14981,N16434,N16446);
or or1310(N14982,N16458,N16470);
or or1311(N14983,N16482,N16494);
or or1312(N14984,N16506,N16518);
or or1313(N14985,N16530,N16542);
or or1314(N14986,N16554,N16566);
or or1315(N14987,N16578,N16590);
or or1316(N14988,N16602,N16614);
or or1317(N14989,N16626,N16638);
or or1318(N14990,N16650,N16662);
or or1319(N14991,N16674,N16686);
or or1320(N14992,N16698,N16710);
or or1321(N14993,N16722,N16734);
or or1322(N14994,N16746,N16758);
or or1323(N14995,N16770,N16782);
or or1324(N14996,N16794,N16806);
or or1325(N14997,N16818,N16830);
or or1326(N14998,N16842,N16854);
or or1327(N14999,N16866,N16878);
or or1328(N15000,N16890,N16901);
or or1329(N15001,N16912,N16923);
or or1330(N15002,N16934,N16945);
or or1331(N15003,N16955,N16965);
or or1332(N15004,N16975,N16985);
or or1333(N15005,N16995,N17005);
or or1334(N15006,N17015,N17025);
or or1335(N15007,N17041,N17057);
or or1336(N15008,N17072,N17087);
or or1337(N15009,N17102,N17117);
or or1338(N15010,N17132,N17147);
or or1339(N15011,N17162,N17177);
or or1340(N15012,N17192,N17207);
or or1341(N15013,N17222,N17237);
or or1342(N15014,N17252,N17267);
or or1343(N15015,N17282,N17297);
or or1344(N15016,N17311,N17325);
or or1345(N15017,N17339,N17353);
or or1346(N15018,N17367,N17381);
or or1347(N15019,N17395,N17409);
or or1348(N15020,N17423,N17437);
or or1349(N15021,N17451,N17465);
or or1350(N15022,N17479,N17493);
or or1351(N15023,N17507,N17521);
or or1352(N15024,N17535,N17549);
or or1353(N15025,N17563,N17577);
or or1354(N15026,N17591,N17605);
or or1355(N15027,N17619,N17633);
or or1356(N15028,N17647,N17661);
or or1357(N15029,N17675,N17689);
or or1358(N15030,N17703,N17717);
or or1359(N15031,N17731,N17745);
or or1360(N15032,N17759,N17772);
or or1361(N15033,N17785,N17798);
or or1362(N15034,N17811,N17824);
or or1363(N15035,N17837,N17850);
or or1364(N15036,N17863,N17876);
or or1365(N15037,N17889,N17902);
or or1366(N15038,N17915,N17928);
or or1367(N15039,N17941,N17954);
or or1368(N15040,N17967,N17980);
or or1369(N15041,N17993,N18006);
or or1370(N15042,N18019,N18032);
or or1371(N15043,N18045,N18058);
or or1372(N15044,N18071,N18084);
or or1373(N15045,N18097,N18110);
or or1374(N15046,N18123,N18136);
or or1375(N15047,N18149,N18162);
or or1376(N15048,N18175,N18188);
or or1377(N15049,N18201,N18214);
or or1378(N15050,N18227,N18240);
or or1379(N15051,N18253,N18266);
or or1380(N15052,N18279,N18292);
or or1381(N15053,N18305,N18318);
or or1382(N15054,N18331,N18344);
or or1383(N15055,N18357,N18370);
or or1384(N15056,N18383,N18396);
or or1385(N15057,N18409,N18422);
or or1386(N15058,N18435,N18448);
or or1387(N15059,N18461,N18474);
or or1388(N15060,N18487,N18500);
or or1389(N15061,N18513,N18526);
or or1390(N15062,N18539,N18552);
or or1391(N15063,N18565,N18578);
or or1392(N15064,N18591,N18603);
or or1393(N15065,N18615,N18627);
or or1394(N15066,N18639,N18651);
or or1395(N15067,N18663,N18675);
or or1396(N15068,N18687,N18699);
or or1397(N15069,N18711,N18723);
or or1398(N15070,N18735,N18747);
or or1399(N15071,N18759,N18771);
or or1400(N15072,N18783,N18795);
or or1401(N15073,N18807,N18819);
or or1402(N15074,N18831,N18843);
or or1403(N15075,N18855,N18867);
or or1404(N15076,N18879,N18891);
or or1405(N15077,N18903,N18915);
or or1406(N15078,N18927,N18939);
or or1407(N15079,N18951,N18963);
or or1408(N15080,N18975,N18987);
or or1409(N15081,N18999,N19011);
or or1410(N15082,N19023,N19035);
or or1411(N15083,N19047,N19059);
or or1412(N15084,N19071,N19083);
or or1413(N15085,N19095,N19107);
or or1414(N15086,N19119,N19131);
or or1415(N15087,N19143,N19155);
or or1416(N15088,N19166,N19177);
or or1417(N15089,N19188,N19199);
or or1418(N15090,N19210,N19221);
or or1419(N15091,N19232,N19243);
or or1420(N15092,N19254,N19265);
or or1421(N15093,N19276,N19287);
or or1422(N15094,N19298,N19309);
or or1423(N15095,N19320,N19331);
or or1424(N15096,N19342,N19353);
or or1425(N15097,N19364,N19375);
or or1426(N15098,N19386,N19397);
or or1427(N15099,N19408,N19419);
or or1428(N15100,N19430,N19441);
or or1429(N15101,N19452,N19463);
or or1430(N15102,N19474,N19485);
or or1431(N15103,N19496,N19507);
or or1432(N15104,N19518,N19529);
or or1433(N15105,N19540,N19551);
or or1434(N15106,N19562,N19573);
or or1435(N15107,N19583,N19593);
or or1436(N15108,N19603,N19613);
or or1437(N15109,N19623,N19633);
or or1438(N15110,N19643,N19653);
or or1439(N15111,N19663,N19673);
or or1440(N15112,N19683,N19693);
or or1441(N15113,N19703,N19713);
or or1442(N15114,N19723,N19733);
or or1443(N15115,N19743,N19753);
or or1444(N15116,N19763,N19772);
or or1445(N15117,N19781,N19790);
or or1446(N15118,N19799,N19808);
or or1447(N15119,N19817,N19826);
or or1448(N15120,N19835,N19844);
or or1449(N15121,N19852,N19866);
or or1450(N15122,N19880,N19894);
or or1451(N15123,N19908,N19922);
or or1452(N15124,N19935,N19948);
or or1453(N15125,N19961,N19973);
or or1454(N15126,N19985,N19997);
or or1455(N15127,N20009,N20021);
or or1456(N15128,N20033,N20045);
or or1457(N15129,N20057,N20069);
or or1458(N15130,N20081,N20092);
or or1459(N15131,N20103,N20114);
or or1460(N15132,N20125,N20136);
or or1461(N15133,N20147,N20158);
or or1462(N15134,N20169,N20180);
or or1463(N15135,N20191,N20202);
or or1464(N15136,N20213,N20224);
or or1465(N15137,N20234,N20244);
or or1466(N15138,N20254,N20264);
or or1467(N15139,N20274,N20284);
or or1468(N15140,N20294,N20304);
or or1469(N15141,N20314,N20324);
or or1470(N15142,N20334,N20343);
or or1471(N15143,N20352,N20361);
or or1472(N15144,N20370,N20378);
or or1473(N15145,N20386,N20394);
or or1474(N20402,N20403,N20404);
or or1475(N20403,N20405,N20406);
or or1476(N20404,N20407,N20408);
or or1477(N20405,N20409,N20410);
or or1478(N20406,N20411,N20412);
or or1479(N20407,N20413,N20414);
or or1480(N20408,N20415,N20416);
or or1481(N20409,N20417,N20418);
or or1482(N20410,N20419,N20420);
or or1483(N20411,N20421,N20422);
or or1484(N20412,N20423,N20424);
or or1485(N20413,N20425,N20426);
or or1486(N20414,N20427,N20428);
or or1487(N20415,N20429,N20430);
or or1488(N20416,N20431,N20432);
or or1489(N20417,N20433,N20434);
or or1490(N20418,N20435,N20436);
or or1491(N20419,N20437,N20438);
or or1492(N20420,N20439,N20440);
or or1493(N20421,N20441,N20442);
or or1494(N20422,N20443,N20444);
or or1495(N20423,N20445,N20446);
or or1496(N20424,N20447,N20448);
or or1497(N20425,N20449,N20450);
or or1498(N20426,N20451,N20452);
or or1499(N20427,N20453,N20454);
or or1500(N20428,N20455,N20456);
or or1501(N20429,N20457,N20458);
or or1502(N20430,N20459,N20460);
or or1503(N20431,N20461,N20462);
or or1504(N20432,N20463,N20464);
or or1505(N20433,N20465,N20466);
or or1506(N20434,N20467,N20468);
or or1507(N20435,N20469,N20470);
or or1508(N20436,N20471,N20472);
or or1509(N20437,N20473,N20474);
or or1510(N20438,N20475,N20476);
or or1511(N20439,N20477,N20478);
or or1512(N20440,N20479,N20480);
or or1513(N20441,N20481,N20482);
or or1514(N20442,N20483,N20484);
or or1515(N20443,N20485,N20486);
or or1516(N20444,N20487,N20488);
or or1517(N20445,N20489,N20490);
or or1518(N20446,N20491,N20492);
or or1519(N20447,N20493,N20494);
or or1520(N20448,N20495,N20496);
or or1521(N20449,N20497,N20498);
or or1522(N20450,N20499,N20500);
or or1523(N20451,N20501,N20502);
or or1524(N20452,N20503,N20504);
or or1525(N20453,N20505,N20506);
or or1526(N20454,N20507,N20508);
or or1527(N20455,N20509,N20510);
or or1528(N20456,N20511,N20512);
or or1529(N20457,N20513,N20514);
or or1530(N20458,N20515,N20516);
or or1531(N20459,N20517,N20518);
or or1532(N20460,N20519,N20520);
or or1533(N20461,N20521,N20522);
or or1534(N20462,N20523,N20524);
or or1535(N20463,N20525,N20526);
or or1536(N20464,N20527,N20528);
or or1537(N20465,N20529,N20530);
or or1538(N20466,N20531,N20532);
or or1539(N20467,N20533,N20534);
or or1540(N20468,N20535,N20536);
or or1541(N20469,N20537,N20538);
or or1542(N20470,N20539,N20540);
or or1543(N20471,N20541,N20542);
or or1544(N20472,N20543,N20544);
or or1545(N20473,N20545,N20546);
or or1546(N20474,N20547,N20548);
or or1547(N20475,N20549,N20550);
or or1548(N20476,N20551,N20552);
or or1549(N20477,N20553,N20554);
or or1550(N20478,N20555,N20556);
or or1551(N20479,N20557,N20558);
or or1552(N20480,N20559,N20560);
or or1553(N20481,N20561,N20562);
or or1554(N20482,N20563,N20564);
or or1555(N20483,N20565,N20566);
or or1556(N20484,N20567,N20568);
or or1557(N20485,N20569,N20570);
or or1558(N20486,N20571,N20572);
or or1559(N20487,N20573,N20574);
or or1560(N20488,N20575,N20576);
or or1561(N20489,N20577,N20578);
or or1562(N20490,N20579,N20580);
or or1563(N20491,N20581,N20582);
or or1564(N20492,N20583,N20584);
or or1565(N20493,N20585,N20586);
or or1566(N20494,N20587,N20588);
or or1567(N20495,N20589,N20590);
or or1568(N20496,N20591,N20592);
or or1569(N20497,N20593,N20594);
or or1570(N20498,N20595,N20596);
or or1571(N20499,N20597,N20598);
or or1572(N20500,N20599,N20600);
or or1573(N20501,N20601,N20602);
or or1574(N20502,N20603,N20604);
or or1575(N20503,N20605,N20606);
or or1576(N20504,N20607,N20608);
or or1577(N20505,N20609,N20610);
or or1578(N20506,N20611,N20612);
or or1579(N20507,N20613,N20614);
or or1580(N20508,N20615,N20616);
or or1581(N20509,N20617,N20618);
or or1582(N20510,N20619,N20620);
or or1583(N20511,N20621,N20622);
or or1584(N20512,N20623,N20624);
or or1585(N20513,N20625,N20626);
or or1586(N20514,N20627,N20628);
or or1587(N20515,N20629,N20630);
or or1588(N20516,N20631,N20632);
or or1589(N20517,N20633,N20634);
or or1590(N20518,N20635,N20651);
or or1591(N20519,N20669,N20687);
or or1592(N20520,N20704,N20721);
or or1593(N20521,N20738,N20755);
or or1594(N20522,N20772,N20789);
or or1595(N20523,N20806,N20823);
or or1596(N20524,N20840,N20857);
or or1597(N20525,N20874,N20891);
or or1598(N20526,N20908,N20924);
or or1599(N20527,N20940,N20956);
or or1600(N20528,N20972,N20988);
or or1601(N20529,N21004,N21020);
or or1602(N20530,N21036,N21052);
or or1603(N20531,N21068,N21084);
or or1604(N20532,N21100,N21116);
or or1605(N20533,N21132,N21148);
or or1606(N20534,N21164,N21180);
or or1607(N20535,N21196,N21212);
or or1608(N20536,N21228,N21244);
or or1609(N20537,N21260,N21276);
or or1610(N20538,N21292,N21308);
or or1611(N20539,N21323,N21338);
or or1612(N20540,N21353,N21368);
or or1613(N20541,N21383,N21398);
or or1614(N20542,N21413,N21428);
or or1615(N20543,N21443,N21458);
or or1616(N20544,N21473,N21488);
or or1617(N20545,N21503,N21518);
or or1618(N20546,N21533,N21548);
or or1619(N20547,N21563,N21578);
or or1620(N20548,N21593,N21608);
or or1621(N20549,N21623,N21638);
or or1622(N20550,N21653,N21668);
or or1623(N20551,N21683,N21697);
or or1624(N20552,N21711,N21725);
or or1625(N20553,N21739,N21753);
or or1626(N20554,N21767,N21781);
or or1627(N20555,N21795,N21809);
or or1628(N20556,N21823,N21837);
or or1629(N20557,N21851,N21865);
or or1630(N20558,N21879,N21893);
or or1631(N20559,N21907,N21921);
or or1632(N20560,N21935,N21949);
or or1633(N20561,N21963,N21977);
or or1634(N20562,N21991,N22005);
or or1635(N20563,N22019,N22033);
or or1636(N20564,N22047,N22061);
or or1637(N20565,N22075,N22089);
or or1638(N20566,N22103,N22117);
or or1639(N20567,N22131,N22145);
or or1640(N20568,N22159,N22173);
or or1641(N20569,N22187,N22201);
or or1642(N20570,N22214,N22227);
or or1643(N20571,N22240,N22253);
or or1644(N20572,N22266,N22279);
or or1645(N20573,N22292,N22305);
or or1646(N20574,N22318,N22331);
or or1647(N20575,N22344,N22357);
or or1648(N20576,N22370,N22383);
or or1649(N20577,N22396,N22409);
or or1650(N20578,N22422,N22435);
or or1651(N20579,N22448,N22461);
or or1652(N20580,N22474,N22487);
or or1653(N20581,N22500,N22513);
or or1654(N20582,N22526,N22539);
or or1655(N20583,N22552,N22565);
or or1656(N20584,N22578,N22591);
or or1657(N20585,N22604,N22617);
or or1658(N20586,N22630,N22643);
or or1659(N20587,N22656,N22669);
or or1660(N20588,N22682,N22694);
or or1661(N20589,N22706,N22718);
or or1662(N20590,N22730,N22742);
or or1663(N20591,N22754,N22766);
or or1664(N20592,N22778,N22790);
or or1665(N20593,N22802,N22814);
or or1666(N20594,N22826,N22838);
or or1667(N20595,N22850,N22862);
or or1668(N20596,N22874,N22886);
or or1669(N20597,N22898,N22910);
or or1670(N20598,N22922,N22933);
or or1671(N20599,N22944,N22955);
or or1672(N20600,N22966,N22977);
or or1673(N20601,N22988,N22999);
or or1674(N20602,N23010,N23020);
or or1675(N20603,N23030,N23046);
or or1676(N20604,N23062,N23078);
or or1677(N20605,N23093,N23108);
or or1678(N20606,N23123,N23137);
or or1679(N20607,N23151,N23165);
or or1680(N20608,N23179,N23193);
or or1681(N20609,N23207,N23221);
or or1682(N20610,N23235,N23248);
or or1683(N20611,N23261,N23274);
or or1684(N20612,N23287,N23300);
or or1685(N20613,N23313,N23326);
or or1686(N20614,N23339,N23352);
or or1687(N20615,N23365,N23378);
or or1688(N20616,N23391,N23404);
or or1689(N20617,N23417,N23430);
or or1690(N20618,N23443,N23455);
or or1691(N20619,N23467,N23479);
or or1692(N20620,N23491,N23503);
or or1693(N20621,N23515,N23527);
or or1694(N20622,N23539,N23551);
or or1695(N20623,N23563,N23575);
or or1696(N20624,N23587,N23599);
or or1697(N20625,N23611,N23622);
or or1698(N20626,N23633,N23644);
or or1699(N20627,N23655,N23666);
or or1700(N20628,N23677,N23688);
or or1701(N20629,N23699,N23710);
or or1702(N20630,N23721,N23731);
or or1703(N20631,N23740,N23753);
or or1704(N20632,N23765,N23776);
or or1705(N20633,N23787,N23797);
or or1706(N20634,N23807,N23815);
or or1707(N23823,N23824,N23825);
or or1708(N23824,N23826,N23827);
or or1709(N23825,N23828,N23829);
or or1710(N23826,N23830,N23831);
or or1711(N23827,N23832,N23833);
or or1712(N23828,N23834,N23835);
or or1713(N23829,N23836,N23837);
or or1714(N23830,N23838,N23839);
or or1715(N23831,N23840,N23841);
or or1716(N23832,N23842,N23843);
or or1717(N23833,N23844,N23845);
or or1718(N23834,N23846,N23847);
or or1719(N23835,N23848,N23849);
or or1720(N23836,N23850,N23851);
or or1721(N23837,N23852,N23853);
or or1722(N23838,N23854,N23855);
or or1723(N23839,N23856,N23857);
or or1724(N23840,N23858,N23859);
or or1725(N23841,N23860,N23861);
or or1726(N23842,N23862,N23863);
or or1727(N23843,N23864,N23865);
or or1728(N23844,N23866,N23867);
or or1729(N23845,N23868,N23869);
or or1730(N23846,N23870,N23871);
or or1731(N23847,N23872,N23873);
or or1732(N23848,N23874,N23875);
or or1733(N23849,N23876,N23877);
or or1734(N23850,N23878,N23879);
or or1735(N23851,N23880,N23881);
or or1736(N23852,N23882,N23883);
or or1737(N23853,N23884,N23885);
or or1738(N23854,N23886,N23887);
or or1739(N23855,N23888,N23889);
or or1740(N23856,N23890,N23891);
or or1741(N23857,N23892,N23893);
or or1742(N23858,N23894,N23895);
or or1743(N23859,N23896,N23897);
or or1744(N23860,N23898,N23899);
or or1745(N23861,N23900,N23901);
or or1746(N23862,N23902,N23903);
or or1747(N23863,N23904,N23905);
or or1748(N23864,N23906,N23907);
or or1749(N23865,N23908,N23909);
or or1750(N23866,N23910,N23911);
or or1751(N23867,N23912,N23913);
or or1752(N23868,N23914,N23915);
or or1753(N23869,N23916,N23917);
or or1754(N23870,N23918,N23919);
or or1755(N23871,N23920,N23921);
or or1756(N23872,N23922,N23923);
or or1757(N23873,N23924,N23925);
or or1758(N23874,N23926,N23927);
or or1759(N23875,N23928,N23929);
or or1760(N23876,N23930,N23931);
or or1761(N23877,N23932,N23933);
or or1762(N23878,N23934,N23935);
or or1763(N23879,N23936,N23937);
or or1764(N23880,N23938,N23939);
or or1765(N23881,N23940,N23941);
or or1766(N23882,N23942,N23943);
or or1767(N23883,N23944,N23945);
or or1768(N23884,N23946,N23947);
or or1769(N23885,N23948,N23949);
or or1770(N23886,N23950,N23951);
or or1771(N23887,N23952,N23953);
or or1772(N23888,N23954,N23955);
or or1773(N23889,N23956,N23957);
or or1774(N23890,N23958,N23959);
or or1775(N23891,N23960,N23961);
or or1776(N23892,N23962,N23963);
or or1777(N23893,N23964,N23965);
or or1778(N23894,N23966,N23967);
or or1779(N23895,N23968,N23969);
or or1780(N23896,N23970,N23971);
or or1781(N23897,N23972,N23973);
or or1782(N23898,N23974,N23975);
or or1783(N23899,N23976,N23977);
or or1784(N23900,N23978,N23979);
or or1785(N23901,N23980,N23981);
or or1786(N23902,N23982,N23983);
or or1787(N23903,N23984,N23985);
or or1788(N23904,N23986,N23987);
or or1789(N23905,N23988,N23989);
or or1790(N23906,N23990,N23991);
or or1791(N23907,N23992,N23993);
or or1792(N23908,N23994,N23995);
or or1793(N23909,N23996,N23997);
or or1794(N23910,N23998,N23999);
or or1795(N23911,N24000,N24001);
or or1796(N23912,N24002,N24003);
or or1797(N23913,N24004,N24005);
or or1798(N23914,N24006,N24007);
or or1799(N23915,N24008,N24009);
or or1800(N23916,N24010,N24011);
or or1801(N23917,N24012,N24013);
or or1802(N23918,N24014,N24015);
or or1803(N23919,N24016,N24017);
or or1804(N23920,N24018,N24019);
or or1805(N23921,N24020,N24021);
or or1806(N23922,N24022,N24023);
or or1807(N23923,N24024,N24025);
or or1808(N23924,N24026,N24027);
or or1809(N23925,N24028,N24029);
or or1810(N23926,N24030,N24031);
or or1811(N23927,N24032,N24033);
or or1812(N23928,N24034,N24035);
or or1813(N23929,N24036,N24037);
or or1814(N23930,N24038,N24039);
or or1815(N23931,N24040,N24041);
or or1816(N23932,N24042,N24043);
or or1817(N23933,N24044,N24045);
or or1818(N23934,N24046,N24047);
or or1819(N23935,N24048,N24049);
or or1820(N23936,N24050,N24051);
or or1821(N23937,N24052,N24053);
or or1822(N23938,N24054,N24055);
or or1823(N23939,N24056,N24057);
or or1824(N23940,N24058,N24059);
or or1825(N23941,N24060,N24061);
or or1826(N23942,N24062,N24063);
or or1827(N23943,N24064,N24065);
or or1828(N23944,N24066,N24067);
or or1829(N23945,N24068,N24069);
or or1830(N23946,N24070,N24071);
or or1831(N23947,N24072,N24073);
or or1832(N23948,N24074,N24075);
or or1833(N23949,N24076,N24077);
or or1834(N23950,N24078,N24079);
or or1835(N23951,N24080,N24081);
or or1836(N23952,N24082,N24083);
or or1837(N23953,N24084,N24085);
or or1838(N23954,N24086,N24087);
or or1839(N23955,N24088,N24089);
or or1840(N23956,N24090,N24091);
or or1841(N23957,N24092,N24093);
or or1842(N23958,N24094,N24095);
or or1843(N23959,N24096,N24097);
or or1844(N23960,N24098,N24099);
or or1845(N23961,N24100,N24101);
or or1846(N23962,N24102,N24103);
or or1847(N23963,N24104,N24105);
or or1848(N23964,N24106,N24107);
or or1849(N23965,N24108,N24109);
or or1850(N23966,N24110,N24111);
or or1851(N23967,N24112,N24113);
or or1852(N23968,N24114,N24115);
or or1853(N23969,N24116,N24117);
or or1854(N23970,N24118,N24119);
or or1855(N23971,N24120,N24121);
or or1856(N23972,N24122,N24123);
or or1857(N23973,N24124,N24125);
or or1858(N23974,N24126,N24127);
or or1859(N23975,N24128,N24129);
or or1860(N23976,N24130,N24131);
or or1861(N23977,N24132,N24133);
or or1862(N23978,N24134,N24135);
or or1863(N23979,N24136,N24137);
or or1864(N23980,N24138,N24139);
or or1865(N23981,N24140,N24141);
or or1866(N23982,N24142,N24143);
or or1867(N23983,N24144,N24145);
or or1868(N23984,N24146,N24147);
or or1869(N23985,N24148,N24149);
or or1870(N23986,N24150,N24151);
or or1871(N23987,N24152,N24153);
or or1872(N23988,N24154,N24155);
or or1873(N23989,N24156,N24157);
or or1874(N23990,N24158,N24159);
or or1875(N23991,N24160,N24161);
or or1876(N23992,N24162,N24163);
or or1877(N23993,N24164,N24165);
or or1878(N23994,N24166,N24167);
or or1879(N23995,N24168,N24169);
or or1880(N23996,N24170,N24171);
or or1881(N23997,N24172,N24173);
or or1882(N23998,N24174,N24175);
or or1883(N23999,N24176,N24177);
or or1884(N24000,N24178,N24179);
or or1885(N24001,N24180,N24181);
or or1886(N24002,N24182,N24183);
or or1887(N24003,N24184,N24185);
or or1888(N24004,N24186,N24187);
or or1889(N24005,N24188,N24189);
or or1890(N24006,N24190,N24191);
or or1891(N24007,N24209,N24227);
or or1892(N24008,N24245,N24263);
or or1893(N24009,N24281,N24299);
or or1894(N24010,N24317,N24334);
or or1895(N24011,N24351,N24368);
or or1896(N24012,N24385,N24402);
or or1897(N24013,N24419,N24436);
or or1898(N24014,N24453,N24470);
or or1899(N24015,N24486,N24502);
or or1900(N24016,N24518,N24534);
or or1901(N24017,N24550,N24566);
or or1902(N24018,N24582,N24598);
or or1903(N24019,N24614,N24630);
or or1904(N24020,N24646,N24662);
or or1905(N24021,N24678,N24694);
or or1906(N24022,N24710,N24726);
or or1907(N24023,N24742,N24758);
or or1908(N24024,N24774,N24790);
or or1909(N24025,N24806,N24822);
or or1910(N24026,N24838,N24854);
or or1911(N24027,N24870,N24886);
or or1912(N24028,N24902,N24918);
or or1913(N24029,N24934,N24950);
or or1914(N24030,N24965,N24980);
or or1915(N24031,N24995,N25010);
or or1916(N24032,N25025,N25040);
or or1917(N24033,N25055,N25070);
or or1918(N24034,N25085,N25100);
or or1919(N24035,N25115,N25130);
or or1920(N24036,N25145,N25160);
or or1921(N24037,N25175,N25190);
or or1922(N24038,N25205,N25220);
or or1923(N24039,N25235,N25250);
or or1924(N24040,N25265,N25280);
or or1925(N24041,N25295,N25310);
or or1926(N24042,N25325,N25340);
or or1927(N24043,N25355,N25370);
or or1928(N24044,N25385,N25400);
or or1929(N24045,N25415,N25429);
or or1930(N24046,N25443,N25457);
or or1931(N24047,N25471,N25485);
or or1932(N24048,N25499,N25513);
or or1933(N24049,N25527,N25541);
or or1934(N24050,N25555,N25569);
or or1935(N24051,N25583,N25597);
or or1936(N24052,N25611,N25625);
or or1937(N24053,N25639,N25653);
or or1938(N24054,N25667,N25681);
or or1939(N24055,N25695,N25709);
or or1940(N24056,N25723,N25737);
or or1941(N24057,N25751,N25765);
or or1942(N24058,N25779,N25793);
or or1943(N24059,N25807,N25821);
or or1944(N24060,N25835,N25849);
or or1945(N24061,N25863,N25877);
or or1946(N24062,N25891,N25905);
or or1947(N24063,N25919,N25933);
or or1948(N24064,N25947,N25961);
or or1949(N24065,N25975,N25989);
or or1950(N24066,N26003,N26017);
or or1951(N24067,N26031,N26045);
or or1952(N24068,N26059,N26073);
or or1953(N24069,N26087,N26101);
or or1954(N24070,N26115,N26129);
or or1955(N24071,N26143,N26157);
or or1956(N24072,N26171,N26184);
or or1957(N24073,N26197,N26210);
or or1958(N24074,N26223,N26236);
or or1959(N24075,N26249,N26262);
or or1960(N24076,N26275,N26288);
or or1961(N24077,N26301,N26314);
or or1962(N24078,N26327,N26340);
or or1963(N24079,N26353,N26366);
or or1964(N24080,N26379,N26392);
or or1965(N24081,N26405,N26418);
or or1966(N24082,N26431,N26444);
or or1967(N24083,N26457,N26470);
or or1968(N24084,N26483,N26496);
or or1969(N24085,N26509,N26522);
or or1970(N24086,N26535,N26548);
or or1971(N24087,N26561,N26574);
or or1972(N24088,N26587,N26600);
or or1973(N24089,N26613,N26625);
or or1974(N24090,N26637,N26649);
or or1975(N24091,N26661,N26673);
or or1976(N24092,N26685,N26697);
or or1977(N24093,N26709,N26721);
or or1978(N24094,N26733,N26745);
or or1979(N24095,N26757,N26769);
or or1980(N24096,N26781,N26793);
or or1981(N24097,N26805,N26817);
or or1982(N24098,N26829,N26841);
or or1983(N24099,N26853,N26865);
or or1984(N24100,N26877,N26889);
or or1985(N24101,N26901,N26913);
or or1986(N24102,N26925,N26937);
or or1987(N24103,N26949,N26961);
or or1988(N24104,N26973,N26985);
or or1989(N24105,N26997,N27009);
or or1990(N24106,N27021,N27033);
or or1991(N24107,N27045,N27057);
or or1992(N24108,N27068,N27079);
or or1993(N24109,N27090,N27101);
or or1994(N24110,N27111,N27121);
or or1995(N24111,N27131,N27141);
or or1996(N24112,N27151,N27161);
or or1997(N24113,N27171,N27181);
or or1998(N24114,N27191,N27201);
or or1999(N24115,N27217,N27233);
or or2000(N24116,N27248,N27263);
or or2001(N24117,N27278,N27292);
or or2002(N24118,N27306,N27320);
or or2003(N24119,N27334,N27348);
or or2004(N24120,N27362,N27376);
or or2005(N24121,N27390,N27404);
or or2006(N24122,N27418,N27432);
or or2007(N24123,N27446,N27460);
or or2008(N24124,N27474,N27488);
or or2009(N24125,N27502,N27516);
or or2010(N24126,N27530,N27544);
or or2011(N24127,N27558,N27572);
or or2012(N24128,N27586,N27600);
or or2013(N24129,N27613,N27626);
or or2014(N24130,N27639,N27652);
or or2015(N24131,N27665,N27678);
or or2016(N24132,N27691,N27704);
or or2017(N24133,N27717,N27730);
or or2018(N24134,N27743,N27756);
or or2019(N24135,N27769,N27782);
or or2020(N24136,N27795,N27808);
or or2021(N24137,N27821,N27834);
or or2022(N24138,N27847,N27860);
or or2023(N24139,N27873,N27886);
or or2024(N24140,N27899,N27912);
or or2025(N24141,N27925,N27938);
or or2026(N24142,N27951,N27964);
or or2027(N24143,N27977,N27990);
or or2028(N24144,N28003,N28016);
or or2029(N24145,N28029,N28042);
or or2030(N24146,N28055,N28068);
or or2031(N24147,N28081,N28094);
or or2032(N24148,N28106,N28118);
or or2033(N24149,N28130,N28142);
or or2034(N24150,N28154,N28166);
or or2035(N24151,N28178,N28190);
or or2036(N24152,N28202,N28214);
or or2037(N24153,N28226,N28238);
or or2038(N24154,N28250,N28262);
or or2039(N24155,N28274,N28286);
or or2040(N24156,N28298,N28310);
or or2041(N24157,N28322,N28334);
or or2042(N24158,N28346,N28358);
or or2043(N24159,N28370,N28382);
or or2044(N24160,N28394,N28406);
or or2045(N24161,N28418,N28430);
or or2046(N24162,N28442,N28454);
or or2047(N24163,N28465,N28476);
or or2048(N24164,N28487,N28498);
or or2049(N24165,N28509,N28520);
or or2050(N24166,N28531,N28542);
or or2051(N24167,N28553,N28564);
or or2052(N24168,N28575,N28586);
or or2053(N24169,N28597,N28608);
or or2054(N24170,N28619,N28630);
or or2055(N24171,N28641,N28652);
or or2056(N24172,N28663,N28674);
or or2057(N24173,N28685,N28695);
or or2058(N24174,N28705,N28715);
or or2059(N24175,N28725,N28735);
or or2060(N24176,N28745,N28755);
or or2061(N24177,N28765,N28775);
or or2062(N24178,N28785,N28795);
or or2063(N24179,N28805,N28815);
or or2064(N24180,N28825,N28835);
or or2065(N24181,N28844,N28852);
or or2066(N24182,N28860,N28873);
or or2067(N24183,N28885,N28897);
or or2068(N24184,N28909,N28921);
or or2069(N24185,N28932,N28943);
or or2070(N24186,N28954,N28965);
or or2071(N24187,N28975,N28985);
or or2072(N24188,N28995,N29005);
or or2073(N24189,N29015,N29025);
or or2074(N24190,N29035,N29044);
or or2075(N29051,N29052,N29053);
or or2076(N29052,N29054,N29055);
or or2077(N29053,N29056,N29057);
or or2078(N29054,N29058,N29059);
or or2079(N29055,N29060,N29061);
or or2080(N29056,N29062,N29063);
or or2081(N29057,N29064,N29065);
or or2082(N29058,N29066,N29067);
or or2083(N29059,N29068,N29069);
or or2084(N29060,N29070,N29071);
or or2085(N29061,N29072,N29073);
or or2086(N29062,N29074,N29075);
or or2087(N29063,N29076,N29077);
or or2088(N29064,N29078,N29079);
or or2089(N29065,N29080,N29081);
or or2090(N29066,N29082,N29083);
or or2091(N29067,N29084,N29085);
or or2092(N29068,N29086,N29087);
or or2093(N29069,N29088,N29089);
or or2094(N29070,N29090,N29091);
or or2095(N29071,N29092,N29093);
or or2096(N29072,N29094,N29095);
or or2097(N29073,N29096,N29097);
or or2098(N29074,N29098,N29099);
or or2099(N29075,N29100,N29101);
or or2100(N29076,N29102,N29103);
or or2101(N29077,N29104,N29105);
or or2102(N29078,N29106,N29107);
or or2103(N29079,N29108,N29109);
or or2104(N29080,N29110,N29111);
or or2105(N29081,N29112,N29113);
or or2106(N29082,N29114,N29115);
or or2107(N29083,N29116,N29117);
or or2108(N29084,N29118,N29119);
or or2109(N29085,N29120,N29121);
or or2110(N29086,N29122,N29123);
or or2111(N29087,N29124,N29125);
or or2112(N29088,N29126,N29127);
or or2113(N29089,N29128,N29129);
or or2114(N29090,N29130,N29131);
or or2115(N29091,N29132,N29133);
or or2116(N29092,N29134,N29135);
or or2117(N29093,N29136,N29137);
or or2118(N29094,N29138,N29139);
or or2119(N29095,N29140,N29141);
or or2120(N29096,N29142,N29143);
or or2121(N29097,N29144,N29145);
or or2122(N29098,N29146,N29147);
or or2123(N29099,N29148,N29149);
or or2124(N29100,N29150,N29151);
or or2125(N29101,N29152,N29153);
or or2126(N29102,N29154,N29155);
or or2127(N29103,N29156,N29157);
or or2128(N29104,N29158,N29159);
or or2129(N29105,N29160,N29161);
or or2130(N29106,N29162,N29163);
or or2131(N29107,N29164,N29165);
or or2132(N29108,N29166,N29167);
or or2133(N29109,N29168,N29169);
or or2134(N29110,N29170,N29171);
or or2135(N29111,N29172,N29173);
or or2136(N29112,N29174,N29175);
or or2137(N29113,N29176,N29177);
or or2138(N29114,N29178,N29179);
or or2139(N29115,N29180,N29181);
or or2140(N29116,N29182,N29183);
or or2141(N29117,N29184,N29185);
or or2142(N29118,N29186,N29187);
or or2143(N29119,N29188,N29189);
or or2144(N29120,N29190,N29191);
or or2145(N29121,N29192,N29193);
or or2146(N29122,N29194,N29195);
or or2147(N29123,N29196,N29197);
or or2148(N29124,N29198,N29199);
or or2149(N29125,N29200,N29201);
or or2150(N29126,N29202,N29203);
or or2151(N29127,N29204,N29205);
or or2152(N29128,N29206,N29207);
or or2153(N29129,N29208,N29209);
or or2154(N29130,N29210,N29211);
or or2155(N29131,N29212,N29213);
or or2156(N29132,N29214,N29215);
or or2157(N29133,N29216,N29234);
or or2158(N29134,N29252,N29267);
or or2159(N29135,N29285,N29303);
or or2160(N29136,N29321,N29339);
or or2161(N29137,N29357,N29374);
or or2162(N29138,N29391,N29408);
or or2163(N29139,N29425,N29442);
or or2164(N29140,N29459,N29476);
or or2165(N29141,N29493,N29510);
or or2166(N29142,N29527,N29543);
or or2167(N29143,N29559,N29575);
or or2168(N29144,N29591,N29607);
or or2169(N29145,N29623,N29639);
or or2170(N29146,N29655,N29671);
or or2171(N29147,N29687,N29703);
or or2172(N29148,N29719,N29735);
or or2173(N29149,N29751,N29766);
or or2174(N29150,N29781,N29796);
or or2175(N29151,N29811,N29826);
or or2176(N29152,N29841,N29856);
or or2177(N29153,N29871,N29886);
or or2178(N29154,N29901,N29916);
or or2179(N29155,N29931,N29946);
or or2180(N29156,N29961,N29976);
or or2181(N29157,N29991,N30006);
or or2182(N29158,N30021,N30036);
or or2183(N29159,N30051,N30066);
or or2184(N29160,N30080,N30094);
or or2185(N29161,N30108,N30122);
or or2186(N29162,N30136,N30150);
or or2187(N29163,N30164,N30178);
or or2188(N29164,N30192,N30206);
or or2189(N29165,N30220,N30234);
or or2190(N29166,N30248,N30262);
or or2191(N29167,N30276,N30290);
or or2192(N29168,N30304,N30318);
or or2193(N29169,N30332,N30346);
or or2194(N29170,N30360,N30374);
or or2195(N29171,N30388,N30402);
or or2196(N29172,N30416,N30430);
or or2197(N29173,N30444,N30458);
or or2198(N29174,N30472,N30486);
or or2199(N29175,N30500,N30514);
or or2200(N29176,N30528,N30542);
or or2201(N29177,N30556,N30570);
or or2202(N29178,N30584,N30598);
or or2203(N29179,N30612,N30626);
or or2204(N29180,N30640,N30654);
or or2205(N29181,N30668,N30682);
or or2206(N29182,N30696,N30710);
or or2207(N29183,N30723,N30736);
or or2208(N29184,N30749,N30762);
or or2209(N29185,N30775,N30788);
or or2210(N29186,N30801,N30814);
or or2211(N29187,N30827,N30840);
or or2212(N29188,N30853,N30866);
or or2213(N29189,N30879,N30892);
or or2214(N29190,N30905,N30918);
or or2215(N29191,N30931,N30944);
or or2216(N29192,N30957,N30970);
or or2217(N29193,N30983,N30996);
or or2218(N29194,N31009,N31022);
or or2219(N29195,N31034,N31046);
or or2220(N29196,N31058,N31070);
or or2221(N29197,N31082,N31094);
or or2222(N29198,N31106,N31118);
or or2223(N29199,N31130,N31142);
or or2224(N29200,N31154,N31166);
or or2225(N29201,N31178,N31190);
or or2226(N29202,N31202,N31213);
or or2227(N29203,N31224,N31235);
or or2228(N29204,N31250,N31265);
or or2229(N29205,N31280,N31295);
or or2230(N29206,N31309,N31323);
or or2231(N29207,N31337,N31351);
or or2232(N29208,N31365,N31379);
or or2233(N29209,N31393,N31406);
or or2234(N29210,N31419,N31432);
or or2235(N29211,N31445,N31458);
or or2236(N29212,N31471,N31484);
or or2237(N29213,N31496,N31508);
or or2238(N29214,N31520,N31532);
or or2239(N29215,N31543,N31554);
or or2240(N31564,N31565,N31566);
or or2241(N31565,N31567,N31568);
or or2242(N31566,N31569,N31570);
or or2243(N31567,N31571,N31572);
or or2244(N31568,N31573,N31574);
or or2245(N31569,N31575,N31576);
or or2246(N31570,N31577,N31578);
or or2247(N31571,N31579,N31580);
or or2248(N31572,N31581,N31582);
or or2249(N31573,N31583,N31584);
or or2250(N31574,N31585,N31586);
or or2251(N31575,N31587,N31588);
or or2252(N31576,N31589,N31590);
or or2253(N31577,N31591,N31592);
or or2254(N31578,N31593,N31594);
or or2255(N31579,N31595,N31596);
or or2256(N31580,N31597,N31598);
or or2257(N31581,N31599,N31600);
or or2258(N31582,N31601,N31602);
or or2259(N31583,N31603,N31604);
or or2260(N31584,N31605,N31606);
or or2261(N31585,N31607,N31608);
or or2262(N31586,N31609,N31610);
or or2263(N31587,N31611,N31612);
or or2264(N31588,N31613,N31614);
or or2265(N31589,N31615,N31616);
or or2266(N31590,N31617,N31618);
or or2267(N31591,N31619,N31620);
or or2268(N31592,N31621,N31622);
or or2269(N31593,N31623,N31624);
or or2270(N31594,N31625,N31626);
or or2271(N31595,N31627,N31628);
or or2272(N31596,N31629,N31630);
or or2273(N31597,N31631,N31632);
or or2274(N31598,N31633,N31634);
or or2275(N31599,N31635,N31636);
or or2276(N31600,N31637,N31638);
or or2277(N31601,N31639,N31640);
or or2278(N31602,N31641,N31642);
or or2279(N31603,N31643,N31644);
or or2280(N31604,N31645,N31646);
or or2281(N31605,N31647,N31648);
or or2282(N31606,N31649,N31650);
or or2283(N31607,N31651,N31652);
or or2284(N31608,N31653,N31654);
or or2285(N31609,N31655,N31656);
or or2286(N31610,N31657,N31658);
or or2287(N31611,N31659,N31660);
or or2288(N31612,N31661,N31662);
or or2289(N31613,N31663,N31664);
or or2290(N31614,N31665,N31666);
or or2291(N31615,N31667,N31668);
or or2292(N31616,N31669,N31670);
or or2293(N31617,N31671,N31672);
or or2294(N31618,N31673,N31674);
or or2295(N31619,N31675,N31676);
or or2296(N31620,N31677,N31678);
or or2297(N31621,N31679,N31680);
or or2298(N31622,N31681,N31682);
or or2299(N31623,N31683,N31684);
or or2300(N31624,N31685,N31686);
or or2301(N31625,N31687,N31688);
or or2302(N31626,N31689,N31690);
or or2303(N31627,N31691,N31692);
or or2304(N31628,N31693,N31694);
or or2305(N31629,N31695,N31696);
or or2306(N31630,N31697,N31698);
or or2307(N31631,N31699,N31700);
or or2308(N31632,N31701,N31702);
or or2309(N31633,N31703,N31704);
or or2310(N31634,N31705,N31706);
or or2311(N31635,N31707,N31708);
or or2312(N31636,N31709,N31710);
or or2313(N31637,N31711,N31712);
or or2314(N31638,N31713,N31714);
or or2315(N31639,N31715,N31716);
or or2316(N31640,N31717,N31718);
or or2317(N31641,N31719,N31720);
or or2318(N31642,N31721,N31722);
or or2319(N31643,N31723,N31724);
or or2320(N31644,N31725,N31726);
or or2321(N31645,N31727,N31728);
or or2322(N31646,N31729,N31730);
or or2323(N31647,N31731,N31732);
or or2324(N31648,N31733,N31734);
or or2325(N31649,N31735,N31736);
or or2326(N31650,N31737,N31738);
or or2327(N31651,N31739,N31740);
or or2328(N31652,N31741,N31742);
or or2329(N31653,N31743,N31744);
or or2330(N31654,N31745,N31746);
or or2331(N31655,N31747,N31748);
or or2332(N31656,N31749,N31750);
or or2333(N31657,N31751,N31752);
or or2334(N31658,N31753,N31754);
or or2335(N31659,N31755,N31756);
or or2336(N31660,N31757,N31758);
or or2337(N31661,N31759,N31760);
or or2338(N31662,N31761,N31762);
or or2339(N31663,N31763,N31764);
or or2340(N31664,N31765,N31766);
or or2341(N31665,N31767,N31768);
or or2342(N31666,N31769,N31770);
or or2343(N31667,N31771,N31772);
or or2344(N31668,N31773,N31774);
or or2345(N31669,N31775,N31776);
or or2346(N31670,N31777,N31778);
or or2347(N31671,N31779,N31780);
or or2348(N31672,N31781,N31782);
or or2349(N31673,N31783,N31784);
or or2350(N31674,N31799,N31817);
or or2351(N31675,N31835,N31853);
or or2352(N31676,N31871,N31889);
or or2353(N31677,N31907,N31925);
or or2354(N31678,N31942,N31959);
or or2355(N31679,N31976,N31993);
or or2356(N31680,N32010,N32027);
or or2357(N31681,N32043,N32059);
or or2358(N31682,N32075,N32091);
or or2359(N31683,N32107,N32123);
or or2360(N31684,N32139,N32155);
or or2361(N31685,N32171,N32187);
or or2362(N31686,N32203,N32219);
or or2363(N31687,N32235,N32251);
or or2364(N31688,N32267,N32283);
or or2365(N31689,N32299,N32315);
or or2366(N31690,N32331,N32347);
or or2367(N31691,N32363,N32379);
or or2368(N31692,N32395,N32411);
or or2369(N31693,N32427,N32442);
or or2370(N31694,N32457,N32472);
or or2371(N31695,N32487,N32502);
or or2372(N31696,N32517,N32532);
or or2373(N31697,N32547,N32562);
or or2374(N31698,N32577,N32592);
or or2375(N31699,N32607,N32622);
or or2376(N31700,N32637,N32652);
or or2377(N31701,N32667,N32682);
or or2378(N31702,N32697,N32712);
or or2379(N31703,N32727,N32742);
or or2380(N31704,N32757,N32772);
or or2381(N31705,N32787,N32802);
or or2382(N31706,N32817,N32831);
or or2383(N31707,N32845,N32859);
or or2384(N31708,N32873,N32887);
or or2385(N31709,N32901,N32915);
or or2386(N31710,N32929,N32943);
or or2387(N31711,N32957,N32971);
or or2388(N31712,N32985,N32999);
or or2389(N31713,N33013,N33027);
or or2390(N31714,N33041,N33055);
or or2391(N31715,N33069,N33083);
or or2392(N31716,N33097,N33111);
or or2393(N31717,N33125,N33139);
or or2394(N31718,N33153,N33167);
or or2395(N31719,N33181,N33195);
or or2396(N31720,N33209,N33223);
or or2397(N31721,N33237,N33251);
or or2398(N31722,N33265,N33279);
or or2399(N31723,N33293,N33307);
or or2400(N31724,N33321,N33335);
or or2401(N31725,N33349,N33363);
or or2402(N31726,N33377,N33391);
or or2403(N31727,N33405,N33418);
or or2404(N31728,N33431,N33444);
or or2405(N31729,N33457,N33470);
or or2406(N31730,N33483,N33496);
or or2407(N31731,N33509,N33522);
or or2408(N31732,N33535,N33548);
or or2409(N31733,N33561,N33574);
or or2410(N31734,N33587,N33600);
or or2411(N31735,N33613,N33626);
or or2412(N31736,N33639,N33652);
or or2413(N31737,N33665,N33678);
or or2414(N31738,N33691,N33704);
or or2415(N31739,N33717,N33729);
or or2416(N31740,N33741,N33753);
or or2417(N31741,N33765,N33777);
or or2418(N31742,N33789,N33801);
or or2419(N31743,N33813,N33825);
or or2420(N31744,N33837,N33849);
or or2421(N31745,N33861,N33873);
or or2422(N31746,N33885,N33897);
or or2423(N31747,N33909,N33921);
or or2424(N31748,N33933,N33945);
or or2425(N31749,N33957,N33969);
or or2426(N31750,N33980,N33991);
or or2427(N31751,N34002,N34013);
or or2428(N31752,N34024,N34035);
or or2429(N31753,N34045,N34061);
or or2430(N31754,N34076,N34091);
or or2431(N31755,N34106,N34120);
or or2432(N31756,N34134,N34148);
or or2433(N31757,N34162,N34176);
or or2434(N31758,N34190,N34204);
or or2435(N31759,N34218,N34232);
or or2436(N31760,N34246,N34260);
or or2437(N31761,N34274,N34288);
or or2438(N31762,N34302,N34316);
or or2439(N31763,N34329,N34342);
or or2440(N31764,N34355,N34368);
or or2441(N31765,N34381,N34394);
or or2442(N31766,N34407,N34420);
or or2443(N31767,N34433,N34445);
or or2444(N31768,N34457,N34469);
or or2445(N31769,N34481,N34493);
or or2446(N31770,N34505,N34517);
or or2447(N31771,N34529,N34541);
or or2448(N31772,N34553,N34565);
or or2449(N31773,N34577,N34589);
or or2450(N31774,N34601,N34613);
or or2451(N31775,N34625,N34637);
or or2452(N31776,N34649,N34661);
or or2453(N31777,N34673,N34685);
or or2454(N31778,N34697,N34708);
or or2455(N31779,N34719,N34730);
or or2456(N31780,N34741,N34752);
or or2457(N31781,N34762,N34772);
or or2458(N31782,N34782,N34791);
or or2459(N31783,N34802,N34813);
or or2460(N34824,N34825,N34826);
or or2461(N34825,N34827,N34828);
or or2462(N34826,N34829,N34830);
or or2463(N34827,N34831,N34832);
or or2464(N34828,N34833,N34834);
or or2465(N34829,N34835,N34836);
or or2466(N34830,N34837,N34838);
or or2467(N34831,N34839,N34840);
or or2468(N34832,N34841,N34842);
or or2469(N34833,N34843,N34844);
or or2470(N34834,N34845,N34846);
or or2471(N34835,N34847,N34848);
or or2472(N34836,N34849,N34850);
or or2473(N34837,N34851,N34852);
or or2474(N34838,N34853,N34854);
or or2475(N34839,N34855,N34856);
or or2476(N34840,N34857,N34858);
or or2477(N34841,N34859,N34860);
or or2478(N34842,N34861,N34862);
or or2479(N34843,N34863,N34864);
or or2480(N34844,N34865,N34866);
or or2481(N34845,N34867,N34868);
or or2482(N34846,N34869,N34870);
or or2483(N34847,N34871,N34872);
or or2484(N34848,N34873,N34874);
or or2485(N34849,N34875,N34876);
or or2486(N34850,N34877,N34889);
or or2487(N34851,N34901,N34913);
or or2488(N34852,N34925,N34937);
or or2489(N34853,N34948,N34959);
or or2490(N34854,N34970,N34981);
or or2491(N34855,N34992,N35002);
or or2492(N34856,N35012,N35022);
or or2493(N34857,N35032,N35042);
or or2494(N34858,N35052,N35062);
or or2495(N34859,N35072,N35082);
or or2496(N34860,N35092,N35102);
or or2497(N34861,N35112,N35122);
or or2498(N34862,N35131,N35140);
or or2499(N34863,N35149,N35158);
or or2500(N34864,N35167,N35176);
or or2501(N34865,N35185,N35194);
or or2502(N34866,N35203,N35212);
or or2503(N34867,N35221,N35230);
or or2504(N34868,N35238,N35246);
or or2505(N34869,N35254,N35262);
or or2506(N34870,N35270,N35278);
or or2507(N34871,N35285,N35292);
or or2508(N34872,N35299,N35306);
or or2509(N34873,N35313,N35320);
or or2510(N34874,N35327,N35337);
or or2511(N34875,N35345,N35353);
or or2512(N34876,N35361,N35369);
or or2513(N35375,N35376,N35377);
or or2514(N35376,N35378,N35379);
or or2515(N35377,N35380,N35381);
or or2516(N35378,N35382,N35383);
or or2517(N35379,N35384,N35385);
or or2518(N35380,N35386,N35387);
or or2519(N35381,N35388,N35389);
or or2520(N35382,N35390,N35391);
or or2521(N35383,N35392,N35393);
or or2522(N35384,N35394,N35395);
or or2523(N35385,N35396,N35397);
or or2524(N35386,N35398,N35399);
or or2525(N35387,N35400,N35401);
or or2526(N35388,N35402,N35403);
or or2527(N35389,N35404,N35405);
or or2528(N35390,N35406,N35407);
or or2529(N35391,N35408,N35409);
or or2530(N35392,N35410,N35411);
or or2531(N35393,N35423,N35435);
or or2532(N35394,N35446,N35456);
or or2533(N35395,N35465,N35477);
or or2534(N35396,N35489,N35500);
or or2535(N35397,N35510,N35520);
or or2536(N35398,N35530,N35540);
or or2537(N35399,N35550,N35560);
or or2538(N35400,N35570,N35580);
or or2539(N35401,N35590,N35600);
or or2540(N35402,N35609,N35618);
or or2541(N35403,N35627,N35636);
or or2542(N35404,N35645,N35654);
or or2543(N35405,N35663,N35672);
or or2544(N35406,N35681,N35690);
or or2545(N35407,N35698,N35706);
or or2546(N35408,N35714,N35722);
or or2547(N35409,N35730,N35738);
or or2548(N35410,N35745,N35752);
or or2549(N35759,N35760,N35761);
or or2550(N35760,N35762,N35763);
or or2551(N35761,N35764,N35765);
or or2552(N35762,N35766,N35767);
or or2553(N35763,N35768,N35769);
or or2554(N35764,N35770,N35771);
or or2555(N35765,N35772,N35785);
or or2556(N35766,N35798,N35810);
or or2557(N35767,N35822,N35834);
or or2558(N35768,N35846,N35857);
or or2559(N35769,N35868,N35878);
or or2560(N35770,N35887,N35896);
or or2561(N35771,N35905,N35914);
or or2562(N35922,N35923,N35924);
or or2563(N35923,N35925,N35926);
or or2564(N35924,N35927,N35928);
or or2565(N35925,N35929,N35930);
or or2566(N35926,N35931,N35932);
or or2567(N35927,N35933,N35934);
or or2568(N35928,N35935,N35936);
or or2569(N35929,N35937,N35938);
or or2570(N35930,N35939,N35940);
or or2571(N35931,N35941,N35942);
or or2572(N35932,N35943,N35944);
or or2573(N35933,N35945,N35946);
or or2574(N35934,N35947,N35948);
or or2575(N35935,N35949,N35950);
or or2576(N35936,N35951,N35952);
or or2577(N35937,N35953,N35954);
or or2578(N35938,N35955,N35956);
or or2579(N35939,N35957,N35958);
or or2580(N35940,N35959,N35960);
or or2581(N35941,N35961,N35962);
or or2582(N35942,N35963,N35964);
or or2583(N35943,N35965,N35966);
or or2584(N35944,N35979,N35991);
or or2585(N35945,N36003,N36014);
or or2586(N35946,N36024,N36033);
or or2587(N35947,N36045,N36057);
or or2588(N35948,N36068,N36079);
or or2589(N35949,N36089,N36099);
or or2590(N35950,N36109,N36119);
or or2591(N35951,N36129,N36139);
or or2592(N35952,N36149,N36159);
or or2593(N35953,N36169,N36179);
or or2594(N35954,N36189,N36199);
or or2595(N35955,N36209,N36218);
or or2596(N35956,N36227,N36236);
or or2597(N35957,N36245,N36254);
or or2598(N35958,N36262,N36270);
or or2599(N35959,N36278,N36286);
or or2600(N35960,N36294,N36302);
or or2601(N35961,N36310,N36318);
or or2602(N35962,N36326,N36334);
or or2603(N35963,N36342,N36350);
or or2604(N35964,N36358,N36365);
or or2605(N35965,N36372,N36379);
or or2606(N36387,N36388,N36389);
or or2607(N36388,N36390,N36391);
or or2608(N36389,N36392,N36393);
or or2609(N36390,N36394,N36395);
or or2610(N36391,N36396,N36397);
or or2611(N36392,N36398,N36399);
or or2612(N36393,N36400,N36401);
or or2613(N36394,N36402,N36403);
or or2614(N36395,N36404,N36405);
or or2615(N36396,N36406,N36407);
or or2616(N36397,N36408,N36422);
or or2617(N36398,N36435,N36448);
or or2618(N36399,N36461,N36473);
or or2619(N36400,N36485,N36496);
or or2620(N36401,N36507,N36518);
or or2621(N36402,N36529,N36540);
or or2622(N36403,N36551,N36561);
or or2623(N36404,N36569,N36580);
or or2624(N36405,N36591,N36601);
or or2625(N36406,N36611,N36620);
or or2626(N36407,N36629,N36638);
or or2627(N36646,N36647,N36648);
or or2628(N36647,N36649,N36650);
or or2629(N36648,N36651,N36652);
or or2630(N36649,N36653,N36654);
or or2631(N36650,N36655,N36656);
or or2632(N36651,N36657,N36658);
or or2633(N36652,N36659,N36660);
or or2634(N36653,N36661,N36662);
or or2635(N36654,N36663,N36664);
or or2636(N36655,N36665,N36666);
or or2637(N36656,N36667,N36668);
or or2638(N36657,N36669,N36670);
or or2639(N36658,N36671,N36672);
or or2640(N36659,N36673,N36674);
or or2641(N36660,N36675,N36676);
or or2642(N36661,N36677,N36678);
or or2643(N36662,N36679,N36680);
or or2644(N36663,N36681,N36682);
or or2645(N36664,N36683,N36684);
or or2646(N36665,N36685,N36686);
or or2647(N36666,N36687,N36688);
or or2648(N36667,N36689,N36690);
or or2649(N36668,N36691,N36692);
or or2650(N36669,N36693,N36707);
or or2651(N36670,N36719,N36731);
or or2652(N36671,N36742,N36752);
or or2653(N36672,N36764,N36776);
or or2654(N36673,N36788,N36799);
or or2655(N36674,N36810,N36821);
or or2656(N36675,N36832,N36842);
or or2657(N36676,N36852,N36862);
or or2658(N36677,N36872,N36882);
or or2659(N36678,N36892,N36902);
or or2660(N36679,N36912,N36922);
or or2661(N36680,N36932,N36942);
or or2662(N36681,N36952,N36961);
or or2663(N36682,N36970,N36979);
or or2664(N36683,N36988,N36997);
or or2665(N36684,N37006,N37015);
or or2666(N36685,N37023,N37031);
or or2667(N36686,N37039,N37047);
or or2668(N36687,N37055,N37063);
or or2669(N36688,N37071,N37079);
or or2670(N36689,N37087,N37095);
or or2671(N36690,N37103,N37111);
or or2672(N36691,N37118,N37125);
or or2673(N36692,N37132,N37139);

not not0(N420,in0);
not not1(N421,in1);
not not2(N422,R0);
not not3(N423,R2);
not not4(N437,in1);
not not5(N438,R0);
not not6(N439,R1);
not not7(N440,R2);
not not8(N441,R3);
not not9(N454,in1);
not not10(N455,in2);
not not11(N456,R1);
not not12(N457,R2);
not not13(N458,R3);
not not14(N471,in2);
not not15(N472,R0);
not not16(N473,R1);
not not17(N474,R2);
not not18(N475,R3);
not not19(N488,in2);
not not20(N489,R0);
not not21(N490,R1);
not not22(N491,R2);
not not23(N505,in1);
not not24(N506,R0);
not not25(N507,R1);
not not26(N508,R2);
not not27(N522,in0);
not not28(N523,in1);
not not29(N524,in2);
not not30(N525,R0);
not not31(N526,R1);
not not32(N539,in0);
not not33(N540,in1);
not not34(N541,in2);
not not35(N542,R0);
not not36(N543,R1);
not not37(N556,in0);
not not38(N557,in1);
not not39(N558,in2);
not not40(N559,R0);
not not41(N560,R1);
not not42(N561,R2);
not not43(N573,in0);
not not44(N574,in1);
not not45(N575,in2);
not not46(N576,R0);
not not47(N577,R1);
not not48(N578,R3);
not not49(N590,in0);
not not50(N591,in1);
not not51(N592,in2);
not not52(N593,R0);
not not53(N594,R1);
not not54(N607,in0);
not not55(N608,in1);
not not56(N609,in2);
not not57(N610,R0);
not not58(N611,R1);
not not59(N624,in0);
not not60(N625,R1);
not not61(N626,R2);
not not62(N640,R0);
not not63(N641,R1);
not not64(N642,R2);
not not65(N643,R3);
not not66(N656,in0);
not not67(N657,R0);
not not68(N658,R1);
not not69(N659,R2);
not not70(N672,in0);
not not71(N673,in1);
not not72(N674,R0);
not not73(N675,R3);
not not74(N688,in0);
not not75(N689,in1);
not not76(N690,R3);
not not77(N704,in0);
not not78(N705,R1);
not not79(N706,R2);
not not80(N720,in0);
not not81(N721,in1);
not not82(N722,R1);
not not83(N723,R2);
not not84(N724,R3);
not not85(N736,in1);
not not86(N737,in2);
not not87(N738,R0);
not not88(N739,R1);
not not89(N740,R2);
not not90(N752,in0);
not not91(N753,in2);
not not92(N754,R0);
not not93(N755,R1);
not not94(N756,R2);
not not95(N768,in0);
not not96(N769,in1);
not not97(N770,R0);
not not98(N771,R3);
not not99(N784,in1);
not not100(N785,in2);
not not101(N786,R0);
not not102(N787,R1);
not not103(N788,R2);
not not104(N800,in0);
not not105(N801,in1);
not not106(N802,R0);
not not107(N803,R1);
not not108(N816,in1);
not not109(N817,in2);
not not110(N818,R0);
not not111(N819,R3);
not not112(N831,R1);
not not113(N832,R2);
not not114(N833,R3);
not not115(N846,R1);
not not116(N847,R2);
not not117(N848,R3);
not not118(N861,in0);
not not119(N862,in1);
not not120(N863,R1);
not not121(N864,R2);
not not122(N876,in1);
not not123(N877,R2);
not not124(N878,R3);
not not125(N891,in0);
not not126(N892,R1);
not not127(N893,R2);
not not128(N906,in0);
not not129(N907,R0);
not not130(N921,in0);
not not131(N922,R0);
not not132(N923,R1);
not not133(N924,R2);
not not134(N925,R3);
not not135(N936,in0);
not not136(N937,in1);
not not137(N938,R1);
not not138(N951,in2);
not not139(N952,R0);
not not140(N953,R1);
not not141(N954,R3);
not not142(N966,in1);
not not143(N967,R0);
not not144(N968,R1);
not not145(N969,R3);
not not146(N981,in2);
not not147(N982,R0);
not not148(N983,R1);
not not149(N984,R2);
not not150(N996,in0);
not not151(N997,in1);
not not152(N998,R1);
not not153(N1011,in1);
not not154(N1012,R0);
not not155(N1013,R1);
not not156(N1026,in0);
not not157(N1027,in2);
not not158(N1028,R0);
not not159(N1029,R3);
not not160(N1041,in0);
not not161(N1042,R0);
not not162(N1043,R1);
not not163(N1044,R3);
not not164(N1056,in0);
not not165(N1057,in1);
not not166(N1058,R1);
not not167(N1071,in0);
not not168(N1072,in2);
not not169(N1073,R1);
not not170(N1086,in0);
not not171(N1087,in2);
not not172(N1088,R1);
not not173(N1089,R3);
not not174(N1101,in0);
not not175(N1102,R0);
not not176(N1103,R1);
not not177(N1104,R2);
not not178(N1116,in0);
not not179(N1117,in1);
not not180(N1118,in2);
not not181(N1119,R1);
not not182(N1131,in0);
not not183(N1132,R1);
not not184(N1133,R2);
not not185(N1134,R3);
not not186(N1146,in0);
not not187(N1147,in1);
not not188(N1148,R0);
not not189(N1161,in0);
not not190(N1162,in1);
not not191(N1163,R1);
not not192(N1176,in1);
not not193(N1177,in2);
not not194(N1178,R2);
not not195(N1179,R3);
not not196(N1191,in0);
not not197(N1192,in1);
not not198(N1193,in2);
not not199(N1194,R0);
not not200(N1195,R1);
not not201(N1206,in0);
not not202(N1207,in2);
not not203(N1208,R2);
not not204(N1209,R3);
not not205(N1221,in0);
not not206(N1222,in1);
not not207(N1223,R1);
not not208(N1224,R2);
not not209(N1236,in0);
not not210(N1237,in1);
not not211(N1238,R2);
not not212(N1251,in2);
not not213(N1252,R0);
not not214(N1253,R1);
not not215(N1254,R2);
not not216(N1266,in0);
not not217(N1267,in1);
not not218(N1268,in2);
not not219(N1269,R0);
not not220(N1270,R2);
not not221(N1281,in1);
not not222(N1282,R0);
not not223(N1283,R1);
not not224(N1284,R2);
not not225(N1296,in0);
not not226(N1297,R0);
not not227(N1298,R1);
not not228(N1299,R2);
not not229(N1311,in0);
not not230(N1312,in1);
not not231(N1313,R0);
not not232(N1314,R1);
not not233(N1326,in0);
not not234(N1327,in2);
not not235(N1328,R0);
not not236(N1329,R1);
not not237(N1341,in0);
not not238(N1342,in1);
not not239(N1343,in2);
not not240(N1344,R2);
not not241(N1356,in0);
not not242(N1357,R0);
not not243(N1358,R1);
not not244(N1370,in0);
not not245(N1384,in0);
not not246(N1385,in1);
not not247(N1386,R1);
not not248(N1398,in0);
not not249(N1399,R0);
not not250(N1400,R1);
not not251(N1401,R2);
not not252(N1412,in2);
not not253(N1413,R0);
not not254(N1414,R3);
not not255(N1426,in0);
not not256(N1427,in1);
not not257(N1428,R0);
not not258(N1440,in0);
not not259(N1441,R0);
not not260(N1454,in0);
not not261(N1455,in1);
not not262(N1456,R2);
not not263(N1468,R0);
not not264(N1469,R1);
not not265(N1470,R2);
not not266(N1482,in0);
not not267(N1483,R1);
not not268(N1484,R2);
not not269(N1496,in0);
not not270(N1497,in1);
not not271(N1498,in2);
not not272(N1510,in1);
not not273(N1511,in2);
not not274(N1512,R1);
not not275(N1513,R3);
not not276(N1524,in0);
not not277(N1525,R0);
not not278(N1526,R2);
not not279(N1538,in1);
not not280(N1539,R0);
not not281(N1540,R1);
not not282(N1541,R3);
not not283(N1552,in0);
not not284(N1553,in1);
not not285(N1554,R0);
not not286(N1566,in0);
not not287(N1567,R1);
not not288(N1580,in0);
not not289(N1581,in1);
not not290(N1594,in0);
not not291(N1595,R1);
not not292(N1596,R3);
not not293(N1608,in0);
not not294(N1609,in2);
not not295(N1610,R1);
not not296(N1611,R2);
not not297(N1622,in0);
not not298(N1623,R0);
not not299(N1624,R1);
not not300(N1625,R3);
not not301(N1636,in0);
not not302(N1637,in1);
not not303(N1638,R2);
not not304(N1650,in0);
not not305(N1651,in2);
not not306(N1652,R1);
not not307(N1653,R2);
not not308(N1664,in0);
not not309(N1665,R1);
not not310(N1666,R2);
not not311(N1678,in1);
not not312(N1679,in2);
not not313(N1680,R0);
not not314(N1692,in1);
not not315(N1693,in2);
not not316(N1694,R0);
not not317(N1695,R1);
not not318(N1706,in0);
not not319(N1707,in2);
not not320(N1708,R2);
not not321(N1720,in0);
not not322(N1721,in1);
not not323(N1722,R2);
not not324(N1734,in1);
not not325(N1735,R1);
not not326(N1747,R0);
not not327(N1748,R1);
not not328(N1760,in1);
not not329(N1761,R3);
not not330(N1773,R0);
not not331(N1774,R1);
not not332(N1786,in1);
not not333(N1787,R1);
not not334(N1788,R3);
not not335(N1799,in0);
not not336(N1800,in2);
not not337(N1801,R1);
not not338(N1812,R3);
not not339(N1825,in1);
not not340(N1826,R0);
not not341(N1838,R0);
not not342(N1839,R3);
not not343(N1851,in2);
not not344(N1852,R1);
not not345(N1864,R0);
not not346(N1865,R3);
not not347(N1877,in0);
not not348(N1878,in1);
not not349(N1879,R1);
not not350(N1890,in0);
not not351(N1891,in1);
not not352(N1892,R1);
not not353(N1893,R2);
not not354(N1903,R2);
not not355(N1916,R1);
not not356(N1917,R3);
not not357(N1929,in0);
not not358(N1942,R0);
not not359(N1943,R3);
not not360(N1955,in1);
not not361(N1968,R1);
not not362(N1981,R1);
not not363(N1982,R2);
not not364(N1994,in0);
not not365(N1995,R1);
not not366(N2007,in1);
not not367(N2008,R1);
not not368(N2020,in2);
not not369(N2021,R1);
not not370(N2033,in0);
not not371(N2034,R2);
not not372(N2046,in0);
not not373(N2047,R1);
not not374(N2048,R2);
not not375(N2059,in0);
not not376(N2060,in1);
not not377(N2061,R1);
not not378(N2062,R2);
not not379(N2072,in0);
not not380(N2073,in2);
not not381(N2074,R2);
not not382(N2085,R1);
not not383(N2086,R2);
not not384(N2098,in1);
not not385(N2099,R2);
not not386(N2111,in1);
not not387(N2112,R2);
not not388(N2124,R2);
not not389(N2125,R3);
not not390(N2137,in0);
not not391(N2138,R2);
not not392(N2150,in1);
not not393(N2151,in2);
not not394(N2152,R3);
not not395(N2163,in0);
not not396(N2164,in1);
not not397(N2165,R3);
not not398(N2176,in0);
not not399(N2177,R0);
not not400(N2178,R1);
not not401(N2189,in0);
not not402(N2190,in1);
not not403(N2191,R1);
not not404(N2202,in0);
not not405(N2203,in2);
not not406(N2204,R0);
not not407(N2205,R1);
not not408(N2215,in2);
not not409(N2216,R0);
not not410(N2228,in2);
not not411(N2229,R0);
not not412(N2230,R1);
not not413(N2241,R2);
not not414(N2242,R3);
not not415(N2254,in0);
not not416(N2255,R0);
not not417(N2256,R1);
not not418(N2267,in0);
not not419(N2268,R0);
not not420(N2269,R1);
not not421(N2270,R2);
not not422(N2280,in1);
not not423(N2281,R0);
not not424(N2282,R1);
not not425(N2293,in2);
not not426(N2294,R0);
not not427(N2295,R1);
not not428(N2306,in1);
not not429(N2307,R0);
not not430(N2308,R1);
not not431(N2319,in2);
not not432(N2320,R0);
not not433(N2321,R1);
not not434(N2332,in0);
not not435(N2333,R2);
not not436(N2345,in2);
not not437(N2357,in2);
not not438(N2358,R0);
not not439(N2369,in0);
not not440(N2370,R0);
not not441(N2393,in0);
not not442(N2394,R1);
not not443(N2395,R2);
not not444(N2405,in0);
not not445(N2406,R1);
not not446(N2417,in0);
not not447(N2418,in1);
not not448(N2429,R1);
not not449(N2430,R2);
not not450(N2441,in0);
not not451(N2442,R1);
not not452(N2453,in1);
not not453(N2454,R2);
not not454(N2465,in0);
not not455(N2466,R2);
not not456(N2489,in2);
not not457(N2490,R0);
not not458(N2501,in0);
not not459(N2513,R2);
not not460(N2525,R1);
not not461(N2526,R2);
not not462(N2537,R0);
not not463(N2549,in0);
not not464(N2550,R2);
not not465(N2561,in1);
not not466(N2562,in2);
not not467(N2584,R0);
not not468(N2606,R0);
not not469(N2617,in2);
not not470(N2618,R0);
not not471(N2628,R1);
not not472(N2639,R2);
not not473(N2661,in0);
not not474(N2662,R2);
not not475(N2672,R0);
not not476(N2694,R1);
not not477(N2705,R0);
not not478(N2706,R2);
not not479(N2716,in1);
not not480(N2727,R3);
not not481(N2738,R3);
not not482(N2749,in2);
not not483(N2760,R0);
not not484(N2761,R1);
not not485(N2771,R1);
not not486(N2810,in1);
not not487(N2811,R0);
not not488(N2812,R1);
not not489(N2813,R2);
not not490(N2814,R3);
not not491(N2815,R4);
not not492(N2816,R5);
not not493(N2826,in1);
not not494(N2827,R0);
not not495(N2828,R1);
not not496(N2829,R3);
not not497(N2830,R4);
not not498(N2831,R5);
not not499(N2842,in1);
not not500(N2843,R0);
not not501(N2844,R1);
not not502(N2845,R2);
not not503(N2846,R3);
not not504(N2847,R4);
not not505(N2858,in1);
not not506(N2859,in2);
not not507(N2860,R0);
not not508(N2861,R2);
not not509(N2862,R4);
not not510(N2863,R5);
not not511(N2874,in0);
not not512(N2875,R0);
not not513(N2876,R2);
not not514(N2877,R3);
not not515(N2878,R4);
not not516(N2879,R5);
not not517(N2889,in2);
not not518(N2890,R1);
not not519(N2891,R2);
not not520(N2892,R3);
not not521(N2893,R5);
not not522(N2904,in0);
not not523(N2905,in1);
not not524(N2906,in2);
not not525(N2907,R3);
not not526(N2908,R4);
not not527(N2919,in1);
not not528(N2920,in2);
not not529(N2921,R1);
not not530(N2922,R2);
not not531(N2923,R4);
not not532(N2934,in0);
not not533(N2935,in1);
not not534(N2936,R1);
not not535(N2937,R2);
not not536(N2938,R3);
not not537(N2939,R5);
not not538(N2949,in1);
not not539(N2950,in2);
not not540(N2951,R0);
not not541(N2952,R2);
not not542(N2953,R4);
not not543(N2964,in1);
not not544(N2965,in2);
not not545(N2966,R0);
not not546(N2967,R1);
not not547(N2968,R2);
not not548(N2969,R4);
not not549(N2979,R2);
not not550(N2980,R3);
not not551(N2981,R4);
not not552(N2982,R5);
not not553(N2993,in0);
not not554(N2994,R0);
not not555(N2995,R1);
not not556(N2996,R3);
not not557(N2997,R4);
not not558(N3007,in1);
not not559(N3008,R1);
not not560(N3009,R2);
not not561(N3010,R3);
not not562(N3011,R4);
not not563(N3021,in1);
not not564(N3022,in2);
not not565(N3023,R0);
not not566(N3024,R4);
not not567(N3035,in1);
not not568(N3036,R0);
not not569(N3037,R3);
not not570(N3038,R4);
not not571(N3049,in1);
not not572(N3050,R1);
not not573(N3051,R4);
not not574(N3052,R5);
not not575(N3063,in2);
not not576(N3064,R0);
not not577(N3065,R1);
not not578(N3066,R2);
not not579(N3067,R5);
not not580(N3077,in1);
not not581(N3078,R0);
not not582(N3079,R1);
not not583(N3080,R4);
not not584(N3081,R5);
not not585(N3091,in2);
not not586(N3092,R0);
not not587(N3093,R1);
not not588(N3094,R4);
not not589(N3095,R5);
not not590(N3105,in1);
not not591(N3106,R0);
not not592(N3107,R1);
not not593(N3108,R4);
not not594(N3109,R5);
not not595(N3119,in0);
not not596(N3120,in1);
not not597(N3121,in2);
not not598(N3122,R3);
not not599(N3123,R4);
not not600(N3133,in1);
not not601(N3134,R0);
not not602(N3135,R1);
not not603(N3136,R3);
not not604(N3147,in2);
not not605(N3148,R0);
not not606(N3149,R1);
not not607(N3150,R3);
not not608(N3161,in1);
not not609(N3162,in2);
not not610(N3163,R0);
not not611(N3164,R5);
not not612(N3175,in0);
not not613(N3176,in2);
not not614(N3177,R1);
not not615(N3178,R2);
not not616(N3179,R3);
not not617(N3189,in0);
not not618(N3190,in1);
not not619(N3191,R1);
not not620(N3192,R2);
not not621(N3193,R3);
not not622(N3194,R4);
not not623(N3203,R0);
not not624(N3204,R1);
not not625(N3205,R2);
not not626(N3206,R3);
not not627(N3217,in0);
not not628(N3218,in2);
not not629(N3219,R3);
not not630(N3220,R5);
not not631(N3231,in0);
not not632(N3232,in2);
not not633(N3233,R3);
not not634(N3234,R4);
not not635(N3245,in1);
not not636(N3246,in2);
not not637(N3247,R3);
not not638(N3248,R4);
not not639(N3259,in0);
not not640(N3260,in1);
not not641(N3261,R2);
not not642(N3262,R4);
not not643(N3263,R5);
not not644(N3273,in0);
not not645(N3274,in2);
not not646(N3275,R0);
not not647(N3276,R1);
not not648(N3277,R3);
not not649(N3287,in1);
not not650(N3288,R0);
not not651(N3289,R3);
not not652(N3290,R5);
not not653(N3301,in0);
not not654(N3302,in1);
not not655(N3303,R3);
not not656(N3304,R4);
not not657(N3305,R5);
not not658(N3315,in0);
not not659(N3316,in2);
not not660(N3317,R2);
not not661(N3318,R4);
not not662(N3319,R5);
not not663(N3329,in1);
not not664(N3330,in2);
not not665(N3331,R4);
not not666(N3332,R5);
not not667(N3343,in2);
not not668(N3344,R0);
not not669(N3345,R1);
not not670(N3346,R4);
not not671(N3357,in1);
not not672(N3358,in2);
not not673(N3359,R0);
not not674(N3360,R1);
not not675(N3361,R3);
not not676(N3371,in2);
not not677(N3372,R1);
not not678(N3373,R2);
not not679(N3374,R3);
not not680(N3375,R4);
not not681(N3385,in1);
not not682(N3386,in2);
not not683(N3387,R0);
not not684(N3388,R3);
not not685(N3399,in0);
not not686(N3400,R2);
not not687(N3401,R3);
not not688(N3402,R4);
not not689(N3403,R5);
not not690(N3413,in1);
not not691(N3414,R1);
not not692(N3415,R2);
not not693(N3416,R4);
not not694(N3427,in2);
not not695(N3428,R1);
not not696(N3429,R2);
not not697(N3430,R4);
not not698(N3441,in0);
not not699(N3442,R0);
not not700(N3443,R1);
not not701(N3444,R3);
not not702(N3455,in0);
not not703(N3456,in1);
not not704(N3457,R3);
not not705(N3458,R5);
not not706(N3469,in2);
not not707(N3470,R1);
not not708(N3471,R2);
not not709(N3472,R3);
not not710(N3473,R4);
not not711(N3474,R5);
not not712(N3483,R0);
not not713(N3484,R4);
not not714(N3485,R5);
not not715(N3496,in1);
not not716(N3497,R4);
not not717(N3498,R5);
not not718(N3509,in2);
not not719(N3510,R0);
not not720(N3511,R5);
not not721(N3522,R0);
not not722(N3523,R1);
not not723(N3524,R4);
not not724(N3535,R1);
not not725(N3536,R2);
not not726(N3537,R3);
not not727(N3538,R4);
not not728(N3548,in1);
not not729(N3549,R3);
not not730(N3550,R4);
not not731(N3561,R1);
not not732(N3562,R2);
not not733(N3563,R4);
not not734(N3574,in0);
not not735(N3575,R0);
not not736(N3576,R2);
not not737(N3577,R4);
not not738(N3587,in0);
not not739(N3588,in1);
not not740(N3589,R0);
not not741(N3590,R4);
not not742(N3600,in1);
not not743(N3601,R1);
not not744(N3602,R2);
not not745(N3603,R3);
not not746(N3613,in0);
not not747(N3614,in2);
not not748(N3615,R0);
not not749(N3626,in0);
not not750(N3627,in1);
not not751(N3628,R0);
not not752(N3639,in1);
not not753(N3640,R1);
not not754(N3641,R4);
not not755(N3652,in1);
not not756(N3653,R1);
not not757(N3654,R3);
not not758(N3655,R4);
not not759(N3665,in1);
not not760(N3666,in2);
not not761(N3667,R2);
not not762(N3678,in1);
not not763(N3679,R2);
not not764(N3680,R3);
not not765(N3681,R5);
not not766(N3691,in0);
not not767(N3692,in2);
not not768(N3693,R1);
not not769(N3694,R2);
not not770(N3695,R3);
not not771(N3704,in0);
not not772(N3705,R1);
not not773(N3706,R2);
not not774(N3717,in0);
not not775(N3718,R1);
not not776(N3719,R2);
not not777(N3730,in1);
not not778(N3731,in2);
not not779(N3732,R0);
not not780(N3733,R1);
not not781(N3734,R2);
not not782(N3743,R0);
not not783(N3744,R2);
not not784(N3745,R4);
not not785(N3756,R0);
not not786(N3757,R2);
not not787(N3758,R4);
not not788(N3769,in0);
not not789(N3770,R0);
not not790(N3771,R2);
not not791(N3772,R4);
not not792(N3782,in0);
not not793(N3783,in2);
not not794(N3784,R1);
not not795(N3785,R3);
not not796(N3786,R4);
not not797(N3795,R0);
not not798(N3796,R1);
not not799(N3797,R2);
not not800(N3798,R4);
not not801(N3808,R0);
not not802(N3809,R1);
not not803(N3810,R2);
not not804(N3811,R5);
not not805(N3821,in2);
not not806(N3822,R0);
not not807(N3823,R1);
not not808(N3824,R3);
not not809(N3834,in0);
not not810(N3835,R0);
not not811(N3836,R3);
not not812(N3847,in1);
not not813(N3848,R1);
not not814(N3849,R3);
not not815(N3850,R4);
not not816(N3860,R1);
not not817(N3861,R3);
not not818(N3862,R4);
not not819(N3863,R5);
not not820(N3873,in1);
not not821(N3874,in2);
not not822(N3875,R1);
not not823(N3876,R3);
not not824(N3886,in0);
not not825(N3887,in2);
not not826(N3888,R0);
not not827(N3889,R5);
not not828(N3899,in1);
not not829(N3900,R0);
not not830(N3901,R2);
not not831(N3902,R4);
not not832(N3912,in2);
not not833(N3913,R3);
not not834(N3914,R4);
not not835(N3925,R0);
not not836(N3926,R1);
not not837(N3927,R4);
not not838(N3928,R5);
not not839(N3938,in0);
not not840(N3939,in1);
not not841(N3940,R3);
not not842(N3941,R4);
not not843(N3951,in2);
not not844(N3952,R1);
not not845(N3953,R4);
not not846(N3964,in0);
not not847(N3965,in1);
not not848(N3966,in2);
not not849(N3967,R4);
not not850(N3977,in2);
not not851(N3978,R1);
not not852(N3989,R0);
not not853(N3990,R3);
not not854(N3991,R4);
not not855(N4001,R3);
not not856(N4002,R5);
not not857(N4013,R0);
not not858(N4014,R1);
not not859(N4015,R2);
not not860(N4016,R4);
not not861(N4025,in1);
not not862(N4026,in2);
not not863(N4027,R5);
not not864(N4037,in1);
not not865(N4038,in2);
not not866(N4039,R1);
not not867(N4040,R5);
not not868(N4049,in1);
not not869(N4050,R3);
not not870(N4051,R4);
not not871(N4061,in1);
not not872(N4062,in2);
not not873(N4063,R1);
not not874(N4064,R2);
not not875(N4073,R0);
not not876(N4074,R3);
not not877(N4085,R0);
not not878(N4086,R3);
not not879(N4097,R1);
not not880(N4098,R2);
not not881(N4099,R3);
not not882(N4109,in2);
not not883(N4110,R2);
not not884(N4111,R3);
not not885(N4121,in2);
not not886(N4122,R3);
not not887(N4133,in2);
not not888(N4134,R1);
not not889(N4135,R5);
not not890(N4145,in1);
not not891(N4146,R2);
not not892(N4157,in0);
not not893(N4158,R2);
not not894(N4169,in2);
not not895(N4170,R0);
not not896(N4171,R5);
not not897(N4181,in0);
not not898(N4182,in1);
not not899(N4183,R0);
not not900(N4184,R5);
not not901(N4193,in2);
not not902(N4194,R1);
not not903(N4195,R4);
not not904(N4205,R1);
not not905(N4206,R2);
not not906(N4207,R5);
not not907(N4217,in2);
not not908(N4218,R2);
not not909(N4219,R3);
not not910(N4229,in1);
not not911(N4230,R5);
not not912(N4241,in0);
not not913(N4242,R4);
not not914(N4253,in0);
not not915(N4254,in2);
not not916(N4255,R2);
not not917(N4256,R5);
not not918(N4265,in2);
not not919(N4266,R0);
not not920(N4267,R1);
not not921(N4268,R5);
not not922(N4277,R2);
not not923(N4278,R4);
not not924(N4279,R5);
not not925(N4289,in1);
not not926(N4290,in2);
not not927(N4291,R0);
not not928(N4301,in1);
not not929(N4302,R0);
not not930(N4303,R1);
not not931(N4313,R3);
not not932(N4314,R4);
not not933(N4325,R3);
not not934(N4326,R4);
not not935(N4337,in2);
not not936(N4338,R0);
not not937(N4339,R5);
not not938(N4349,in1);
not not939(N4350,R0);
not not940(N4351,R4);
not not941(N4361,in1);
not not942(N4362,R3);
not not943(N4363,R4);
not not944(N4373,R0);
not not945(N4374,R1);
not not946(N4375,R3);
not not947(N4385,in1);
not not948(N4386,R0);
not not949(N4387,R1);
not not950(N4397,in0);
not not951(N4398,in2);
not not952(N4399,R0);
not not953(N4409,in1);
not not954(N4410,R0);
not not955(N4411,R2);
not not956(N4421,R1);
not not957(N4422,R4);
not not958(N4423,R5);
not not959(N4433,R0);
not not960(N4434,R2);
not not961(N4435,R5);
not not962(N4445,in2);
not not963(N4446,R0);
not not964(N4447,R1);
not not965(N4457,in1);
not not966(N4458,R4);
not not967(N4469,R0);
not not968(N4470,R5);
not not969(N4481,in2);
not not970(N4482,R3);
not not971(N4483,R4);
not not972(N4493,R2);
not not973(N4494,R5);
not not974(N4505,R0);
not not975(N4506,R2);
not not976(N4507,R4);
not not977(N4517,R0);
not not978(N4518,R2);
not not979(N4529,R0);
not not980(N4530,R1);
not not981(N4531,R2);
not not982(N4541,in0);
not not983(N4542,R0);
not not984(N4543,R4);
not not985(N4553,in2);
not not986(N4554,R2);
not not987(N4565,in0);
not not988(N4566,in1);
not not989(N4567,R0);
not not990(N4577,in1);
not not991(N4578,in2);
not not992(N4579,R0);
not not993(N4589,in2);
not not994(N4590,R0);
not not995(N4591,R2);
not not996(N4601,R1);
not not997(N4602,R3);
not not998(N4612,in1);
not not999(N4613,in2);
not not1000(N4614,R1);
not not1001(N4623,R2);
not not1002(N4624,R5);
not not1003(N4634,R2);
not not1004(N4635,R4);
not not1005(N4645,R1);
not not1006(N4646,R3);
not not1007(N4656,R1);
not not1008(N4657,R4);
not not1009(N4667,in0);
not not1010(N4668,in1);
not not1011(N4669,R2);
not not1012(N4678,in0);
not not1013(N4679,in2);
not not1014(N4689,in1);
not not1015(N4700,in2);
not not1016(N4711,in0);
not not1017(N4712,R4);
not not1018(N4722,in0);
not not1019(N4723,in2);
not not1020(N4724,R5);
not not1021(N4733,in2);
not not1022(N4734,R1);
not not1023(N4735,R2);
not not1024(N4744,R0);
not not1025(N4745,R1);
not not1026(N4746,R2);
not not1027(N4755,R0);
not not1028(N4756,R1);
not not1029(N4757,R2);
not not1030(N4766,in1);
not not1031(N4767,R5);
not not1032(N4777,in1);
not not1033(N4778,in2);
not not1034(N4788,R4);
not not1035(N4789,R5);
not not1036(N4799,in1);
not not1037(N4800,R3);
not not1038(N4810,in1);
not not1039(N4811,R5);
not not1040(N4821,in1);
not not1041(N4822,R1);
not not1042(N4823,R5);
not not1043(N4832,R2);
not not1044(N4833,R5);
not not1045(N4843,in0);
not not1046(N4844,in1);
not not1047(N4854,in1);
not not1048(N4855,R0);
not not1049(N4865,in2);
not not1050(N4866,R4);
not not1051(N4876,R0);
not not1052(N4877,R1);
not not1053(N4878,R5);
not not1054(N4887,in2);
not not1055(N4888,R3);
not not1056(N4898,in1);
not not1057(N4899,R0);
not not1058(N4908,in1);
not not1059(N4909,R4);
not not1060(N4918,R1);
not not1061(N4919,R2);
not not1062(N4928,in0);
not not1063(N4929,R0);
not not1064(N4938,in0);
not not1065(N4939,R3);
not not1066(N4948,R0);
not not1067(N4949,R2);
not not1068(N4958,in2);
not not1069(N4968,R1);
not not1070(N4978,in1);
not not1071(N4988,in0);
not not1072(N4998,in1);
not not1073(N5008,R0);
not not1074(N5018,R0);
not not1075(N5028,R1);
not not1076(N5038,R0);
not not1077(N5058,in2);
not not1078(N5068,R5);
not not1079(N5078,R4);
not not1080(N5087,R5);
not not1081(N5096,R1);
not not1082(N5105,in0);
not not1083(N5114,in0);
not not1084(N5131,in2);
not not1085(N5132,R2);
not not1086(N5133,R3);
not not1087(N5134,R4);
not not1088(N5135,R5);
not not1089(N5136,R6);
not not1090(N5137,R7);
not not1091(N5145,in1);
not not1092(N5146,R0);
not not1093(N5147,R2);
not not1094(N5148,R3);
not not1095(N5149,R4);
not not1096(N5150,R5);
not not1097(N5151,R6);
not not1098(N5159,R0);
not not1099(N5160,R2);
not not1100(N5161,R3);
not not1101(N5162,R4);
not not1102(N5163,R5);
not not1103(N5164,R6);
not not1104(N5165,R7);
not not1105(N5173,in1);
not not1106(N5174,R1);
not not1107(N5175,R2);
not not1108(N5176,R3);
not not1109(N5177,R4);
not not1110(N5178,R5);
not not1111(N5186,in2);
not not1112(N5187,R0);
not not1113(N5188,R3);
not not1114(N5189,R5);
not not1115(N5190,R6);
not not1116(N5191,R7);
not not1117(N5199,in1);
not not1118(N5200,R0);
not not1119(N5201,R1);
not not1120(N5202,R2);
not not1121(N5203,R6);
not not1122(N5204,R7);
not not1123(N5212,R0);
not not1124(N5213,R2);
not not1125(N5214,R3);
not not1126(N5215,R4);
not not1127(N5216,R5);
not not1128(N5217,R6);
not not1129(N5225,in1);
not not1130(N5226,R0);
not not1131(N5227,R2);
not not1132(N5228,R3);
not not1133(N5229,R4);
not not1134(N5230,R6);
not not1135(N5238,in2);
not not1136(N5239,R1);
not not1137(N5240,R3);
not not1138(N5241,R4);
not not1139(N5242,R6);
not not1140(N5250,in1);
not not1141(N5251,R1);
not not1142(N5252,R3);
not not1143(N5253,R4);
not not1144(N5254,R6);
not not1145(N5262,R1);
not not1146(N5263,R4);
not not1147(N5264,R5);
not not1148(N5265,R6);
not not1149(N5266,R7);
not not1150(N5274,in2);
not not1151(N5275,R2);
not not1152(N5276,R5);
not not1153(N5277,R6);
not not1154(N5278,R7);
not not1155(N5286,R0);
not not1156(N5287,R1);
not not1157(N5288,R4);
not not1158(N5289,R5);
not not1159(N5290,R6);
not not1160(N5298,R0);
not not1161(N5299,R1);
not not1162(N5300,R2);
not not1163(N5301,R5);
not not1164(N5302,R7);
not not1165(N5310,in2);
not not1166(N5311,R0);
not not1167(N5312,R2);
not not1168(N5313,R4);
not not1169(N5314,R6);
not not1170(N5322,R0);
not not1171(N5323,R1);
not not1172(N5324,R2);
not not1173(N5325,R6);
not not1174(N5326,R7);
not not1175(N5334,in2);
not not1176(N5335,R3);
not not1177(N5336,R4);
not not1178(N5337,R6);
not not1179(N5345,in1);
not not1180(N5346,R4);
not not1181(N5347,R5);
not not1182(N5348,R6);
not not1183(N5356,in1);
not not1184(N5357,R2);
not not1185(N5358,R5);
not not1186(N5359,R6);
not not1187(N5367,in0);
not not1188(N5368,in2);
not not1189(N5369,R0);
not not1190(N5370,R4);
not not1191(N5378,R1);
not not1192(N5379,R2);
not not1193(N5380,R5);
not not1194(N5381,R7);
not not1195(N5389,R1);
not not1196(N5390,R4);
not not1197(N5391,R5);
not not1198(N5392,R6);
not not1199(N5400,R1);
not not1200(N5401,R5);
not not1201(N5402,R6);
not not1202(N5403,R7);
not not1203(N5411,R1);
not not1204(N5412,R3);
not not1205(N5413,R5);
not not1206(N5414,R7);
not not1207(N5422,R2);
not not1208(N5423,R4);
not not1209(N5424,R5);
not not1210(N5425,R7);
not not1211(N5433,R1);
not not1212(N5434,R2);
not not1213(N5435,R6);
not not1214(N5436,R7);
not not1215(N5444,in0);
not not1216(N5445,R0);
not not1217(N5446,R5);
not not1218(N5447,R7);
not not1219(N5455,in1);
not not1220(N5456,R1);
not not1221(N5457,R4);
not not1222(N5458,R5);
not not1223(N5466,R0);
not not1224(N5467,R1);
not not1225(N5468,R3);
not not1226(N5469,R6);
not not1227(N5477,in2);
not not1228(N5478,R2);
not not1229(N5479,R5);
not not1230(N5480,R6);
not not1231(N5488,R0);
not not1232(N5489,R4);
not not1233(N5490,R6);
not not1234(N5498,R3);
not not1235(N5499,R4);
not not1236(N5500,R5);
not not1237(N5508,R0);
not not1238(N5509,R4);
not not1239(N5510,R7);
not not1240(N5518,R3);
not not1241(N5519,R5);
not not1242(N5520,R7);
not not1243(N5528,in2);
not not1244(N5529,R4);
not not1245(N5530,R6);
not not1246(N5538,in1);
not not1247(N5539,R1);
not not1248(N5540,R3);
not not1249(N5548,in1);
not not1250(N5549,in2);
not not1251(N5550,R6);
not not1252(N5558,in1);
not not1253(N5559,R1);
not not1254(N5560,R7);
not not1255(N5568,in2);
not not1256(N5569,R1);
not not1257(N5570,R6);
not not1258(N5578,R4);
not not1259(N5579,R5);
not not1260(N5580,R6);
not not1261(N5588,in1);
not not1262(N5589,R1);
not not1263(N5590,R6);
not not1264(N5598,in2);
not not1265(N5599,R1);
not not1266(N5600,R3);
not not1267(N5608,R0);
not not1268(N5609,R2);
not not1269(N5617,R4);
not not1270(N5618,R6);
not not1271(N5626,R0);
not not1272(N5627,R4);
not not1273(N5635,R1);
not not1274(N5636,R3);
not not1275(N5644,in2);
not not1276(N5645,R1);
not not1277(N5653,R3);
not not1278(N424,R4);
not not1279(N425,R5);
not not1280(N426,R6);
not not1281(N427,R7);
not not1282(N442,R5);
not not1283(N443,R6);
not not1284(N444,R7);
not not1285(N459,R5);
not not1286(N460,R6);
not not1287(N461,R7);
not not1288(N476,R4);
not not1289(N477,R6);
not not1290(N478,R7);
not not1291(N492,R4);
not not1292(N493,R5);
not not1293(N494,R6);
not not1294(N495,R7);
not not1295(N509,R4);
not not1296(N510,R5);
not not1297(N511,R6);
not not1298(N512,R7);
not not1299(N527,R3);
not not1300(N528,R4);
not not1301(N529,R7);
not not1302(N544,R3);
not not1303(N545,R4);
not not1304(N546,R6);
not not1305(N562,R3);
not not1306(N563,R6);
not not1307(N579,R6);
not not1308(N580,R7);
not not1309(N595,R4);
not not1310(N596,R5);
not not1311(N597,R6);
not not1312(N612,R5);
not not1313(N613,R6);
not not1314(N614,R7);
not not1315(N627,R3);
not not1316(N628,R4);
not not1317(N629,R5);
not not1318(N630,R6);
not not1319(N644,R4);
not not1320(N645,R5);
not not1321(N646,R7);
not not1322(N660,R4);
not not1323(N661,R5);
not not1324(N662,R7);
not not1325(N676,R4);
not not1326(N677,R5);
not not1327(N678,R6);
not not1328(N691,R4);
not not1329(N692,R5);
not not1330(N693,R6);
not not1331(N694,R7);
not not1332(N707,R4);
not not1333(N708,R5);
not not1334(N709,R6);
not not1335(N710,R7);
not not1336(N725,R5);
not not1337(N726,R6);
not not1338(N741,R4);
not not1339(N742,R6);
not not1340(N757,R6);
not not1341(N758,R7);
not not1342(N772,R4);
not not1343(N773,R6);
not not1344(N774,R7);
not not1345(N789,R4);
not not1346(N790,R5);
not not1347(N804,R3);
not not1348(N805,R6);
not not1349(N806,R7);
not not1350(N820,R6);
not not1351(N821,R7);
not not1352(N834,R5);
not not1353(N835,R6);
not not1354(N836,R7);
not not1355(N849,R4);
not not1356(N850,R5);
not not1357(N851,R6);
not not1358(N865,R3);
not not1359(N866,R6);
not not1360(N879,R5);
not not1361(N880,R6);
not not1362(N881,R7);
not not1363(N894,R3);
not not1364(N895,R4);
not not1365(N896,R7);
not not1366(N908,R3);
not not1367(N909,R4);
not not1368(N910,R5);
not not1369(N911,R6);
not not1370(N926,R6);
not not1371(N939,R4);
not not1372(N940,R6);
not not1373(N941,R7);
not not1374(N955,R4);
not not1375(N956,R7);
not not1376(N970,R4);
not not1377(N971,R7);
not not1378(N985,R4);
not not1379(N986,R7);
not not1380(N999,R3);
not not1381(N1000,R4);
not not1382(N1001,R5);
not not1383(N1014,R4);
not not1384(N1015,R6);
not not1385(N1016,R7);
not not1386(N1030,R5);
not not1387(N1031,R6);
not not1388(N1045,R4);
not not1389(N1046,R5);
not not1390(N1059,R3);
not not1391(N1060,R6);
not not1392(N1061,R7);
not not1393(N1074,R3);
not not1394(N1075,R4);
not not1395(N1076,R7);
not not1396(N1090,R5);
not not1397(N1091,R7);
not not1398(N1105,R5);
not not1399(N1106,R6);
not not1400(N1120,R4);
not not1401(N1121,R7);
not not1402(N1135,R6);
not not1403(N1136,R7);
not not1404(N1149,R3);
not not1405(N1150,R5);
not not1406(N1151,R6);
not not1407(N1164,R5);
not not1408(N1165,R6);
not not1409(N1166,R7);
not not1410(N1180,R6);
not not1411(N1181,R7);
not not1412(N1196,R5);
not not1413(N1210,R6);
not not1414(N1211,R7);
not not1415(N1225,R3);
not not1416(N1226,R7);
not not1417(N1239,R3);
not not1418(N1240,R6);
not not1419(N1241,R7);
not not1420(N1255,R4);
not not1421(N1256,R5);
not not1422(N1271,R6);
not not1423(N1285,R4);
not not1424(N1286,R6);
not not1425(N1300,R4);
not not1426(N1301,R7);
not not1427(N1315,R5);
not not1428(N1316,R6);
not not1429(N1330,R5);
not not1430(N1331,R6);
not not1431(N1345,R4);
not not1432(N1346,R7);
not not1433(N1359,R6);
not not1434(N1360,R7);
not not1435(N1371,R3);
not not1436(N1372,R4);
not not1437(N1373,R5);
not not1438(N1374,R7);
not not1439(N1387,R4);
not not1440(N1388,R6);
not not1441(N1402,R4);
not not1442(N1415,R4);
not not1443(N1416,R6);
not not1444(N1429,R4);
not not1445(N1430,R7);
not not1446(N1442,R3);
not not1447(N1443,R4);
not not1448(N1444,R7);
not not1449(N1457,R4);
not not1450(N1458,R7);
not not1451(N1471,R4);
not not1452(N1472,R5);
not not1453(N1485,R4);
not not1454(N1486,R5);
not not1455(N1499,R5);
not not1456(N1500,R6);
not not1457(N1514,R6);
not not1458(N1527,R6);
not not1459(N1528,R7);
not not1460(N1542,R7);
not not1461(N1555,R4);
not not1462(N1556,R7);
not not1463(N1568,R3);
not not1464(N1569,R6);
not not1465(N1570,R7);
not not1466(N1582,R4);
not not1467(N1583,R5);
not not1468(N1584,R6);
not not1469(N1597,R4);
not not1470(N1598,R5);
not not1471(N1612,R7);
not not1472(N1626,R4);
not not1473(N1639,R4);
not not1474(N1640,R5);
not not1475(N1654,R4);
not not1476(N1667,R4);
not not1477(N1668,R7);
not not1478(N1681,R4);
not not1479(N1682,R5);
not not1480(N1696,R4);
not not1481(N1709,R4);
not not1482(N1710,R6);
not not1483(N1723,R4);
not not1484(N1724,R6);
not not1485(N1736,R6);
not not1486(N1737,R7);
not not1487(N1749,R6);
not not1488(N1750,R7);
not not1489(N1762,R6);
not not1490(N1763,R7);
not not1491(N1775,R4);
not not1492(N1776,R6);
not not1493(N1789,R5);
not not1494(N1802,R3);
not not1495(N1813,R4);
not not1496(N1814,R5);
not not1497(N1815,R6);
not not1498(N1827,R5);
not not1499(N1828,R6);
not not1500(N1840,R4);
not not1501(N1841,R7);
not not1502(N1853,R4);
not not1503(N1854,R5);
not not1504(N1866,R4);
not not1505(N1867,R6);
not not1506(N1880,R4);
not not1507(N1904,R3);
not not1508(N1905,R5);
not not1509(N1906,R6);
not not1510(N1918,R6);
not not1511(N1919,R7);
not not1512(N1930,R4);
not not1513(N1931,R5);
not not1514(N1932,R6);
not not1515(N1944,R5);
not not1516(N1945,R6);
not not1517(N1956,R4);
not not1518(N1957,R5);
not not1519(N1958,R7);
not not1520(N1969,R3);
not not1521(N1970,R4);
not not1522(N1971,R7);
not not1523(N1983,R4);
not not1524(N1984,R7);
not not1525(N1996,R5);
not not1526(N1997,R7);
not not1527(N2009,R5);
not not1528(N2010,R7);
not not1529(N2022,R5);
not not1530(N2023,R7);
not not1531(N2035,R5);
not not1532(N2036,R6);
not not1533(N2049,R3);
not not1534(N2075,R6);
not not1535(N2087,R4);
not not1536(N2088,R5);
not not1537(N2100,R4);
not not1538(N2101,R5);
not not1539(N2113,R3);
not not1540(N2114,R6);
not not1541(N2126,R6);
not not1542(N2127,R7);
not not1543(N2139,R3);
not not1544(N2140,R6);
not not1545(N2153,R4);
not not1546(N2166,R6);
not not1547(N2179,R5);
not not1548(N2192,R6);
not not1549(N2217,R4);
not not1550(N2218,R5);
not not1551(N2231,R3);
not not1552(N2243,R4);
not not1553(N2244,R6);
not not1554(N2257,R7);
not not1555(N2283,R4);
not not1556(N2296,R4);
not not1557(N2309,R7);
not not1558(N2322,R7);
not not1559(N2334,R4);
not not1560(N2335,R7);
not not1561(N2346,R6);
not not1562(N2347,R7);
not not1563(N2359,R5);
not not1564(N2371,R5);
not not1565(N2381,R3);
not not1566(N2382,R4);
not not1567(N2383,R7);
not not1568(N2407,R5);
not not1569(N2419,R4);
not not1570(N2431,R5);
not not1571(N2443,R4);
not not1572(N2455,R6);
not not1573(N2467,R5);
not not1574(N2477,R4);
not not1575(N2478,R5);
not not1576(N2479,R7);
not not1577(N2491,R7);
not not1578(N2502,R5);
not not1579(N2503,R6);
not not1580(N2514,R4);
not not1581(N2515,R5);
not not1582(N2527,R6);
not not1583(N2538,R4);
not not1584(N2539,R5);
not not1585(N2551,R6);
not not1586(N2563,R5);
not not1587(N2573,R6);
not not1588(N2574,R7);
not not1589(N2585,R7);
not not1590(N2595,R3);
not not1591(N2596,R7);
not not1592(N2607,R5);
not not1593(N2629,R4);
not not1594(N2640,R6);
not not1595(N2650,R4);
not not1596(N2651,R6);
not not1597(N2673,R6);
not not1598(N2683,R5);
not not1599(N2684,R7);
not not1600(N2695,R7);
not not1601(N2717,R5);
not not1602(N2728,R6);
not not1603(N2739,R4);
not not1604(N2750,R4);
not not1605(N2772,R3);
not not1606(N2782,R4);
not not1607(N2783,R5);
not not1608(N2817,R7);
not not1609(N2832,R6);
not not1610(N2833,R7);
not not1611(N2848,R6);
not not1612(N2849,R7);
not not1613(N2864,R6);
not not1614(N2865,R7);
not not1615(N2880,R6);
not not1616(N2894,R6);
not not1617(N2895,R7);
not not1618(N2909,R5);
not not1619(N2910,R6);
not not1620(N2924,R6);
not not1621(N2925,R7);
not not1622(N2940,R7);
not not1623(N2954,R6);
not not1624(N2955,R7);
not not1625(N2970,R7);
not not1626(N2983,R6);
not not1627(N2984,R7);
not not1628(N2998,R6);
not not1629(N3012,R6);
not not1630(N3025,R5);
not not1631(N3026,R6);
not not1632(N3039,R5);
not not1633(N3040,R6);
not not1634(N3053,R6);
not not1635(N3054,R7);
not not1636(N3068,R6);
not not1637(N3082,R7);
not not1638(N3096,R7);
not not1639(N3110,R7);
not not1640(N3124,R6);
not not1641(N3137,R6);
not not1642(N3138,R7);
not not1643(N3151,R6);
not not1644(N3152,R7);
not not1645(N3165,R6);
not not1646(N3166,R7);
not not1647(N3180,R6);
not not1648(N3207,R6);
not not1649(N3208,R7);
not not1650(N3221,R6);
not not1651(N3222,R7);
not not1652(N3235,R6);
not not1653(N3236,R7);
not not1654(N3249,R6);
not not1655(N3250,R7);
not not1656(N3264,R7);
not not1657(N3278,R5);
not not1658(N3291,R6);
not not1659(N3292,R7);
not not1660(N3306,R7);
not not1661(N3320,R7);
not not1662(N3333,R6);
not not1663(N3334,R7);
not not1664(N3347,R6);
not not1665(N3348,R7);
not not1666(N3362,R6);
not not1667(N3376,R6);
not not1668(N3389,R4);
not not1669(N3390,R6);
not not1670(N3404,R6);
not not1671(N3417,R6);
not not1672(N3418,R7);
not not1673(N3431,R6);
not not1674(N3432,R7);
not not1675(N3445,R6);
not not1676(N3446,R7);
not not1677(N3459,R6);
not not1678(N3460,R7);
not not1679(N3486,R6);
not not1680(N3487,R7);
not not1681(N3499,R6);
not not1682(N3500,R7);
not not1683(N3512,R6);
not not1684(N3513,R7);
not not1685(N3525,R5);
not not1686(N3526,R6);
not not1687(N3539,R6);
not not1688(N3551,R5);
not not1689(N3552,R7);
not not1690(N3564,R6);
not not1691(N3565,R7);
not not1692(N3578,R6);
not not1693(N3591,R6);
not not1694(N3604,R6);
not not1695(N3616,R6);
not not1696(N3617,R7);
not not1697(N3629,R5);
not not1698(N3630,R6);
not not1699(N3642,R6);
not not1700(N3643,R7);
not not1701(N3656,R7);
not not1702(N3668,R6);
not not1703(N3669,R7);
not not1704(N3682,R6);
not not1705(N3707,R6);
not not1706(N3708,R7);
not not1707(N3720,R6);
not not1708(N3721,R7);
not not1709(N3746,R6);
not not1710(N3747,R7);
not not1711(N3759,R6);
not not1712(N3760,R7);
not not1713(N3773,R6);
not not1714(N3799,R7);
not not1715(N3812,R6);
not not1716(N3825,R7);
not not1717(N3837,R5);
not not1718(N3838,R6);
not not1719(N3851,R5);
not not1720(N3864,R7);
not not1721(N3877,R5);
not not1722(N3890,R6);
not not1723(N3903,R6);
not not1724(N3915,R5);
not not1725(N3916,R7);
not not1726(N3929,R7);
not not1727(N3942,R7);
not not1728(N3954,R6);
not not1729(N3955,R7);
not not1730(N3968,R6);
not not1731(N3979,R6);
not not1732(N3980,R7);
not not1733(N3992,R5);
not not1734(N4003,R6);
not not1735(N4004,R7);
not not1736(N4028,R7);
not not1737(N4052,R7);
not not1738(N4075,R6);
not not1739(N4076,R7);
not not1740(N4087,R6);
not not1741(N4088,R7);
not not1742(N4100,R6);
not not1743(N4112,R6);
not not1744(N4123,R6);
not not1745(N4124,R7);
not not1746(N4136,R6);
not not1747(N4147,R6);
not not1748(N4148,R7);
not not1749(N4159,R5);
not not1750(N4160,R6);
not not1751(N4172,R6);
not not1752(N4196,R7);
not not1753(N4208,R7);
not not1754(N4220,R6);
not not1755(N4231,R6);
not not1756(N4232,R7);
not not1757(N4243,R6);
not not1758(N4244,R7);
not not1759(N4280,R7);
not not1760(N4292,R6);
not not1761(N4304,R6);
not not1762(N4315,R6);
not not1763(N4316,R7);
not not1764(N4327,R6);
not not1765(N4328,R7);
not not1766(N4340,R7);
not not1767(N4352,R5);
not not1768(N4364,R6);
not not1769(N4376,R7);
not not1770(N4388,R5);
not not1771(N4400,R7);
not not1772(N4412,R6);
not not1773(N4424,R7);
not not1774(N4436,R6);
not not1775(N4448,R6);
not not1776(N4459,R6);
not not1777(N4460,R7);
not not1778(N4471,R6);
not not1779(N4472,R7);
not not1780(N4484,R7);
not not1781(N4495,R6);
not not1782(N4496,R7);
not not1783(N4508,R6);
not not1784(N4519,R6);
not not1785(N4520,R7);
not not1786(N4532,R6);
not not1787(N4544,R7);
not not1788(N4555,R6);
not not1789(N4556,R7);
not not1790(N4568,R6);
not not1791(N4580,R7);
not not1792(N4592,R6);
not not1793(N4603,R6);
not not1794(N4625,R7);
not not1795(N4636,R7);
not not1796(N4647,R5);
not not1797(N4658,R7);
not not1798(N4680,R7);
not not1799(N4690,R6);
not not1800(N4691,R7);
not not1801(N4701,R5);
not not1802(N4702,R6);
not not1803(N4713,R7);
not not1804(N4768,R6);
not not1805(N4779,R6);
not not1806(N4790,R6);
not not1807(N4801,R7);
not not1808(N4812,R7);
not not1809(N4834,R6);
not not1810(N4845,R7);
not not1811(N4856,R7);
not not1812(N4867,R5);
not not1813(N4889,R7);
not not1814(N4959,R7);
not not1815(N4969,R7);
not not1816(N4979,R7);
not not1817(N4989,R6);
not not1818(N4999,R6);
not not1819(N5009,R6);
not not1820(N5019,R6);
not not1821(N5029,R6);
not not1822(N5039,R7);
not not1823(N5048,R6);
not not1824(N5049,R7);
not not1825(N5059,R6);
not not1826(N5069,R6);
not not1827(N5123,R7);
not not1828(N5854,in0);
not not1829(N5855,R0);
not not1830(N5856,R1);
not not1831(N5870,in0);
not not1832(N5871,in1);
not not1833(N5884,in0);
not not1834(N5885,in1);
not not1835(N5886,R0);
not not1836(N5887,R2);
not not1837(N5901,in0);
not not1838(N5902,R0);
not not1839(N5903,R1);
not not1840(N5904,R2);
not not1841(N5905,R3);
not not1842(N5918,in0);
not not1843(N5919,R0);
not not1844(N5920,R2);
not not1845(N5921,R3);
not not1846(N5935,in0);
not not1847(N5936,in1);
not not1848(N5937,R0);
not not1849(N5938,R1);
not not1850(N5952,in0);
not not1851(N5953,in2);
not not1852(N5954,R0);
not not1853(N5955,R1);
not not1854(N5969,in0);
not not1855(N5970,in1);
not not1856(N5971,R0);
not not1857(N5972,R1);
not not1858(N5973,R3);
not not1859(N5986,in0);
not not1860(N5987,in2);
not not1861(N5988,R0);
not not1862(N5989,R1);
not not1863(N5990,R3);
not not1864(N6003,in0);
not not1865(N6004,in1);
not not1866(N6005,in2);
not not1867(N6006,R1);
not not1868(N6007,R2);
not not1869(N6020,in0);
not not1870(N6021,in1);
not not1871(N6022,in2);
not not1872(N6023,R0);
not not1873(N6024,R2);
not not1874(N6037,in0);
not not1875(N6038,in1);
not not1876(N6039,in2);
not not1877(N6040,R0);
not not1878(N6041,R1);
not not1879(N6054,in0);
not not1880(N6055,in1);
not not1881(N6056,in2);
not not1882(N6057,R0);
not not1883(N6058,R1);
not not1884(N6071,in0);
not not1885(N6072,R0);
not not1886(N6073,R1);
not not1887(N6074,R2);
not not1888(N6087,in0);
not not1889(N6088,in2);
not not1890(N6089,R2);
not not1891(N6090,R3);
not not1892(N6103,in0);
not not1893(N6104,in1);
not not1894(N6105,R2);
not not1895(N6106,R3);
not not1896(N6119,in0);
not not1897(N6120,in1);
not not1898(N6121,R0);
not not1899(N6135,in0);
not not1900(N6136,in1);
not not1901(N6137,R0);
not not1902(N6138,R1);
not not1903(N6151,in0);
not not1904(N6152,in2);
not not1905(N6153,R0);
not not1906(N6154,R1);
not not1907(N6167,in0);
not not1908(N6168,in1);
not not1909(N6169,in2);
not not1910(N6170,R2);
not not1911(N6183,in0);
not not1912(N6184,in1);
not not1913(N6185,R1);
not not1914(N6186,R2);
not not1915(N6199,in0);
not not1916(N6200,in1);
not not1917(N6201,in2);
not not1918(N6202,R1);
not not1919(N6203,R3);
not not1920(N6215,in0);
not not1921(N6216,in1);
not not1922(N6217,R0);
not not1923(N6218,R2);
not not1924(N6231,in0);
not not1925(N6232,in1);
not not1926(N6233,R0);
not not1927(N6234,R1);
not not1928(N6235,R2);
not not1929(N6247,in0);
not not1930(N6248,in1);
not not1931(N6249,in2);
not not1932(N6250,R2);
not not1933(N6263,in0);
not not1934(N6264,in2);
not not1935(N6265,R0);
not not1936(N6266,R2);
not not1937(N6279,in0);
not not1938(N6280,in1);
not not1939(N6281,in2);
not not1940(N6282,R0);
not not1941(N6283,R2);
not not1942(N6295,in0);
not not1943(N6296,in1);
not not1944(N6297,R0);
not not1945(N6298,R1);
not not1946(N6310,in0);
not not1947(N6311,in1);
not not1948(N6312,R0);
not not1949(N6313,R1);
not not1950(N6314,R3);
not not1951(N6325,in0);
not not1952(N6326,R2);
not not1953(N6327,R3);
not not1954(N6340,in0);
not not1955(N6341,in1);
not not1956(N6342,in2);
not not1957(N6343,R3);
not not1958(N6355,in0);
not not1959(N6356,in1);
not not1960(N6357,R1);
not not1961(N6370,in0);
not not1962(N6371,R1);
not not1963(N6372,R3);
not not1964(N6385,in0);
not not1965(N6386,in1);
not not1966(N6387,in2);
not not1967(N6400,in0);
not not1968(N6401,R0);
not not1969(N6402,R2);
not not1970(N6415,in0);
not not1971(N6416,in2);
not not1972(N6417,R1);
not not1973(N6430,in0);
not not1974(N6431,in1);
not not1975(N6432,in2);
not not1976(N6433,R1);
not not1977(N6434,R2);
not not1978(N6445,in0);
not not1979(N6446,in1);
not not1980(N6447,R1);
not not1981(N6448,R3);
not not1982(N6460,in0);
not not1983(N6461,in2);
not not1984(N6462,R0);
not not1985(N6463,R1);
not not1986(N6475,in0);
not not1987(N6476,in2);
not not1988(N6477,R0);
not not1989(N6478,R3);
not not1990(N6490,in0);
not not1991(N6491,in1);
not not1992(N6492,in2);
not not1993(N6493,R0);
not not1994(N6505,in0);
not not1995(N6506,in2);
not not1996(N6507,R2);
not not1997(N6520,in0);
not not1998(N6521,in2);
not not1999(N6522,R1);
not not2000(N6535,in0);
not not2001(N6536,in1);
not not2002(N6537,R1);
not not2003(N6550,in0);
not not2004(N6551,R0);
not not2005(N6552,R2);
not not2006(N6553,R3);
not not2007(N6565,in0);
not not2008(N6566,R0);
not not2009(N6567,R3);
not not2010(N6580,in0);
not not2011(N6581,in1);
not not2012(N6582,in2);
not not2013(N6583,R1);
not not2014(N6595,in0);
not not2015(N6596,in2);
not not2016(N6597,R0);
not not2017(N6598,R3);
not not2018(N6610,in0);
not not2019(N6611,R0);
not not2020(N6612,R2);
not not2021(N6613,R3);
not not2022(N6625,in0);
not not2023(N6626,in1);
not not2024(N6627,R1);
not not2025(N6628,R2);
not not2026(N6629,R3);
not not2027(N6640,in0);
not not2028(N6641,in1);
not not2029(N6642,in2);
not not2030(N6643,R1);
not not2031(N6655,in0);
not not2032(N6656,R0);
not not2033(N6657,R1);
not not2034(N6658,R2);
not not2035(N6670,in0);
not not2036(N6671,R1);
not not2037(N6672,R3);
not not2038(N6685,in0);
not not2039(N6686,in1);
not not2040(N6687,R1);
not not2041(N6700,in0);
not not2042(N6701,in1);
not not2043(N6702,R0);
not not2044(N6703,R1);
not not2045(N6715,in0);
not not2046(N6716,in2);
not not2047(N6717,R0);
not not2048(N6718,R1);
not not2049(N6730,in0);
not not2050(N6731,in1);
not not2051(N6732,in2);
not not2052(N6733,R0);
not not2053(N6745,in0);
not not2054(N6746,in1);
not not2055(N6747,R1);
not not2056(N6748,R2);
not not2057(N6760,in0);
not not2058(N6761,in1);
not not2059(N6762,R1);
not not2060(N6763,R2);
not not2061(N6775,in0);
not not2062(N6776,in1);
not not2063(N6777,R1);
not not2064(N6778,R2);
not not2065(N6790,in0);
not not2066(N6791,in2);
not not2067(N6792,R2);
not not2068(N6805,in0);
not not2069(N6806,in1);
not not2070(N6807,in2);
not not2071(N6820,in0);
not not2072(N6821,in2);
not not2073(N6822,R1);
not not2074(N6823,R3);
not not2075(N6835,in0);
not not2076(N6836,in1);
not not2077(N6837,in2);
not not2078(N6838,R0);
not not2079(N6839,R1);
not not2080(N6850,in0);
not not2081(N6851,in2);
not not2082(N6852,R1);
not not2083(N6853,R2);
not not2084(N6865,in0);
not not2085(N6866,R0);
not not2086(N6867,R1);
not not2087(N6868,R2);
not not2088(N6880,in0);
not not2089(N6881,in1);
not not2090(N6882,R0);
not not2091(N6883,R1);
not not2092(N6895,in0);
not not2093(N6896,in2);
not not2094(N6897,R0);
not not2095(N6898,R1);
not not2096(N6910,in0);
not not2097(N6911,in1);
not not2098(N6912,in2);
not not2099(N6913,R0);
not not2100(N6925,in0);
not not2101(N6926,in1);
not not2102(N6940,in0);
not not2103(N6941,in2);
not not2104(N6942,R2);
not not2105(N6955,in0);
not not2106(N6956,in2);
not not2107(N6957,R0);
not not2108(N6958,R1);
not not2109(N6969,in0);
not not2110(N6983,in0);
not not2111(N6984,R0);
not not2112(N6997,in0);
not not2113(N6998,R0);
not not2114(N7011,in0);
not not2115(N7012,R0);
not not2116(N7025,in0);
not not2117(N7026,in1);
not not2118(N7027,in2);
not not2119(N7028,R1);
not not2120(N7029,R3);
not not2121(N7039,in0);
not not2122(N7040,R1);
not not2123(N7041,R2);
not not2124(N7053,in0);
not not2125(N7054,in1);
not not2126(N7055,in2);
not not2127(N7067,in0);
not not2128(N7068,in1);
not not2129(N7069,in2);
not not2130(N7070,R1);
not not2131(N7081,in0);
not not2132(N7082,R1);
not not2133(N7083,R2);
not not2134(N7095,in0);
not not2135(N7096,in2);
not not2136(N7097,R1);
not not2137(N7109,in0);
not not2138(N7110,in2);
not not2139(N7123,in0);
not not2140(N7124,in1);
not not2141(N7137,in0);
not not2142(N7138,R1);
not not2143(N7151,in0);
not not2144(N7152,in1);
not not2145(N7153,in2);
not not2146(N7154,R2);
not not2147(N7165,in0);
not not2148(N7166,in2);
not not2149(N7167,R1);
not not2150(N7168,R2);
not not2151(N7179,in0);
not not2152(N7180,R3);
not not2153(N7193,in0);
not not2154(N7194,in1);
not not2155(N7195,R2);
not not2156(N7207,in0);
not not2157(N7208,in1);
not not2158(N7209,in2);
not not2159(N7210,R0);
not not2160(N7211,R1);
not not2161(N7221,in0);
not not2162(N7222,R0);
not not2163(N7223,R2);
not not2164(N7235,in0);
not not2165(N7236,in1);
not not2166(N7237,in2);
not not2167(N7249,in0);
not not2168(N7250,R2);
not not2169(N7263,in0);
not not2170(N7264,R1);
not not2171(N7277,in0);
not not2172(N7278,in2);
not not2173(N7290,in0);
not not2174(N7291,in2);
not not2175(N7292,R0);
not not2176(N7303,in0);
not not2177(N7304,in2);
not not2178(N7305,R0);
not not2179(N7306,R2);
not not2180(N7316,in0);
not not2181(N7317,R0);
not not2182(N7318,R1);
not not2183(N7329,in0);
not not2184(N7330,R3);
not not2185(N7342,in0);
not not2186(N7343,R0);
not not2187(N7355,in0);
not not2188(N7356,R2);
not not2189(N7368,in0);
not not2190(N7369,in1);
not not2191(N7370,R0);
not not2192(N7381,in0);
not not2193(N7382,in2);
not not2194(N7383,R1);
not not2195(N7394,in0);
not not2196(N7395,in1);
not not2197(N7407,in0);
not not2198(N7408,in2);
not not2199(N7420,in0);
not not2200(N7421,in1);
not not2201(N7433,in0);
not not2202(N7434,R0);
not not2203(N7435,R1);
not not2204(N7436,R2);
not not2205(N7446,in0);
not not2206(N7447,R1);
not not2207(N7448,R2);
not not2208(N7459,in0);
not not2209(N7460,in1);
not not2210(N7461,in2);
not not2211(N7472,in0);
not not2212(N7473,in2);
not not2213(N7474,R1);
not not2214(N7485,in0);
not not2215(N7486,R2);
not not2216(N7498,in0);
not not2217(N7499,R2);
not not2218(N7511,in0);
not not2219(N7512,in2);
not not2220(N7513,R0);
not not2221(N7524,in0);
not not2222(N7525,R3);
not not2223(N7537,in0);
not not2224(N7538,R0);
not not2225(N7539,R1);
not not2226(N7540,R3);
not not2227(N7550,in0);
not not2228(N7551,R0);
not not2229(N7552,R1);
not not2230(N7553,R3);
not not2231(N7563,in0);
not not2232(N7576,in0);
not not2233(N7577,in1);
not not2234(N7578,R1);
not not2235(N7589,in0);
not not2236(N7590,in1);
not not2237(N7591,R0);
not not2238(N7602,in0);
not not2239(N7603,in2);
not not2240(N7615,in0);
not not2241(N7628,in0);
not not2242(N7629,in1);
not not2243(N7630,R3);
not not2244(N7641,in0);
not not2245(N7642,in2);
not not2246(N7643,R0);
not not2247(N7644,R2);
not not2248(N7654,in0);
not not2249(N7655,R1);
not not2250(N7656,R3);
not not2251(N7667,in0);
not not2252(N7668,in2);
not not2253(N7669,R3);
not not2254(N7680,in0);
not not2255(N7681,in1);
not not2256(N7682,R0);
not not2257(N7693,in0);
not not2258(N7694,in2);
not not2259(N7695,R0);
not not2260(N7706,in0);
not not2261(N7707,R0);
not not2262(N7719,in0);
not not2263(N7720,in1);
not not2264(N7721,R1);
not not2265(N7732,in0);
not not2266(N7733,in1);
not not2267(N7734,R1);
not not2268(N7745,in0);
not not2269(N7746,in1);
not not2270(N7747,R0);
not not2271(N7758,in0);
not not2272(N7759,R0);
not not2273(N7760,R1);
not not2274(N7771,in0);
not not2275(N7772,R1);
not not2276(N7784,in0);
not not2277(N7785,R1);
not not2278(N7786,R3);
not not2279(N7797,in0);
not not2280(N7798,in1);
not not2281(N7810,in0);
not not2282(N7811,R0);
not not2283(N7812,R2);
not not2284(N7823,in0);
not not2285(N7824,in1);
not not2286(N7825,R0);
not not2287(N7835,in0);
not not2288(N7847,in0);
not not2289(N7848,R1);
not not2290(N7859,in0);
not not2291(N7860,R3);
not not2292(N7871,in0);
not not2293(N7872,in2);
not not2294(N7883,in0);
not not2295(N7895,in0);
not not2296(N7896,R3);
not not2297(N7907,in0);
not not2298(N7908,in1);
not not2299(N7919,in0);
not not2300(N7920,in2);
not not2301(N7931,in0);
not not2302(N7943,in0);
not not2303(N7944,in2);
not not2304(N7955,in0);
not not2305(N7956,in2);
not not2306(N7967,in0);
not not2307(N7968,R3);
not not2308(N7979,in0);
not not2309(N7980,R1);
not not2310(N7990,in0);
not not2311(N7991,R1);
not not2312(N8001,in0);
not not2313(N8002,R1);
not not2314(N8012,in0);
not not2315(N8013,R2);
not not2316(N8023,in0);
not not2317(N8024,R0);
not not2318(N8034,in0);
not not2319(N8035,R0);
not not2320(N8045,in0);
not not2321(N8046,R1);
not not2322(N8056,in0);
not not2323(N8057,R2);
not not2324(N8067,in0);
not not2325(N8076,in0);
not not2326(N8077,in2);
not not2327(N8078,R1);
not not2328(N8079,R2);
not not2329(N8080,R4);
not not2330(N8081,R5);
not not2331(N8092,in0);
not not2332(N8093,R0);
not not2333(N8094,R1);
not not2334(N8095,R2);
not not2335(N8096,R4);
not not2336(N8097,R5);
not not2337(N8108,in0);
not not2338(N8109,R0);
not not2339(N8110,R1);
not not2340(N8111,R2);
not not2341(N8112,R3);
not not2342(N8113,R4);
not not2343(N8114,R5);
not not2344(N8124,in0);
not not2345(N8125,in1);
not not2346(N8126,R0);
not not2347(N8127,R1);
not not2348(N8128,R2);
not not2349(N8129,R3);
not not2350(N8130,R4);
not not2351(N8140,in0);
not not2352(N8141,in1);
not not2353(N8142,in2);
not not2354(N8143,R3);
not not2355(N8144,R4);
not not2356(N8155,in0);
not not2357(N8156,in1);
not not2358(N8157,in2);
not not2359(N8158,R1);
not not2360(N8159,R2);
not not2361(N8170,in0);
not not2362(N8171,R1);
not not2363(N8172,R2);
not not2364(N8173,R4);
not not2365(N8174,R5);
not not2366(N8185,in0);
not not2367(N8186,R0);
not not2368(N8187,R1);
not not2369(N8188,R4);
not not2370(N8189,R5);
not not2371(N8200,in0);
not not2372(N8201,in2);
not not2373(N8202,R0);
not not2374(N8203,R4);
not not2375(N8214,in0);
not not2376(N8215,in1);
not not2377(N8216,R0);
not not2378(N8217,R3);
not not2379(N8228,in0);
not not2380(N8229,in1);
not not2381(N8230,in2);
not not2382(N8231,R1);
not not2383(N8232,R3);
not not2384(N8242,in0);
not not2385(N8243,in1);
not not2386(N8244,in2);
not not2387(N8245,R0);
not not2388(N8246,R1);
not not2389(N8256,in0);
not not2390(N8257,in2);
not not2391(N8258,R0);
not not2392(N8259,R4);
not not2393(N8270,in0);
not not2394(N8271,R1);
not not2395(N8272,R2);
not not2396(N8283,in0);
not not2397(N8284,in2);
not not2398(N8285,R1);
not not2399(N8286,R2);
not not2400(N8287,R4);
not not2401(N8296,in0);
not not2402(N8297,R1);
not not2403(N8298,R3);
not not2404(N8309,in0);
not not2405(N8310,in2);
not not2406(N8311,R1);
not not2407(N8312,R5);
not not2408(N8322,in0);
not not2409(N8323,R1);
not not2410(N8324,R5);
not not2411(N8335,in0);
not not2412(N8336,in2);
not not2413(N8337,R0);
not not2414(N8338,R1);
not not2415(N8339,R5);
not not2416(N8348,in0);
not not2417(N8349,R3);
not not2418(N8350,R4);
not not2419(N8361,in0);
not not2420(N8362,in1);
not not2421(N8363,R0);
not not2422(N8373,in0);
not not2423(N8374,in1);
not not2424(N8375,R3);
not not2425(N8385,in0);
not not2426(N8386,R1);
not not2427(N8387,R2);
not not2428(N8388,R5);
not not2429(N8397,in0);
not not2430(N8398,R0);
not not2431(N8399,R1);
not not2432(N8400,R2);
not not2433(N8409,in0);
not not2434(N8410,in2);
not not2435(N8411,R1);
not not2436(N8412,R4);
not not2437(N8421,in0);
not not2438(N8422,R1);
not not2439(N8423,R2);
not not2440(N5857,R3);
not not2441(N5858,R4);
not not2442(N5859,R5);
not not2443(N5872,R3);
not not2444(N5873,R5);
not not2445(N5874,R7);
not not2446(N5888,R4);
not not2447(N5889,R5);
not not2448(N5890,R6);
not not2449(N5891,R7);
not not2450(N5906,R5);
not not2451(N5907,R6);
not not2452(N5908,R7);
not not2453(N5922,R4);
not not2454(N5923,R5);
not not2455(N5924,R6);
not not2456(N5925,R7);
not not2457(N5939,R3);
not not2458(N5940,R4);
not not2459(N5941,R5);
not not2460(N5942,R6);
not not2461(N5956,R3);
not not2462(N5957,R4);
not not2463(N5958,R5);
not not2464(N5959,R6);
not not2465(N5974,R4);
not not2466(N5975,R6);
not not2467(N5976,R7);
not not2468(N5991,R4);
not not2469(N5992,R6);
not not2470(N5993,R7);
not not2471(N6008,R3);
not not2472(N6009,R4);
not not2473(N6010,R6);
not not2474(N6025,R4);
not not2475(N6026,R6);
not not2476(N6027,R7);
not not2477(N6042,R4);
not not2478(N6043,R5);
not not2479(N6044,R6);
not not2480(N6059,R5);
not not2481(N6060,R6);
not not2482(N6061,R7);
not not2483(N6075,R4);
not not2484(N6076,R5);
not not2485(N6077,R7);
not not2486(N6091,R5);
not not2487(N6092,R6);
not not2488(N6093,R7);
not not2489(N6107,R5);
not not2490(N6108,R6);
not not2491(N6109,R7);
not not2492(N6122,R4);
not not2493(N6123,R5);
not not2494(N6124,R6);
not not2495(N6125,R7);
not not2496(N6139,R4);
not not2497(N6140,R5);
not not2498(N6141,R7);
not not2499(N6155,R4);
not not2500(N6156,R5);
not not2501(N6157,R7);
not not2502(N6171,R5);
not not2503(N6172,R6);
not not2504(N6173,R7);
not not2505(N6187,R3);
not not2506(N6188,R4);
not not2507(N6189,R5);
not not2508(N6204,R5);
not not2509(N6205,R7);
not not2510(N6219,R4);
not not2511(N6220,R5);
not not2512(N6221,R7);
not not2513(N6236,R4);
not not2514(N6237,R5);
not not2515(N6251,R5);
not not2516(N6252,R6);
not not2517(N6253,R7);
not not2518(N6267,R5);
not not2519(N6268,R6);
not not2520(N6269,R7);
not not2521(N6284,R5);
not not2522(N6285,R6);
not not2523(N6299,R4);
not not2524(N6300,R6);
not not2525(N6315,R6);
not not2526(N6328,R4);
not not2527(N6329,R5);
not not2528(N6330,R6);
not not2529(N6344,R6);
not not2530(N6345,R7);
not not2531(N6358,R5);
not not2532(N6359,R6);
not not2533(N6360,R7);
not not2534(N6373,R4);
not not2535(N6374,R5);
not not2536(N6375,R6);
not not2537(N6388,R3);
not not2538(N6389,R4);
not not2539(N6390,R7);
not not2540(N6403,R4);
not not2541(N6404,R6);
not not2542(N6405,R7);
not not2543(N6418,R4);
not not2544(N6419,R5);
not not2545(N6420,R6);
not not2546(N6435,R4);
not not2547(N6449,R4);
not not2548(N6450,R7);
not not2549(N6464,R3);
not not2550(N6465,R7);
not not2551(N6479,R4);
not not2552(N6480,R6);
not not2553(N6494,R4);
not not2554(N6495,R7);
not not2555(N6508,R4);
not not2556(N6509,R5);
not not2557(N6510,R6);
not not2558(N6523,R4);
not not2559(N6524,R5);
not not2560(N6525,R6);
not not2561(N6538,R3);
not not2562(N6539,R4);
not not2563(N6540,R5);
not not2564(N6554,R4);
not not2565(N6555,R6);
not not2566(N6568,R4);
not not2567(N6569,R6);
not not2568(N6570,R7);
not not2569(N6584,R3);
not not2570(N6585,R6);
not not2571(N6599,R5);
not not2572(N6600,R6);
not not2573(N6614,R4);
not not2574(N6615,R6);
not not2575(N6630,R4);
not not2576(N6644,R4);
not not2577(N6645,R7);
not not2578(N6659,R4);
not not2579(N6660,R5);
not not2580(N6673,R4);
not not2581(N6674,R6);
not not2582(N6675,R7);
not not2583(N6688,R4);
not not2584(N6689,R5);
not not2585(N6690,R6);
not not2586(N6704,R6);
not not2587(N6705,R7);
not not2588(N6719,R5);
not not2589(N6720,R6);
not not2590(N6734,R4);
not not2591(N6735,R7);
not not2592(N6749,R6);
not not2593(N6750,R7);
not not2594(N6764,R5);
not not2595(N6765,R7);
not not2596(N6779,R3);
not not2597(N6780,R6);
not not2598(N6793,R3);
not not2599(N6794,R6);
not not2600(N6795,R7);
not not2601(N6808,R4);
not not2602(N6809,R5);
not not2603(N6810,R6);
not not2604(N6824,R5);
not not2605(N6825,R7);
not not2606(N6840,R6);
not not2607(N6854,R5);
not not2608(N6855,R7);
not not2609(N6869,R6);
not not2610(N6870,R7);
not not2611(N6884,R3);
not not2612(N6885,R5);
not not2613(N6899,R4);
not not2614(N6900,R7);
not not2615(N6914,R3);
not not2616(N6915,R5);
not not2617(N6927,R4);
not not2618(N6928,R5);
not not2619(N6929,R6);
not not2620(N6930,R7);
not not2621(N6943,R4);
not not2622(N6944,R6);
not not2623(N6945,R7);
not not2624(N6959,R6);
not not2625(N6970,R3);
not not2626(N6971,R4);
not not2627(N6972,R5);
not not2628(N6973,R7);
not not2629(N6985,R4);
not not2630(N6986,R5);
not not2631(N6987,R7);
not not2632(N6999,R4);
not not2633(N7000,R5);
not not2634(N7001,R7);
not not2635(N7013,R4);
not not2636(N7014,R5);
not not2637(N7015,R7);
not not2638(N7042,R3);
not not2639(N7043,R6);
not not2640(N7056,R5);
not not2641(N7057,R7);
not not2642(N7071,R7);
not not2643(N7084,R3);
not not2644(N7085,R4);
not not2645(N7098,R5);
not not2646(N7099,R7);
not not2647(N7111,R3);
not not2648(N7112,R6);
not not2649(N7113,R7);
not not2650(N7125,R3);
not not2651(N7126,R6);
not not2652(N7127,R7);
not not2653(N7139,R3);
not not2654(N7140,R5);
not not2655(N7141,R7);
not not2656(N7155,R4);
not not2657(N7169,R4);
not not2658(N7181,R4);
not not2659(N7182,R5);
not not2660(N7183,R7);
not not2661(N7196,R4);
not not2662(N7197,R5);
not not2663(N7224,R6);
not not2664(N7225,R7);
not not2665(N7238,R4);
not not2666(N7239,R7);
not not2667(N7251,R3);
not not2668(N7252,R4);
not not2669(N7253,R6);
not not2670(N7265,R3);
not not2671(N7266,R5);
not not2672(N7267,R6);
not not2673(N7279,R6);
not not2674(N7280,R7);
not not2675(N7293,R7);
not not2676(N7319,R6);
not not2677(N7331,R4);
not not2678(N7332,R7);
not not2679(N7344,R3);
not not2680(N7345,R6);
not not2681(N7357,R5);
not not2682(N7358,R7);
not not2683(N7371,R5);
not not2684(N7384,R3);
not not2685(N7396,R4);
not not2686(N7397,R6);
not not2687(N7409,R4);
not not2688(N7410,R6);
not not2689(N7422,R4);
not not2690(N7423,R6);
not not2691(N7449,R5);
not not2692(N7462,R3);
not not2693(N7475,R4);
not not2694(N7487,R5);
not not2695(N7488,R7);
not not2696(N7500,R5);
not not2697(N7501,R7);
not not2698(N7514,R4);
not not2699(N7526,R4);
not not2700(N7527,R7);
not not2701(N7564,R4);
not not2702(N7565,R5);
not not2703(N7566,R6);
not not2704(N7579,R6);
not not2705(N7592,R6);
not not2706(N7604,R6);
not not2707(N7605,R7);
not not2708(N7616,R5);
not not2709(N7617,R6);
not not2710(N7618,R7);
not not2711(N7631,R6);
not not2712(N7657,R7);
not not2713(N7670,R4);
not not2714(N7683,R6);
not not2715(N7696,R3);
not not2716(N7708,R5);
not not2717(N7709,R6);
not not2718(N7722,R6);
not not2719(N7735,R4);
not not2720(N7748,R7);
not not2721(N7761,R6);
not not2722(N7773,R4);
not not2723(N7774,R7);
not not2724(N7787,R7);
not not2725(N7799,R4);
not not2726(N7800,R6);
not not2727(N7813,R4);
not not2728(N7836,R4);
not not2729(N7837,R5);
not not2730(N7849,R5);
not not2731(N7861,R7);
not not2732(N7873,R4);
not not2733(N7884,R5);
not not2734(N7885,R7);
not not2735(N7897,R5);
not not2736(N7909,R4);
not not2737(N7921,R7);
not not2738(N7932,R5);
not not2739(N7933,R6);
not not2740(N7945,R6);
not not2741(N7957,R5);
not not2742(N7969,R6);
not not2743(N8082,R6);
not not2744(N8083,R7);
not not2745(N8098,R6);
not not2746(N8099,R7);
not not2747(N8115,R6);
not not2748(N8131,R6);
not not2749(N8145,R5);
not not2750(N8146,R6);
not not2751(N8160,R6);
not not2752(N8161,R7);
not not2753(N8175,R6);
not not2754(N8176,R7);
not not2755(N8190,R6);
not not2756(N8191,R7);
not not2757(N8204,R6);
not not2758(N8205,R7);
not not2759(N8218,R6);
not not2760(N8219,R7);
not not2761(N8233,R6);
not not2762(N8247,R5);
not not2763(N8260,R5);
not not2764(N8261,R6);
not not2765(N8273,R6);
not not2766(N8274,R7);
not not2767(N8299,R6);
not not2768(N8300,R7);
not not2769(N8313,R6);
not not2770(N8325,R6);
not not2771(N8326,R7);
not not2772(N8351,R6);
not not2773(N8352,R7);
not not2774(N8364,R7);
not not2775(N8376,R6);
not not2776(N8424,R7);
not not2777(N8894,in0);
not not2778(N8895,in2);
not not2779(N8896,R0);
not not2780(N8897,R1);
not not2781(N8898,R2);
not not2782(N8899,R3);
not not2783(N8912,in0);
not not2784(N8913,in2);
not not2785(N8914,R1);
not not2786(N8915,R2);
not not2787(N8929,in0);
not not2788(N8930,in1);
not not2789(N8931,in2);
not not2790(N8932,R0);
not not2791(N8933,R1);
not not2792(N8946,in0);
not not2793(N8947,in1);
not not2794(N8948,R1);
not not2795(N8949,R2);
not not2796(N8950,R3);
not not2797(N8963,in0);
not not2798(N8964,in1);
not not2799(N8965,in2);
not not2800(N8966,R0);
not not2801(N8967,R1);
not not2802(N8968,R3);
not not2803(N8980,in0);
not not2804(N8981,in1);
not not2805(N8982,in2);
not not2806(N8983,R1);
not not2807(N8984,R3);
not not2808(N8997,in1);
not not2809(N8998,R0);
not not2810(N8999,R2);
not not2811(N9013,R0);
not not2812(N9014,R2);
not not2813(N9015,R3);
not not2814(N9029,in0);
not not2815(N9030,in1);
not not2816(N9031,R0);
not not2817(N9032,R1);
not not2818(N9033,R3);
not not2819(N9045,in2);
not not2820(N9046,R1);
not not2821(N9047,R2);
not not2822(N9048,R3);
not not2823(N9061,in1);
not not2824(N9062,R1);
not not2825(N9063,R2);
not not2826(N9064,R3);
not not2827(N9077,R0);
not not2828(N9078,R1);
not not2829(N9079,R3);
not not2830(N9093,R0);
not not2831(N9094,R1);
not not2832(N9095,R2);
not not2833(N9096,R3);
not not2834(N9109,in1);
not not2835(N9110,R2);
not not2836(N9111,R3);
not not2837(N9125,in0);
not not2838(N9126,R2);
not not2839(N9127,R3);
not not2840(N9141,in0);
not not2841(N9142,in1);
not not2842(N9143,R0);
not not2843(N9144,R1);
not not2844(N9157,in0);
not not2845(N9158,R1);
not not2846(N9159,R2);
not not2847(N9160,R3);
not not2848(N9173,in0);
not not2849(N9174,in1);
not not2850(N9175,in2);
not not2851(N9176,R1);
not not2852(N9177,R3);
not not2853(N9189,in0);
not not2854(N9190,in1);
not not2855(N9191,R0);
not not2856(N9192,R1);
not not2857(N9193,R2);
not not2858(N9205,in1);
not not2859(N9206,in2);
not not2860(N9207,R2);
not not2861(N9208,R3);
not not2862(N9221,in0);
not not2863(N9222,in1);
not not2864(N9223,in2);
not not2865(N9224,R0);
not not2866(N9225,R1);
not not2867(N9237,in0);
not not2868(N9238,in1);
not not2869(N9239,in2);
not not2870(N9240,R1);
not not2871(N9252,in0);
not not2872(N9253,in1);
not not2873(N9254,in2);
not not2874(N9255,R1);
not not2875(N9267,in2);
not not2876(N9268,R0);
not not2877(N9269,R2);
not not2878(N9282,in0);
not not2879(N9283,in2);
not not2880(N9284,R0);
not not2881(N9285,R1);
not not2882(N9286,R2);
not not2883(N9297,in1);
not not2884(N9298,R0);
not not2885(N9299,R1);
not not2886(N9300,R3);
not not2887(N9312,in0);
not not2888(N9313,in1);
not not2889(N9314,in2);
not not2890(N9315,R0);
not not2891(N9327,in1);
not not2892(N9328,R2);
not not2893(N9329,R3);
not not2894(N9342,in0);
not not2895(N9343,R0);
not not2896(N9344,R1);
not not2897(N9357,in0);
not not2898(N9358,in2);
not not2899(N9359,R1);
not not2900(N9372,in0);
not not2901(N9373,R1);
not not2902(N9387,in2);
not not2903(N9388,R0);
not not2904(N9389,R2);
not not2905(N9390,R3);
not not2906(N9402,in0);
not not2907(N9403,in1);
not not2908(N9404,in2);
not not2909(N9405,R3);
not not2910(N9417,in0);
not not2911(N9418,in1);
not not2912(N9419,in2);
not not2913(N9420,R1);
not not2914(N9421,R2);
not not2915(N9432,in0);
not not2916(N9433,in1);
not not2917(N9434,in2);
not not2918(N9435,R3);
not not2919(N9447,in1);
not not2920(N9448,R0);
not not2921(N9449,R1);
not not2922(N9450,R2);
not not2923(N9462,in2);
not not2924(N9463,R0);
not not2925(N9464,R1);
not not2926(N9465,R2);
not not2927(N9477,in2);
not not2928(N9478,R1);
not not2929(N9479,R3);
not not2930(N9492,in1);
not not2931(N9493,in2);
not not2932(N9494,R2);
not not2933(N9495,R3);
not not2934(N9507,in0);
not not2935(N9508,in1);
not not2936(N9509,in2);
not not2937(N9510,R1);
not not2938(N9522,in0);
not not2939(N9523,in1);
not not2940(N9524,in2);
not not2941(N9537,in1);
not not2942(N9538,R0);
not not2943(N9539,R1);
not not2944(N9552,in0);
not not2945(N9553,in1);
not not2946(N9554,R1);
not not2947(N9555,R2);
not not2948(N9567,in0);
not not2949(N9568,in2);
not not2950(N9569,R2);
not not2951(N9582,in0);
not not2952(N9583,in1);
not not2953(N9584,R1);
not not2954(N9585,R2);
not not2955(N9597,in0);
not not2956(N9598,in1);
not not2957(N9599,in2);
not not2958(N9600,R1);
not not2959(N9601,R2);
not not2960(N9612,in0);
not not2961(N9613,in2);
not not2962(N9614,R1);
not not2963(N9615,R2);
not not2964(N9627,in0);
not not2965(N9628,in1);
not not2966(N9629,R2);
not not2967(N9630,R3);
not not2968(N9642,in0);
not not2969(N9643,in1);
not not2970(N9644,in2);
not not2971(N9645,R0);
not not2972(N9657,in0);
not not2973(N9658,in1);
not not2974(N9659,R0);
not not2975(N9660,R1);
not not2976(N9672,in0);
not not2977(N9673,in2);
not not2978(N9674,R3);
not not2979(N9687,in0);
not not2980(N9688,in1);
not not2981(N9689,in2);
not not2982(N9690,R1);
not not2983(N9691,R2);
not not2984(N9702,in1);
not not2985(N9703,in2);
not not2986(N9704,R1);
not not2987(N9705,R2);
not not2988(N9717,in0);
not not2989(N9718,in2);
not not2990(N9719,R0);
not not2991(N9732,in0);
not not2992(N9733,R1);
not not2993(N9734,R2);
not not2994(N9747,in1);
not not2995(N9748,R0);
not not2996(N9749,R1);
not not2997(N9750,R3);
not not2998(N9761,in2);
not not2999(N9762,R0);
not not3000(N9763,R1);
not not3001(N9764,R3);
not not3002(N9775,in0);
not not3003(N9776,in1);
not not3004(N9777,in2);
not not3005(N9778,R0);
not not3006(N9789,in0);
not not3007(N9790,in1);
not not3008(N9791,in2);
not not3009(N9792,R1);
not not3010(N9803,in0);
not not3011(N9804,R0);
not not3012(N9817,in0);
not not3013(N9818,in1);
not not3014(N9831,in2);
not not3015(N9832,R3);
not not3016(N9845,in0);
not not3017(N9846,in2);
not not3018(N9847,R0);
not not3019(N9859,R0);
not not3020(N9860,R1);
not not3021(N9861,R3);
not not3022(N9873,in2);
not not3023(N9874,R0);
not not3024(N9875,R3);
not not3025(N9887,in1);
not not3026(N9888,R2);
not not3027(N9901,in2);
not not3028(N9902,R2);
not not3029(N9915,R0);
not not3030(N9916,R1);
not not3031(N9929,in1);
not not3032(N9930,in2);
not not3033(N9931,R0);
not not3034(N9932,R1);
not not3035(N9933,R3);
not not3036(N9943,R0);
not not3037(N9944,R2);
not not3038(N9957,in2);
not not3039(N9958,R0);
not not3040(N9959,R3);
not not3041(N9971,R0);
not not3042(N9972,R1);
not not3043(N9973,R3);
not not3044(N9985,in0);
not not3045(N9986,in1);
not not3046(N9987,R1);
not not3047(N9999,in0);
not not3048(N10000,R1);
not not3049(N10001,R3);
not not3050(N10013,in0);
not not3051(N10014,R2);
not not3052(N10015,R3);
not not3053(N10027,in0);
not not3054(N10028,in1);
not not3055(N10029,R2);
not not3056(N10041,in0);
not not3057(N10042,in1);
not not3058(N10043,in2);
not not3059(N10044,R1);
not not3060(N10045,R2);
not not3061(N10055,in0);
not not3062(N10056,in2);
not not3063(N10057,R1);
not not3064(N10069,in0);
not not3065(N10070,in1);
not not3066(N10083,R1);
not not3067(N10084,R2);
not not3068(N10085,R3);
not not3069(N10097,in0);
not not3070(N10098,R1);
not not3071(N10111,in0);
not not3072(N10112,in1);
not not3073(N10125,in0);
not not3074(N10126,in2);
not not3075(N10139,in0);
not not3076(N10140,R1);
not not3077(N10141,R2);
not not3078(N10153,in0);
not not3079(N10154,R0);
not not3080(N10155,R1);
not not3081(N10156,R3);
not not3082(N10167,in1);
not not3083(N10168,R2);
not not3084(N10169,R3);
not not3085(N10181,R0);
not not3086(N10182,R1);
not not3087(N10183,R2);
not not3088(N10195,in0);
not not3089(N10196,in2);
not not3090(N10197,R1);
not not3091(N10198,R2);
not not3092(N10209,in0);
not not3093(N10210,in2);
not not3094(N10211,R2);
not not3095(N10223,in0);
not not3096(N10224,in1);
not not3097(N10225,R0);
not not3098(N10226,R2);
not not3099(N10237,in2);
not not3100(N10238,R0);
not not3101(N10239,R2);
not not3102(N10251,in1);
not not3103(N10252,R0);
not not3104(N10253,R3);
not not3105(N10265,in2);
not not3106(N10266,R0);
not not3107(N10267,R1);
not not3108(N10279,in0);
not not3109(N10280,in1);
not not3110(N10281,R0);
not not3111(N10293,in1);
not not3112(N10294,R2);
not not3113(N10307,in0);
not not3114(N10308,in1);
not not3115(N10320,in2);
not not3116(N10321,R1);
not not3117(N10333,in0);
not not3118(N10334,in1);
not not3119(N10335,R0);
not not3120(N10346,in0);
not not3121(N10347,in2);
not not3122(N10348,R0);
not not3123(N10359,in0);
not not3124(N10372,in2);
not not3125(N10373,R0);
not not3126(N10374,R1);
not not3127(N10385,in2);
not not3128(N10386,R1);
not not3129(N10387,R3);
not not3130(N10398,in0);
not not3131(N10399,R1);
not not3132(N10411,R0);
not not3133(N10412,R1);
not not3134(N10413,R2);
not not3135(N10424,in2);
not not3136(N10425,R1);
not not3137(N10426,R2);
not not3138(N10437,in0);
not not3139(N10438,in1);
not not3140(N10439,R3);
not not3141(N10450,in0);
not not3142(N10451,in1);
not not3143(N10452,in2);
not not3144(N10463,in0);
not not3145(N10464,in2);
not not3146(N10465,R1);
not not3147(N10466,R2);
not not3148(N10476,in1);
not not3149(N10477,in2);
not not3150(N10478,R1);
not not3151(N10479,R2);
not not3152(N10489,in0);
not not3153(N10490,in1);
not not3154(N10491,R1);
not not3155(N10492,R2);
not not3156(N10502,in1);
not not3157(N10503,in2);
not not3158(N10504,R2);
not not3159(N10515,in1);
not not3160(N10516,R3);
not not3161(N10528,R1);
not not3162(N10529,R3);
not not3163(N10541,in0);
not not3164(N10542,R1);
not not3165(N10543,R2);
not not3166(N10554,in0);
not not3167(N10555,in2);
not not3168(N10567,in0);
not not3169(N10568,in2);
not not3170(N10580,in1);
not not3171(N10581,R1);
not not3172(N10582,R2);
not not3173(N10583,R3);
not not3174(N10593,in0);
not not3175(N10594,in1);
not not3176(N10595,R1);
not not3177(N10596,R3);
not not3178(N10606,R1);
not not3179(N10619,R1);
not not3180(N10632,in0);
not not3181(N10633,R1);
not not3182(N10634,R2);
not not3183(N10645,in1);
not not3184(N10646,R1);
not not3185(N10647,R2);
not not3186(N10658,in0);
not not3187(N10659,in1);
not not3188(N10660,R0);
not not3189(N10661,R1);
not not3190(N10671,in2);
not not3191(N10672,R0);
not not3192(N10684,in0);
not not3193(N10685,R0);
not not3194(N10697,in1);
not not3195(N10698,R0);
not not3196(N10699,R1);
not not3197(N10700,R2);
not not3198(N10710,R3);
not not3199(N10723,R1);
not not3200(N10724,R2);
not not3201(N10736,R1);
not not3202(N10737,R2);
not not3203(N10749,in0);
not not3204(N10750,R1);
not not3205(N10751,R2);
not not3206(N10762,in2);
not not3207(N10763,R0);
not not3208(N10764,R1);
not not3209(N10775,in0);
not not3210(N10776,R0);
not not3211(N10777,R1);
not not3212(N10788,in2);
not not3213(N10789,R1);
not not3214(N10790,R3);
not not3215(N10801,in1);
not not3216(N10802,R1);
not not3217(N10803,R3);
not not3218(N10814,in2);
not not3219(N10815,R0);
not not3220(N10816,R1);
not not3221(N10827,R1);
not not3222(N10839,R0);
not not3223(N10851,R1);
not not3224(N10852,R3);
not not3225(N10863,in1);
not not3226(N10864,R0);
not not3227(N10875,in0);
not not3228(N10876,in1);
not not3229(N10887,in1);
not not3230(N10899,in1);
not not3231(N10911,R0);
not not3232(N10935,in1);
not not3233(N10936,in2);
not not3234(N10937,R0);
not not3235(N10947,R0);
not not3236(N10959,in1);
not not3237(N10960,in2);
not not3238(N10961,R3);
not not3239(N10971,in1);
not not3240(N10983,in1);
not not3241(N10984,R0);
not not3242(N10995,in0);
not not3243(N11007,in1);
not not3244(N11008,R0);
not not3245(N11019,R1);
not not3246(N11020,R3);
not not3247(N11031,in2);
not not3248(N11043,in1);
not not3249(N11044,R0);
not not3250(N11067,in0);
not not3251(N11068,R3);
not not3252(N11079,in1);
not not3253(N11080,R3);
not not3254(N11091,R0);
not not3255(N11092,R1);
not not3256(N11103,R3);
not not3257(N11115,in2);
not not3258(N11127,R2);
not not3259(N11139,in1);
not not3260(N11140,R2);
not not3261(N11151,R0);
not not3262(N11162,R1);
not not3263(N11163,R2);
not not3264(N11173,in1);
not not3265(N11174,R2);
not not3266(N11184,in0);
not not3267(N11185,R0);
not not3268(N11195,R3);
not not3269(N11206,in1);
not not3270(N11217,in2);
not not3271(N11228,R1);
not not3272(N11239,R2);
not not3273(N11250,in1);
not not3274(N11272,R1);
not not3275(N11273,R3);
not not3276(N11283,in1);
not not3277(N11294,R1);
not not3278(N11305,R1);
not not3279(N11316,in2);
not not3280(N11327,R0);
not not3281(N11337,R3);
not not3282(N11357,in1);
not not3283(N11367,R1);
not not3284(N11376,in0);
not not3285(N11377,in1);
not not3286(N11378,in2);
not not3287(N11379,R0);
not not3288(N11380,R4);
not not3289(N11381,R5);
not not3290(N11392,in1);
not not3291(N11393,R0);
not not3292(N11394,R1);
not not3293(N11395,R2);
not not3294(N11396,R3);
not not3295(N11397,R4);
not not3296(N11398,R5);
not not3297(N11408,in1);
not not3298(N11409,R0);
not not3299(N11410,R2);
not not3300(N11411,R3);
not not3301(N11412,R4);
not not3302(N11413,R5);
not not3303(N11424,in1);
not not3304(N11425,R0);
not not3305(N11426,R2);
not not3306(N11427,R3);
not not3307(N11428,R4);
not not3308(N11429,R5);
not not3309(N11440,in2);
not not3310(N11441,R0);
not not3311(N11442,R1);
not not3312(N11443,R3);
not not3313(N11444,R4);
not not3314(N11445,R5);
not not3315(N11456,in1);
not not3316(N11457,R0);
not not3317(N11458,R1);
not not3318(N11459,R2);
not not3319(N11460,R4);
not not3320(N11461,R5);
not not3321(N11472,in1);
not not3322(N11473,in2);
not not3323(N11474,R0);
not not3324(N11475,R2);
not not3325(N11476,R3);
not not3326(N11477,R4);
not not3327(N11478,R5);
not not3328(N11488,in1);
not not3329(N11489,R1);
not not3330(N11490,R2);
not not3331(N11491,R3);
not not3332(N11492,R5);
not not3333(N11503,in0);
not not3334(N11504,in2);
not not3335(N11505,R1);
not not3336(N11506,R4);
not not3337(N11507,R5);
not not3338(N11518,in0);
not not3339(N11519,in2);
not not3340(N11520,R0);
not not3341(N11521,R1);
not not3342(N11522,R2);
not not3343(N11533,in0);
not not3344(N11534,in2);
not not3345(N11535,R0);
not not3346(N11536,R1);
not not3347(N11537,R2);
not not3348(N11538,R5);
not not3349(N11548,in0);
not not3350(N11549,in1);
not not3351(N11550,in2);
not not3352(N11551,R0);
not not3353(N11552,R1);
not not3354(N11553,R4);
not not3355(N11563,in0);
not not3356(N11564,in2);
not not3357(N11565,R1);
not not3358(N11566,R2);
not not3359(N11567,R3);
not not3360(N11568,R4);
not not3361(N11578,R0);
not not3362(N11579,R1);
not not3363(N11580,R2);
not not3364(N11581,R4);
not not3365(N11582,R5);
not not3366(N11593,in0);
not not3367(N11594,R0);
not not3368(N11595,R3);
not not3369(N11596,R4);
not not3370(N11597,R5);
not not3371(N11607,R1);
not not3372(N11608,R2);
not not3373(N11609,R3);
not not3374(N11610,R4);
not not3375(N11611,R5);
not not3376(N11621,in0);
not not3377(N11622,R0);
not not3378(N11623,R1);
not not3379(N11624,R4);
not not3380(N11625,R5);
not not3381(N11635,R1);
not not3382(N11636,R2);
not not3383(N11637,R3);
not not3384(N11638,R5);
not not3385(N11649,in1);
not not3386(N11650,R0);
not not3387(N11651,R3);
not not3388(N11652,R4);
not not3389(N11663,in2);
not not3390(N11664,R1);
not not3391(N11665,R2);
not not3392(N11666,R3);
not not3393(N11667,R4);
not not3394(N11677,in0);
not not3395(N11678,in1);
not not3396(N11679,R0);
not not3397(N11680,R3);
not not3398(N11681,R4);
not not3399(N11691,in2);
not not3400(N11692,R0);
not not3401(N11693,R1);
not not3402(N11694,R3);
not not3403(N11695,R4);
not not3404(N11705,in0);
not not3405(N11706,R3);
not not3406(N11707,R4);
not not3407(N11708,R5);
not not3408(N11719,in0);
not not3409(N11720,in1);
not not3410(N11721,R1);
not not3411(N11722,R4);
not not3412(N11733,in1);
not not3413(N11734,R0);
not not3414(N11735,R4);
not not3415(N11736,R5);
not not3416(N11747,in1);
not not3417(N11748,R0);
not not3418(N11749,R4);
not not3419(N11750,R5);
not not3420(N11761,in2);
not not3421(N11762,R0);
not not3422(N11763,R1);
not not3423(N11764,R3);
not not3424(N11775,in0);
not not3425(N11776,in2);
not not3426(N11777,R0);
not not3427(N11778,R3);
not not3428(N11779,R4);
not not3429(N11789,in0);
not not3430(N11790,in1);
not not3431(N11791,in2);
not not3432(N11792,R2);
not not3433(N11803,R0);
not not3434(N11804,R2);
not not3435(N11805,R3);
not not3436(N11806,R4);
not not3437(N11807,R5);
not not3438(N11817,R0);
not not3439(N11818,R2);
not not3440(N11819,R3);
not not3441(N11820,R4);
not not3442(N11821,R5);
not not3443(N11831,in0);
not not3444(N11832,in1);
not not3445(N11833,R0);
not not3446(N11834,R2);
not not3447(N11835,R4);
not not3448(N11845,R1);
not not3449(N11846,R2);
not not3450(N11847,R3);
not not3451(N11848,R4);
not not3452(N11849,R5);
not not3453(N11859,in1);
not not3454(N11860,R0);
not not3455(N11861,R1);
not not3456(N11862,R2);
not not3457(N11873,in2);
not not3458(N11874,R0);
not not3459(N11875,R1);
not not3460(N11876,R2);
not not3461(N11877,R3);
not not3462(N11887,in1);
not not3463(N11888,in2);
not not3464(N11889,R1);
not not3465(N11890,R5);
not not3466(N11901,in0);
not not3467(N11902,in1);
not not3468(N11903,R0);
not not3469(N11904,R4);
not not3470(N11905,R5);
not not3471(N11915,in1);
not not3472(N11916,R0);
not not3473(N11917,R1);
not not3474(N11918,R2);
not not3475(N11919,R5);
not not3476(N11929,in1);
not not3477(N11930,in2);
not not3478(N11931,R1);
not not3479(N11932,R2);
not not3480(N11943,in0);
not not3481(N11944,in1);
not not3482(N11945,R0);
not not3483(N11946,R4);
not not3484(N11947,R5);
not not3485(N11957,in0);
not not3486(N11958,R0);
not not3487(N11959,R1);
not not3488(N11960,R4);
not not3489(N11961,R5);
not not3490(N11971,in0);
not not3491(N11972,in2);
not not3492(N11973,R0);
not not3493(N11974,R1);
not not3494(N11975,R3);
not not3495(N11985,in2);
not not3496(N11986,R0);
not not3497(N11987,R3);
not not3498(N11988,R5);
not not3499(N11999,in1);
not not3500(N12000,R0);
not not3501(N12001,R1);
not not3502(N12002,R3);
not not3503(N12013,in1);
not not3504(N12014,in2);
not not3505(N12015,R0);
not not3506(N12016,R1);
not not3507(N12017,R2);
not not3508(N12027,in0);
not not3509(N12028,in2);
not not3510(N12029,R1);
not not3511(N12030,R2);
not not3512(N12031,R5);
not not3513(N12041,in0);
not not3514(N12042,R0);
not not3515(N12043,R1);
not not3516(N12044,R2);
not not3517(N12045,R3);
not not3518(N12055,in0);
not not3519(N12056,in1);
not not3520(N12057,in2);
not not3521(N12058,R0);
not not3522(N12069,in0);
not not3523(N12070,in2);
not not3524(N12071,R0);
not not3525(N12072,R4);
not not3526(N12073,R5);
not not3527(N12083,in2);
not not3528(N12084,R3);
not not3529(N12085,R4);
not not3530(N12096,R0);
not not3531(N12097,R1);
not not3532(N12098,R3);
not not3533(N12099,R4);
not not3534(N12109,in0);
not not3535(N12110,in1);
not not3536(N12111,in2);
not not3537(N12112,R0);
not not3538(N12122,R0);
not not3539(N12123,R1);
not not3540(N12124,R2);
not not3541(N12125,R5);
not not3542(N12135,R0);
not not3543(N12136,R1);
not not3544(N12137,R4);
not not3545(N12138,R5);
not not3546(N12148,in1);
not not3547(N12149,R0);
not not3548(N12150,R3);
not not3549(N12151,R4);
not not3550(N12161,in1);
not not3551(N12162,R0);
not not3552(N12163,R1);
not not3553(N12164,R2);
not not3554(N12174,in2);
not not3555(N12175,R2);
not not3556(N12176,R5);
not not3557(N12187,in1);
not not3558(N12188,R0);
not not3559(N12189,R2);
not not3560(N12190,R4);
not not3561(N12200,in2);
not not3562(N12201,R0);
not not3563(N12202,R5);
not not3564(N12213,in0);
not not3565(N12214,R0);
not not3566(N12215,R1);
not not3567(N12216,R4);
not not3568(N12226,in2);
not not3569(N12227,R0);
not not3570(N12228,R3);
not not3571(N12229,R4);
not not3572(N12230,R5);
not not3573(N12239,in1);
not not3574(N12240,in2);
not not3575(N12241,R1);
not not3576(N12252,in0);
not not3577(N12253,R1);
not not3578(N12254,R2);
not not3579(N12255,R3);
not not3580(N12265,in1);
not not3581(N12266,R1);
not not3582(N12267,R2);
not not3583(N12268,R5);
not not3584(N12278,in2);
not not3585(N12279,R1);
not not3586(N12280,R2);
not not3587(N12281,R5);
not not3588(N12291,R0);
not not3589(N12292,R1);
not not3590(N12293,R2);
not not3591(N12304,in2);
not not3592(N12305,R0);
not not3593(N12306,R1);
not not3594(N12317,in1);
not not3595(N12318,in2);
not not3596(N12319,R0);
not not3597(N12320,R1);
not not3598(N12330,in1);
not not3599(N12331,R1);
not not3600(N12332,R3);
not not3601(N12343,in1);
not not3602(N12344,in2);
not not3603(N12345,R2);
not not3604(N12346,R4);
not not3605(N12356,in2);
not not3606(N12357,R3);
not not3607(N12358,R4);
not not3608(N12369,in0);
not not3609(N12370,R2);
not not3610(N12371,R3);
not not3611(N12382,in1);
not not3612(N12383,R2);
not not3613(N12384,R4);
not not3614(N12385,R5);
not not3615(N12395,in1);
not not3616(N12396,R0);
not not3617(N12397,R1);
not not3618(N12398,R3);
not not3619(N12408,in0);
not not3620(N12409,in1);
not not3621(N12410,in2);
not not3622(N12411,R0);
not not3623(N12421,in1);
not not3624(N12422,R1);
not not3625(N12423,R3);
not not3626(N12424,R4);
not not3627(N12434,in1);
not not3628(N12435,in2);
not not3629(N12436,R1);
not not3630(N12437,R4);
not not3631(N12447,in1);
not not3632(N12448,R0);
not not3633(N12449,R4);
not not3634(N12450,R5);
not not3635(N12460,in1);
not not3636(N12461,in2);
not not3637(N12462,R4);
not not3638(N12463,R5);
not not3639(N12473,in1);
not not3640(N12474,in2);
not not3641(N12475,R0);
not not3642(N12476,R1);
not not3643(N12486,in1);
not not3644(N12487,R3);
not not3645(N12488,R4);
not not3646(N12499,in0);
not not3647(N12500,R0);
not not3648(N12501,R3);
not not3649(N12502,R4);
not not3650(N12512,R2);
not not3651(N12513,R3);
not not3652(N12514,R4);
not not3653(N12515,R5);
not not3654(N12525,R0);
not not3655(N12526,R1);
not not3656(N12527,R2);
not not3657(N12528,R3);
not not3658(N12538,in1);
not not3659(N12539,in2);
not not3660(N12540,R4);
not not3661(N12551,in0);
not not3662(N12552,in2);
not not3663(N12553,R0);
not not3664(N12554,R4);
not not3665(N12564,in1);
not not3666(N12565,R1);
not not3667(N12566,R5);
not not3668(N12577,in2);
not not3669(N12578,R1);
not not3670(N12579,R5);
not not3671(N12590,R0);
not not3672(N12591,R1);
not not3673(N12592,R2);
not not3674(N12593,R5);
not not3675(N12603,R0);
not not3676(N12604,R1);
not not3677(N12605,R2);
not not3678(N12606,R4);
not not3679(N12616,R0);
not not3680(N12617,R3);
not not3681(N12618,R5);
not not3682(N12629,in2);
not not3683(N12630,R1);
not not3684(N12631,R3);
not not3685(N12632,R4);
not not3686(N12642,in1);
not not3687(N12643,in2);
not not3688(N12644,R1);
not not3689(N12645,R4);
not not3690(N12655,in0);
not not3691(N12656,in1);
not not3692(N12657,R1);
not not3693(N12658,R4);
not not3694(N12668,in2);
not not3695(N12669,R1);
not not3696(N12670,R4);
not not3697(N12671,R5);
not not3698(N12681,R4);
not not3699(N12682,R5);
not not3700(N12693,R3);
not not3701(N12694,R4);
not not3702(N12705,in1);
not not3703(N12706,R3);
not not3704(N12707,R5);
not not3705(N12717,R1);
not not3706(N12718,R2);
not not3707(N12719,R3);
not not3708(N12729,in1);
not not3709(N12730,R3);
not not3710(N12731,R4);
not not3711(N12741,in0);
not not3712(N12742,R1);
not not3713(N12743,R3);
not not3714(N12753,R0);
not not3715(N12754,R3);
not not3716(N12765,in1);
not not3717(N12766,R2);
not not3718(N12777,in1);
not not3719(N12778,in2);
not not3720(N12779,R0);
not not3721(N12789,in0);
not not3722(N12790,in1);
not not3723(N12791,R0);
not not3724(N12801,in0);
not not3725(N12802,in1);
not not3726(N12803,R2);
not not3727(N12813,in0);
not not3728(N12814,in2);
not not3729(N12815,R0);
not not3730(N12816,R3);
not not3731(N12825,in1);
not not3732(N12826,R0);
not not3733(N12827,R4);
not not3734(N12828,R5);
not not3735(N12837,in1);
not not3736(N12838,in2);
not not3737(N12839,R0);
not not3738(N12840,R2);
not not3739(N12849,in2);
not not3740(N12850,R2);
not not3741(N12851,R4);
not not3742(N12861,in0);
not not3743(N12862,in1);
not not3744(N12863,R0);
not not3745(N12873,R1);
not not3746(N12874,R4);
not not3747(N12885,R1);
not not3748(N12886,R4);
not not3749(N12897,in0);
not not3750(N12898,in1);
not not3751(N12899,R1);
not not3752(N12909,in1);
not not3753(N12910,in2);
not not3754(N12911,R4);
not not3755(N12912,R5);
not not3756(N12921,in0);
not not3757(N12922,R2);
not not3758(N12933,in1);
not not3759(N12934,in2);
not not3760(N12945,in1);
not not3761(N12946,R1);
not not3762(N12947,R2);
not not3763(N12957,in1);
not not3764(N12958,in2);
not not3765(N12959,R3);
not not3766(N12969,in1);
not not3767(N12970,R5);
not not3768(N12981,in1);
not not3769(N12982,R0);
not not3770(N12983,R4);
not not3771(N12993,in2);
not not3772(N12994,R3);
not not3773(N13005,R1);
not not3774(N13006,R3);
not not3775(N13007,R4);
not not3776(N13008,R5);
not not3777(N13017,in1);
not not3778(N13018,R0);
not not3779(N13019,R1);
not not3780(N13020,R5);
not not3781(N13029,in1);
not not3782(N13030,R2);
not not3783(N13031,R3);
not not3784(N13041,R2);
not not3785(N13042,R4);
not not3786(N13043,R5);
not not3787(N13053,in2);
not not3788(N13054,R0);
not not3789(N13055,R1);
not not3790(N13056,R2);
not not3791(N13065,in2);
not not3792(N13066,R0);
not not3793(N13067,R1);
not not3794(N13068,R2);
not not3795(N13077,in2);
not not3796(N13078,R0);
not not3797(N13079,R1);
not not3798(N13089,in1);
not not3799(N13090,R1);
not not3800(N13091,R2);
not not3801(N13101,in2);
not not3802(N13102,R1);
not not3803(N13103,R2);
not not3804(N13113,R3);
not not3805(N13114,R4);
not not3806(N13125,R0);
not not3807(N13126,R1);
not not3808(N13127,R3);
not not3809(N13137,in0);
not not3810(N13138,R0);
not not3811(N13139,R1);
not not3812(N13149,in2);
not not3813(N13150,R0);
not not3814(N13151,R2);
not not3815(N13161,in2);
not not3816(N13162,R0);
not not3817(N13163,R2);
not not3818(N13173,in0);
not not3819(N13174,in2);
not not3820(N13175,R5);
not not3821(N13185,in0);
not not3822(N13186,R2);
not not3823(N13187,R4);
not not3824(N13197,in0);
not not3825(N13198,in1);
not not3826(N13199,R1);
not not3827(N13209,in1);
not not3828(N13210,in2);
not not3829(N13211,R1);
not not3830(N13212,R3);
not not3831(N13221,in0);
not not3832(N13222,in2);
not not3833(N13223,R1);
not not3834(N13233,R2);
not not3835(N13234,R4);
not not3836(N13235,R5);
not not3837(N13245,R4);
not not3838(N13246,R5);
not not3839(N13257,in1);
not not3840(N13258,R0);
not not3841(N13259,R4);
not not3842(N13260,R5);
not not3843(N13269,in1);
not not3844(N13270,R0);
not not3845(N13271,R1);
not not3846(N13272,R4);
not not3847(N13281,in2);
not not3848(N13282,R2);
not not3849(N13283,R4);
not not3850(N13293,R2);
not not3851(N13294,R5);
not not3852(N13305,in0);
not not3853(N13306,in2);
not not3854(N13307,R0);
not not3855(N13317,R1);
not not3856(N13318,R2);
not not3857(N13329,in2);
not not3858(N13330,R2);
not not3859(N13331,R3);
not not3860(N13341,in0);
not not3861(N13342,R3);
not not3862(N13343,R4);
not not3863(N13353,in1);
not not3864(N13354,in2);
not not3865(N13355,R0);
not not3866(N13365,in1);
not not3867(N13366,R1);
not not3868(N13367,R2);
not not3869(N13368,R4);
not not3870(N13377,in2);
not not3871(N13378,R1);
not not3872(N13379,R4);
not not3873(N13389,in0);
not not3874(N13390,in2);
not not3875(N13391,R4);
not not3876(N13401,R1);
not not3877(N13412,R1);
not not3878(N13423,R0);
not not3879(N13424,R1);
not not3880(N13434,in1);
not not3881(N13435,R1);
not not3882(N13436,R4);
not not3883(N13445,in2);
not not3884(N13456,in0);
not not3885(N13457,R0);
not not3886(N13458,R4);
not not3887(N13467,in2);
not not3888(N13468,R1);
not not3889(N13469,R4);
not not3890(N13478,R0);
not not3891(N13479,R4);
not not3892(N13489,in1);
not not3893(N13490,R5);
not not3894(N13500,in0);
not not3895(N13501,in1);
not not3896(N13511,in2);
not not3897(N13512,R5);
not not3898(N13522,in1);
not not3899(N13523,R1);
not not3900(N13524,R5);
not not3901(N13533,in1);
not not3902(N13534,R1);
not not3903(N13535,R5);
not not3904(N13544,in1);
not not3905(N13545,R1);
not not3906(N13546,R3);
not not3907(N13555,R2);
not not3908(N13556,R4);
not not3909(N13566,in1);
not not3910(N13567,R1);
not not3911(N13577,in0);
not not3912(N13578,R0);
not not3913(N13579,R4);
not not3914(N13588,in0);
not not3915(N13589,R0);
not not3916(N13590,R4);
not not3917(N13599,in1);
not not3918(N13600,in2);
not not3919(N13610,in0);
not not3920(N13611,R0);
not not3921(N13612,R4);
not not3922(N13621,R2);
not not3923(N13622,R4);
not not3924(N13632,R1);
not not3925(N13633,R4);
not not3926(N13634,R5);
not not3927(N13643,in2);
not not3928(N13654,R1);
not not3929(N13655,R2);
not not3930(N13665,in1);
not not3931(N13666,R1);
not not3932(N13676,R4);
not not3933(N13687,in0);
not not3934(N13698,R1);
not not3935(N13699,R3);
not not3936(N13709,in1);
not not3937(N13710,R1);
not not3938(N13711,R5);
not not3939(N13720,in2);
not not3940(N13721,R2);
not not3941(N13722,R5);
not not3942(N13731,R0);
not not3943(N13732,R1);
not not3944(N13733,R5);
not not3945(N13742,in1);
not not3946(N13743,in2);
not not3947(N13753,R0);
not not3948(N13754,R5);
not not3949(N13764,in2);
not not3950(N13765,R1);
not not3951(N13766,R3);
not not3952(N13775,in1);
not not3953(N13776,R3);
not not3954(N13786,in1);
not not3955(N13787,R3);
not not3956(N13797,in2);
not not3957(N13798,R1);
not not3958(N13808,R0);
not not3959(N13809,R5);
not not3960(N13819,R0);
not not3961(N13820,R5);
not not3962(N13830,R0);
not not3963(N13831,R1);
not not3964(N13841,R3);
not not3965(N13842,R4);
not not3966(N13852,R1);
not not3967(N13853,R4);
not not3968(N13863,R2);
not not3969(N13864,R3);
not not3970(N13874,in2);
not not3971(N13875,R1);
not not3972(N13876,R2);
not not3973(N13885,in0);
not not3974(N13886,in2);
not not3975(N13896,R3);
not not3976(N13907,R0);
not not3977(N13908,R1);
not not3978(N13909,R2);
not not3979(N13918,in2);
not not3980(N13919,R2);
not not3981(N13929,R0);
not not3982(N13930,R2);
not not3983(N13940,R0);
not not3984(N13941,R1);
not not3985(N13942,R4);
not not3986(N13951,R4);
not not3987(N13962,R4);
not not3988(N13982,in2);
not not3989(N13983,R4);
not not3990(N13992,R0);
not not3991(N13993,R1);
not not3992(N14002,R0);
not not3993(N14003,R4);
not not3994(N14012,in2);
not not3995(N14013,R0);
not not3996(N14022,R0);
not not3997(N14023,R2);
not not3998(N14032,R0);
not not3999(N14033,R2);
not not4000(N14052,R4);
not not4001(N14053,R5);
not not4002(N14062,in0);
not not4003(N14072,R3);
not not4004(N14073,R4);
not not4005(N14082,in1);
not not4006(N14083,in2);
not not4007(N14092,R1);
not not4008(N14102,R2);
not not4009(N14122,R5);
not not4010(N14131,R5);
not not4011(N14140,in2);
not not4012(N14158,in0);
not not4013(N14185,R4);
not not4014(N14203,in2);
not not4015(N14211,R1);
not not4016(N14212,R2);
not not4017(N14213,R3);
not not4018(N14214,R4);
not not4019(N14215,R5);
not not4020(N14216,R6);
not not4021(N14217,R7);
not not4022(N14225,in2);
not not4023(N14226,R0);
not not4024(N14227,R2);
not not4025(N14228,R4);
not not4026(N14229,R5);
not not4027(N14230,R6);
not not4028(N14231,R7);
not not4029(N14239,in1);
not not4030(N14240,R1);
not not4031(N14241,R2);
not not4032(N14242,R3);
not not4033(N14243,R5);
not not4034(N14244,R6);
not not4035(N14245,R7);
not not4036(N14253,in2);
not not4037(N14254,R2);
not not4038(N14255,R3);
not not4039(N14256,R4);
not not4040(N14257,R5);
not not4041(N14258,R6);
not not4042(N14259,R7);
not not4043(N14267,in1);
not not4044(N14268,R0);
not not4045(N14269,R1);
not not4046(N14270,R2);
not not4047(N14271,R3);
not not4048(N14272,R6);
not not4049(N14280,in1);
not not4050(N14281,R1);
not not4051(N14282,R2);
not not4052(N14283,R3);
not not4053(N14284,R4);
not not4054(N14285,R6);
not not4055(N14293,in2);
not not4056(N14294,R0);
not not4057(N14295,R1);
not not4058(N14296,R4);
not not4059(N14297,R5);
not not4060(N14298,R7);
not not4061(N14306,in1);
not not4062(N14307,R0);
not not4063(N14308,R2);
not not4064(N14309,R4);
not not4065(N14310,R6);
not not4066(N14311,R7);
not not4067(N14319,in2);
not not4068(N14320,R0);
not not4069(N14321,R1);
not not4070(N14322,R2);
not not4071(N14323,R4);
not not4072(N14324,R7);
not not4073(N14332,R1);
not not4074(N14333,R2);
not not4075(N14334,R3);
not not4076(N14335,R4);
not not4077(N14336,R5);
not not4078(N14337,R6);
not not4079(N14345,in2);
not not4080(N14346,R0);
not not4081(N14347,R4);
not not4082(N14348,R5);
not not4083(N14349,R6);
not not4084(N14350,R7);
not not4085(N14358,R0);
not not4086(N14359,R3);
not not4087(N14360,R4);
not not4088(N14361,R5);
not not4089(N14362,R6);
not not4090(N14370,R1);
not not4091(N14371,R4);
not not4092(N14372,R5);
not not4093(N14373,R6);
not not4094(N14374,R7);
not not4095(N14382,in1);
not not4096(N14383,R0);
not not4097(N14384,R3);
not not4098(N14385,R6);
not not4099(N14386,R7);
not not4100(N14394,in1);
not not4101(N14395,in2);
not not4102(N14396,R3);
not not4103(N14397,R4);
not not4104(N14398,R6);
not not4105(N14406,R1);
not not4106(N14407,R2);
not not4107(N14408,R4);
not not4108(N14409,R6);
not not4109(N14410,R7);
not not4110(N14418,in2);
not not4111(N14419,R1);
not not4112(N14420,R3);
not not4113(N14421,R4);
not not4114(N14422,R5);
not not4115(N14430,in1);
not not4116(N14431,R0);
not not4117(N14432,R1);
not not4118(N14433,R4);
not not4119(N14434,R6);
not not4120(N14442,in0);
not not4121(N14443,R3);
not not4122(N14444,R5);
not not4123(N14445,R6);
not not4124(N14446,R7);
not not4125(N14454,in0);
not not4126(N14455,R3);
not not4127(N14456,R5);
not not4128(N14457,R6);
not not4129(N14458,R7);
not not4130(N14466,in1);
not not4131(N14467,in2);
not not4132(N14468,R4);
not not4133(N14469,R5);
not not4134(N14470,R6);
not not4135(N14478,R0);
not not4136(N14479,R1);
not not4137(N14480,R4);
not not4138(N14481,R6);
not not4139(N14482,R7);
not not4140(N14490,R0);
not not4141(N14491,R2);
not not4142(N14492,R4);
not not4143(N14493,R6);
not not4144(N14494,R7);
not not4145(N14502,in2);
not not4146(N14503,R0);
not not4147(N14504,R1);
not not4148(N14505,R4);
not not4149(N14506,R6);
not not4150(N14514,R1);
not not4151(N14515,R3);
not not4152(N14516,R4);
not not4153(N14517,R6);
not not4154(N14525,R1);
not not4155(N14526,R2);
not not4156(N14527,R3);
not not4157(N14528,R4);
not not4158(N14536,R1);
not not4159(N14537,R4);
not not4160(N14538,R5);
not not4161(N14539,R6);
not not4162(N14547,in1);
not not4163(N14548,R1);
not not4164(N14549,R3);
not not4165(N14550,R4);
not not4166(N14558,R0);
not not4167(N14559,R1);
not not4168(N14560,R3);
not not4169(N14561,R7);
not not4170(N14569,in1);
not not4171(N14570,R2);
not not4172(N14571,R5);
not not4173(N14572,R6);
not not4174(N14580,in2);
not not4175(N14581,R3);
not not4176(N14582,R4);
not not4177(N14583,R6);
not not4178(N14591,in1);
not not4179(N14592,R4);
not not4180(N14593,R5);
not not4181(N14594,R6);
not not4182(N14602,in2);
not not4183(N14603,R4);
not not4184(N14604,R5);
not not4185(N14605,R6);
not not4186(N14613,R2);
not not4187(N14614,R6);
not not4188(N14615,R7);
not not4189(N14623,in1);
not not4190(N14624,R2);
not not4191(N14625,R5);
not not4192(N14633,R0);
not not4193(N14634,R1);
not not4194(N14635,R6);
not not4195(N14643,R0);
not not4196(N14644,R5);
not not4197(N14645,R7);
not not4198(N14653,R2);
not not4199(N14654,R5);
not not4200(N14655,R6);
not not4201(N14663,in2);
not not4202(N14664,R2);
not not4203(N14672,R1);
not not4204(N14673,R7);
not not4205(N14681,R4);
not not4206(N14682,R7);
not not4207(N14690,R0);
not not4208(N14691,R6);
not not4209(N14699,R1);
not not4210(N14700,R6);
not not4211(N14714,R1);
not not4212(N14715,R2);
not not4213(N14716,R3);
not not4214(N14717,R6);
not not4215(N14724,R4);
not not4216(N14725,R7);
not not4217(N8900,R4);
not not4218(N8901,R6);
not not4219(N8902,R7);
not not4220(N8916,R4);
not not4221(N8917,R5);
not not4222(N8918,R6);
not not4223(N8919,R7);
not not4224(N8934,R4);
not not4225(N8935,R5);
not not4226(N8936,R6);
not not4227(N8951,R4);
not not4228(N8952,R5);
not not4229(N8953,R6);
not not4230(N8969,R6);
not not4231(N8970,R7);
not not4232(N8985,R5);
not not4233(N8986,R6);
not not4234(N8987,R7);
not not4235(N9000,R4);
not not4236(N9001,R5);
not not4237(N9002,R6);
not not4238(N9003,R7);
not not4239(N9016,R4);
not not4240(N9017,R5);
not not4241(N9018,R6);
not not4242(N9019,R7);
not not4243(N9034,R4);
not not4244(N9035,R6);
not not4245(N9049,R5);
not not4246(N9050,R6);
not not4247(N9051,R7);
not not4248(N9065,R4);
not not4249(N9066,R5);
not not4250(N9067,R6);
not not4251(N9080,R4);
not not4252(N9081,R5);
not not4253(N9082,R6);
not not4254(N9083,R7);
not not4255(N9097,R4);
not not4256(N9098,R6);
not not4257(N9099,R7);
not not4258(N9112,R4);
not not4259(N9113,R5);
not not4260(N9114,R6);
not not4261(N9115,R7);
not not4262(N9128,R4);
not not4263(N9129,R5);
not not4264(N9130,R6);
not not4265(N9131,R7);
not not4266(N9145,R3);
not not4267(N9146,R4);
not not4268(N9147,R7);
not not4269(N9161,R4);
not not4270(N9162,R5);
not not4271(N9163,R7);
not not4272(N9178,R5);
not not4273(N9179,R7);
not not4274(N9194,R5);
not not4275(N9195,R6);
not not4276(N9209,R4);
not not4277(N9210,R6);
not not4278(N9211,R7);
not not4279(N9226,R3);
not not4280(N9227,R5);
not not4281(N9241,R6);
not not4282(N9242,R7);
not not4283(N9256,R4);
not not4284(N9257,R6);
not not4285(N9270,R4);
not not4286(N9271,R6);
not not4287(N9272,R7);
not not4288(N9287,R4);
not not4289(N9301,R4);
not not4290(N9302,R7);
not not4291(N9316,R4);
not not4292(N9317,R7);
not not4293(N9330,R5);
not not4294(N9331,R6);
not not4295(N9332,R7);
not not4296(N9345,R4);
not not4297(N9346,R6);
not not4298(N9347,R7);
not not4299(N9360,R4);
not not4300(N9361,R6);
not not4301(N9362,R7);
not not4302(N9374,R4);
not not4303(N9375,R5);
not not4304(N9376,R6);
not not4305(N9377,R7);
not not4306(N9391,R4);
not not4307(N9392,R6);
not not4308(N9406,R6);
not not4309(N9407,R7);
not not4310(N9422,R5);
not not4311(N9436,R4);
not not4312(N9437,R7);
not not4313(N9451,R4);
not not4314(N9452,R5);
not not4315(N9466,R4);
not not4316(N9467,R5);
not not4317(N9480,R4);
not not4318(N9481,R6);
not not4319(N9482,R7);
not not4320(N9496,R5);
not not4321(N9497,R6);
not not4322(N9511,R4);
not not4323(N9512,R5);
not not4324(N9525,R3);
not not4325(N9526,R5);
not not4326(N9527,R7);
not not4327(N9540,R5);
not not4328(N9541,R6);
not not4329(N9542,R7);
not not4330(N9556,R6);
not not4331(N9557,R7);
not not4332(N9570,R5);
not not4333(N9571,R6);
not not4334(N9572,R7);
not not4335(N9586,R3);
not not4336(N9587,R4);
not not4337(N9602,R4);
not not4338(N9616,R5);
not not4339(N9617,R7);
not not4340(N9631,R6);
not not4341(N9632,R7);
not not4342(N9646,R4);
not not4343(N9647,R5);
not not4344(N9661,R3);
not not4345(N9662,R5);
not not4346(N9675,R4);
not not4347(N9676,R5);
not not4348(N9677,R7);
not not4349(N9692,R7);
not not4350(N9706,R4);
not not4351(N9707,R6);
not not4352(N9720,R4);
not not4353(N9721,R5);
not not4354(N9722,R6);
not not4355(N9735,R4);
not not4356(N9736,R6);
not not4357(N9737,R7);
not not4358(N9751,R6);
not not4359(N9765,R6);
not not4360(N9779,R5);
not not4361(N9793,R5);
not not4362(N9805,R4);
not not4363(N9806,R5);
not not4364(N9807,R7);
not not4365(N9819,R3);
not not4366(N9820,R5);
not not4367(N9821,R6);
not not4368(N9833,R4);
not not4369(N9834,R5);
not not4370(N9835,R6);
not not4371(N9848,R5);
not not4372(N9849,R6);
not not4373(N9862,R4);
not not4374(N9863,R7);
not not4375(N9876,R4);
not not4376(N9877,R7);
not not4377(N9889,R3);
not not4378(N9890,R5);
not not4379(N9891,R6);
not not4380(N9903,R3);
not not4381(N9904,R5);
not not4382(N9905,R6);
not not4383(N9917,R4);
not not4384(N9918,R5);
not not4385(N9919,R6);
not not4386(N9945,R5);
not not4387(N9946,R6);
not not4388(N9947,R7);
not not4389(N9960,R5);
not not4390(N9961,R6);
not not4391(N9974,R4);
not not4392(N9975,R5);
not not4393(N9988,R4);
not not4394(N9989,R7);
not not4395(N10002,R5);
not not4396(N10003,R7);
not not4397(N10016,R5);
not not4398(N10017,R6);
not not4399(N10030,R5);
not not4400(N10031,R6);
not not4401(N10058,R4);
not not4402(N10059,R7);
not not4403(N10071,R4);
not not4404(N10072,R5);
not not4405(N10073,R7);
not not4406(N10086,R6);
not not4407(N10087,R7);
not not4408(N10099,R5);
not not4409(N10100,R6);
not not4410(N10101,R7);
not not4411(N10113,R4);
not not4412(N10114,R6);
not not4413(N10115,R7);
not not4414(N10127,R4);
not not4415(N10128,R5);
not not4416(N10129,R7);
not not4417(N10142,R6);
not not4418(N10143,R7);
not not4419(N10157,R4);
not not4420(N10170,R4);
not not4421(N10171,R6);
not not4422(N10184,R4);
not not4423(N10185,R6);
not not4424(N10199,R4);
not not4425(N10212,R4);
not not4426(N10213,R5);
not not4427(N10227,R6);
not not4428(N10240,R4);
not not4429(N10241,R6);
not not4430(N10254,R5);
not not4431(N10255,R6);
not not4432(N10268,R3);
not not4433(N10269,R5);
not not4434(N10282,R4);
not not4435(N10283,R7);
not not4436(N10295,R4);
not not4437(N10296,R6);
not not4438(N10297,R7);
not not4439(N10309,R6);
not not4440(N10310,R7);
not not4441(N10322,R4);
not not4442(N10323,R7);
not not4443(N10336,R5);
not not4444(N10349,R5);
not not4445(N10360,R3);
not not4446(N10361,R4);
not not4447(N10362,R7);
not not4448(N10375,R5);
not not4449(N10388,R5);
not not4450(N10400,R4);
not not4451(N10401,R6);
not not4452(N10414,R4);
not not4453(N10427,R4);
not not4454(N10440,R7);
not not4455(N10453,R4);
not not4456(N10505,R6);
not not4457(N10517,R6);
not not4458(N10518,R7);
not not4459(N10530,R6);
not not4460(N10531,R7);
not not4461(N10544,R5);
not not4462(N10556,R3);
not not4463(N10557,R7);
not not4464(N10569,R6);
not not4465(N10570,R7);
not not4466(N10607,R4);
not not4467(N10608,R5);
not not4468(N10609,R7);
not not4469(N10620,R5);
not not4470(N10621,R6);
not not4471(N10622,R7);
not not4472(N10635,R7);
not not4473(N10648,R6);
not not4474(N10673,R4);
not not4475(N10674,R5);
not not4476(N10686,R5);
not not4477(N10687,R6);
not not4478(N10711,R4);
not not4479(N10712,R5);
not not4480(N10713,R7);
not not4481(N10725,R4);
not not4482(N10726,R7);
not not4483(N10738,R4);
not not4484(N10739,R6);
not not4485(N10752,R4);
not not4486(N10765,R4);
not not4487(N10778,R4);
not not4488(N10791,R7);
not not4489(N10804,R7);
not not4490(N10817,R7);
not not4491(N10828,R4);
not not4492(N10829,R6);
not not4493(N10840,R4);
not not4494(N10841,R5);
not not4495(N10853,R4);
not not4496(N10865,R5);
not not4497(N10877,R4);
not not4498(N10888,R6);
not not4499(N10889,R7);
not not4500(N10900,R4);
not not4501(N10901,R6);
not not4502(N10912,R4);
not not4503(N10913,R7);
not not4504(N10923,R4);
not not4505(N10924,R5);
not not4506(N10925,R6);
not not4507(N10948,R3);
not not4508(N10949,R5);
not not4509(N10972,R5);
not not4510(N10973,R6);
not not4511(N10985,R3);
not not4512(N10996,R5);
not not4513(N10997,R7);
not not4514(N11009,R7);
not not4515(N11021,R6);
not not4516(N11032,R3);
not not4517(N11033,R5);
not not4518(N11045,R6);
not not4519(N11055,R3);
not not4520(N11056,R6);
not not4521(N11057,R7);
not not4522(N11069,R5);
not not4523(N11081,R6);
not not4524(N11093,R3);
not not4525(N11104,R5);
not not4526(N11105,R6);
not not4527(N11116,R3);
not not4528(N11117,R6);
not not4529(N11128,R4);
not not4530(N11129,R5);
not not4531(N11141,R6);
not not4532(N11152,R7);
not not4533(N11196,R7);
not not4534(N11207,R3);
not not4535(N11218,R3);
not not4536(N11229,R4);
not not4537(N11240,R6);
not not4538(N11251,R4);
not not4539(N11261,R3);
not not4540(N11262,R5);
not not4541(N11284,R5);
not not4542(N11295,R6);
not not4543(N11306,R3);
not not4544(N11317,R4);
not not4545(N11347,R3);
not not4546(N11382,R6);
not not4547(N11383,R7);
not not4548(N11399,R7);
not not4549(N11414,R6);
not not4550(N11415,R7);
not not4551(N11430,R6);
not not4552(N11431,R7);
not not4553(N11446,R6);
not not4554(N11447,R7);
not not4555(N11462,R6);
not not4556(N11463,R7);
not not4557(N11479,R6);
not not4558(N11493,R6);
not not4559(N11494,R7);
not not4560(N11508,R6);
not not4561(N11509,R7);
not not4562(N11523,R6);
not not4563(N11524,R7);
not not4564(N11539,R6);
not not4565(N11554,R6);
not not4566(N11569,R6);
not not4567(N11583,R6);
not not4568(N11584,R7);
not not4569(N11598,R6);
not not4570(N11612,R7);
not not4571(N11626,R7);
not not4572(N11639,R6);
not not4573(N11640,R7);
not not4574(N11653,R5);
not not4575(N11654,R6);
not not4576(N11668,R6);
not not4577(N11682,R5);
not not4578(N11696,R6);
not not4579(N11709,R6);
not not4580(N11710,R7);
not not4581(N11723,R6);
not not4582(N11724,R7);
not not4583(N11737,R6);
not not4584(N11738,R7);
not not4585(N11751,R6);
not not4586(N11752,R7);
not not4587(N11765,R6);
not not4588(N11766,R7);
not not4589(N11780,R6);
not not4590(N11793,R6);
not not4591(N11794,R7);
not not4592(N11808,R6);
not not4593(N11822,R6);
not not4594(N11836,R6);
not not4595(N11850,R7);
not not4596(N11863,R6);
not not4597(N11864,R7);
not not4598(N11878,R6);
not not4599(N11891,R6);
not not4600(N11892,R7);
not not4601(N11906,R7);
not not4602(N11920,R7);
not not4603(N11933,R6);
not not4604(N11934,R7);
not not4605(N11948,R7);
not not4606(N11962,R6);
not not4607(N11976,R7);
not not4608(N11989,R6);
not not4609(N11990,R7);
not not4610(N12003,R4);
not not4611(N12004,R6);
not not4612(N12018,R4);
not not4613(N12032,R6);
not not4614(N12046,R6);
not not4615(N12059,R6);
not not4616(N12060,R7);
not not4617(N12074,R7);
not not4618(N12086,R5);
not not4619(N12087,R7);
not not4620(N12100,R6);
not not4621(N12113,R6);
not not4622(N12126,R6);
not not4623(N12139,R7);
not not4624(N12152,R6);
not not4625(N12165,R7);
not not4626(N12177,R6);
not not4627(N12178,R7);
not not4628(N12191,R6);
not not4629(N12203,R6);
not not4630(N12204,R7);
not not4631(N12217,R6);
not not4632(N12242,R6);
not not4633(N12243,R7);
not not4634(N12256,R7);
not not4635(N12269,R7);
not not4636(N12282,R7);
not not4637(N12294,R6);
not not4638(N12295,R7);
not not4639(N12307,R6);
not not4640(N12308,R7);
not not4641(N12321,R6);
not not4642(N12333,R5);
not not4643(N12334,R7);
not not4644(N12347,R7);
not not4645(N12359,R6);
not not4646(N12360,R7);
not not4647(N12372,R6);
not not4648(N12373,R7);
not not4649(N12386,R7);
not not4650(N12399,R7);
not not4651(N12412,R6);
not not4652(N12425,R7);
not not4653(N12438,R5);
not not4654(N12451,R6);
not not4655(N12464,R6);
not not4656(N12477,R6);
not not4657(N12489,R5);
not not4658(N12490,R6);
not not4659(N12503,R6);
not not4660(N12516,R6);
not not4661(N12529,R6);
not not4662(N12541,R6);
not not4663(N12542,R7);
not not4664(N12555,R6);
not not4665(N12567,R6);
not not4666(N12568,R7);
not not4667(N12580,R6);
not not4668(N12581,R7);
not not4669(N12594,R7);
not not4670(N12607,R7);
not not4671(N12619,R6);
not not4672(N12620,R7);
not not4673(N12633,R7);
not not4674(N12646,R7);
not not4675(N12659,R6);
not not4676(N12672,R7);
not not4677(N12683,R6);
not not4678(N12684,R7);
not not4679(N12695,R6);
not not4680(N12696,R7);
not not4681(N12708,R7);
not not4682(N12720,R4);
not not4683(N12732,R7);
not not4684(N12744,R5);
not not4685(N12755,R6);
not not4686(N12756,R7);
not not4687(N12767,R6);
not not4688(N12768,R7);
not not4689(N12780,R5);
not not4690(N12792,R6);
not not4691(N12804,R6);
not not4692(N12852,R7);
not not4693(N12864,R7);
not not4694(N12875,R6);
not not4695(N12876,R7);
not not4696(N12887,R6);
not not4697(N12888,R7);
not not4698(N12900,R6);
not not4699(N12923,R6);
not not4700(N12924,R7);
not not4701(N12935,R6);
not not4702(N12936,R7);
not not4703(N12948,R7);
not not4704(N12960,R7);
not not4705(N12971,R6);
not not4706(N12972,R7);
not not4707(N12984,R6);
not not4708(N12995,R5);
not not4709(N12996,R7);
not not4710(N13032,R6);
not not4711(N13044,R7);
not not4712(N13080,R6);
not not4713(N13092,R7);
not not4714(N13104,R7);
not not4715(N13115,R6);
not not4716(N13116,R7);
not not4717(N13128,R7);
not not4718(N13140,R7);
not not4719(N13152,R6);
not not4720(N13164,R6);
not not4721(N13176,R6);
not not4722(N13188,R7);
not not4723(N13200,R6);
not not4724(N13224,R6);
not not4725(N13236,R7);
not not4726(N13247,R6);
not not4727(N13248,R7);
not not4728(N13284,R6);
not not4729(N13295,R6);
not not4730(N13296,R7);
not not4731(N13308,R7);
not not4732(N13319,R6);
not not4733(N13320,R7);
not not4734(N13332,R6);
not not4735(N13344,R6);
not not4736(N13356,R7);
not not4737(N13380,R6);
not not4738(N13392,R6);
not not4739(N13402,R6);
not not4740(N13403,R7);
not not4741(N13413,R6);
not not4742(N13414,R7);
not not4743(N13425,R7);
not not4744(N13446,R6);
not not4745(N13447,R7);
not not4746(N13480,R6);
not not4747(N13491,R7);
not not4748(N13502,R7);
not not4749(N13513,R7);
not not4750(N13557,R6);
not not4751(N13568,R6);
not not4752(N13601,R7);
not not4753(N13623,R7);
not not4754(N13644,R5);
not not4755(N13645,R6);
not not4756(N13656,R7);
not not4757(N13667,R7);
not not4758(N13677,R6);
not not4759(N13678,R7);
not not4760(N13688,R6);
not not4761(N13689,R7);
not not4762(N13700,R5);
not not4763(N13744,R6);
not not4764(N13755,R7);
not not4765(N13777,R5);
not not4766(N13788,R5);
not not4767(N13799,R6);
not not4768(N13810,R6);
not not4769(N13821,R6);
not not4770(N13832,R6);
not not4771(N13843,R6);
not not4772(N13854,R7);
not not4773(N13865,R6);
not not4774(N13887,R5);
not not4775(N13897,R6);
not not4776(N13898,R7);
not not4777(N13920,R6);
not not4778(N13931,R6);
not not4779(N13952,R6);
not not4780(N13953,R7);
not not4781(N13963,R7);
not not4782(N13972,R5);
not not4783(N13973,R6);
not not4784(N14042,R5);
not not4785(N14043,R6);
not not4786(N14063,R6);
not not4787(N14093,R7);
not not4788(N14103,R5);
not not4789(N14112,R6);
not not4790(N14113,R7);
not not4791(N14149,R7);
not not4792(N14167,R7);
not not4793(N14176,R7);
not not4794(N14194,R6);
not not4795(N15155,in0);
not not4796(N15156,in2);
not not4797(N15157,R1);
not not4798(N15158,R2);
not not4799(N15159,R3);
not not4800(N15173,in2);
not not4801(N15174,R0);
not not4802(N15175,R1);
not not4803(N15176,R2);
not not4804(N15177,R3);
not not4805(N15190,in2);
not not4806(N15191,R0);
not not4807(N15192,R1);
not not4808(N15193,R2);
not not4809(N15194,R3);
not not4810(N15207,in0);
not not4811(N15208,in2);
not not4812(N15209,R1);
not not4813(N15223,R0);
not not4814(N15224,R1);
not not4815(N15225,R2);
not not4816(N15239,in0);
not not4817(N15240,R1);
not not4818(N15241,R3);
not not4819(N15255,in0);
not not4820(N15256,in1);
not not4821(N15257,R0);
not not4822(N15258,R1);
not not4823(N15271,in0);
not not4824(N15272,in2);
not not4825(N15273,R0);
not not4826(N15274,R1);
not not4827(N15287,in0);
not not4828(N15288,in2);
not not4829(N15289,R0);
not not4830(N15290,R1);
not not4831(N15291,R2);
not not4832(N15303,in0);
not not4833(N15304,in1);
not not4834(N15305,in2);
not not4835(N15306,R1);
not not4836(N15307,R2);
not not4837(N15319,in0);
not not4838(N15320,in1);
not not4839(N15321,in2);
not not4840(N15322,R0);
not not4841(N15323,R2);
not not4842(N15335,in0);
not not4843(N15336,in1);
not not4844(N15337,R0);
not not4845(N15338,R1);
not not4846(N15339,R2);
not not4847(N15351,in0);
not not4848(N15352,in1);
not not4849(N15353,R1);
not not4850(N15354,R2);
not not4851(N15355,R3);
not not4852(N15366,R0);
not not4853(N15367,R2);
not not4854(N15381,in0);
not not4855(N15382,R0);
not not4856(N15383,R1);
not not4857(N15384,R3);
not not4858(N15396,in0);
not not4859(N15397,in1);
not not4860(N15398,R0);
not not4861(N15399,R1);
not not4862(N15400,R3);
not not4863(N15411,R1);
not not4864(N15412,R2);
not not4865(N15413,R3);
not not4866(N15426,in0);
not not4867(N15427,in2);
not not4868(N15428,R1);
not not4869(N15429,R2);
not not4870(N15441,in0);
not not4871(N15442,R0);
not not4872(N15443,R1);
not not4873(N15456,in0);
not not4874(N15457,in1);
not not4875(N15458,R1);
not not4876(N15459,R3);
not not4877(N15471,in0);
not not4878(N15472,in1);
not not4879(N15473,in2);
not not4880(N15474,R0);
not not4881(N15486,in0);
not not4882(N15487,in2);
not not4883(N15488,R3);
not not4884(N15501,in0);
not not4885(N15502,in1);
not not4886(N15503,R1);
not not4887(N15516,in0);
not not4888(N15517,in2);
not not4889(N15518,R0);
not not4890(N15531,in0);
not not4891(N15532,R0);
not not4892(N15533,R2);
not not4893(N15546,in0);
not not4894(N15547,in2);
not not4895(N15548,R0);
not not4896(N15549,R1);
not not4897(N15561,R1);
not not4898(N15575,in1);
not not4899(N15576,R0);
not not4900(N15577,R1);
not not4901(N15589,in1);
not not4902(N15590,in2);
not not4903(N15591,R3);
not not4904(N15603,in0);
not not4905(N15604,in2);
not not4906(N15617,in0);
not not4907(N15618,in1);
not not4908(N15619,in2);
not not4909(N15620,R1);
not not4910(N15631,in0);
not not4911(N15632,in2);
not not4912(N15633,R1);
not not4913(N15645,in0);
not not4914(N15646,R1);
not not4915(N15659,R0);
not not4916(N15660,R1);
not not4917(N15661,R2);
not not4918(N15673,in1);
not not4919(N15674,in2);
not not4920(N15675,R2);
not not4921(N15687,in0);
not not4922(N15688,in1);
not not4923(N15689,R3);
not not4924(N15701,in0);
not not4925(N15702,in2);
not not4926(N15703,R0);
not not4927(N15715,in0);
not not4928(N15716,in1);
not not4929(N15717,in2);
not not4930(N15718,R1);
not not4931(N15719,R2);
not not4932(N15729,in1);
not not4933(N15730,R2);
not not4934(N15743,in1);
not not4935(N15744,in2);
not not4936(N15745,R0);
not not4937(N15746,R1);
not not4938(N15747,R3);
not not4939(N15757,R0);
not not4940(N15758,R1);
not not4941(N15771,in0);
not not4942(N15772,in1);
not not4943(N15773,in2);
not not4944(N15785,in1);
not not4945(N15786,R0);
not not4946(N15799,R0);
not not4947(N15800,R1);
not not4948(N15801,R2);
not not4949(N15813,R0);
not not4950(N15814,R1);
not not4951(N15815,R3);
not not4952(N15827,in1);
not not4953(N15828,in2);
not not4954(N15829,R0);
not not4955(N15830,R2);
not not4956(N15841,in0);
not not4957(N15842,in1);
not not4958(N15843,R1);
not not4959(N15855,in0);
not not4960(N15856,in1);
not not4961(N15857,in2);
not not4962(N15869,in1);
not not4963(N15870,in2);
not not4964(N15871,R1);
not not4965(N15872,R2);
not not4966(N15873,R3);
not not4967(N15883,R0);
not not4968(N15884,R3);
not not4969(N15897,in1);
not not4970(N15898,R0);
not not4971(N15899,R1);
not not4972(N15900,R3);
not not4973(N15911,R1);
not not4974(N15912,R2);
not not4975(N15925,in0);
not not4976(N15926,R1);
not not4977(N15927,R2);
not not4978(N15939,R0);
not not4979(N15940,R2);
not not4980(N15953,in1);
not not4981(N15954,R0);
not not4982(N15955,R1);
not not4983(N15956,R2);
not not4984(N15967,in1);
not not4985(N15968,R1);
not not4986(N15969,R2);
not not4987(N15981,in0);
not not4988(N15982,R1);
not not4989(N15983,R2);
not not4990(N15995,in0);
not not4991(N15996,in2);
not not4992(N15997,R0);
not not4993(N15998,R1);
not not4994(N16009,in2);
not not4995(N16010,R0);
not not4996(N16011,R1);
not not4997(N16012,R3);
not not4998(N16023,in1);
not not4999(N16024,R1);
not not5000(N16025,R3);
not not5001(N16037,in0);
not not5002(N16038,in1);
not not5003(N16039,R1);
not not5004(N16040,R2);
not not5005(N16051,in0);
not not5006(N16052,in2);
not not5007(N16053,R1);
not not5008(N16054,R2);
not not5009(N16065,in2);
not not5010(N16066,R0);
not not5011(N16067,R1);
not not5012(N16079,R0);
not not5013(N16080,R1);
not not5014(N16081,R2);
not not5015(N16093,in0);
not not5016(N16094,in1);
not not5017(N16095,R2);
not not5018(N16107,in2);
not not5019(N16108,R1);
not not5020(N16120,in2);
not not5021(N16121,R3);
not not5022(N16133,in0);
not not5023(N16134,in1);
not not5024(N16135,R0);
not not5025(N16146,in0);
not not5026(N16147,in2);
not not5027(N16148,R0);
not not5028(N16159,R0);
not not5029(N16160,R3);
not not5030(N16172,in0);
not not5031(N16173,in1);
not not5032(N16174,in2);
not not5033(N16185,in1);
not not5034(N16186,R2);
not not5035(N16198,in1);
not not5036(N16199,in2);
not not5037(N16200,R0);
not not5038(N16211,R0);
not not5039(N16212,R3);
not not5040(N16224,in2);
not not5041(N16225,R3);
not not5042(N16237,R0);
not not5043(N16238,R1);
not not5044(N16250,in0);
not not5045(N16251,in2);
not not5046(N16252,R2);
not not5047(N16263,in0);
not not5048(N16264,in2);
not not5049(N16276,in0);
not not5050(N16277,in2);
not not5051(N16278,R0);
not not5052(N16289,in2);
not not5053(N16302,in0);
not not5054(N16303,R0);
not not5055(N16304,R1);
not not5056(N16315,in2);
not not5057(N16316,R2);
not not5058(N16328,in1);
not not5059(N16329,in2);
not not5060(N16330,R1);
not not5061(N16331,R2);
not not5062(N16341,in1);
not not5063(N16342,in2);
not not5064(N16343,R0);
not not5065(N16344,R1);
not not5066(N16354,in0);
not not5067(N16355,in1);
not not5068(N16356,R0);
not not5069(N16357,R1);
not not5070(N16367,R2);
not not5071(N16380,in1);
not not5072(N16381,R0);
not not5073(N16382,R2);
not not5074(N16393,in0);
not not5075(N16394,R1);
not not5076(N16395,R3);
not not5077(N16406,in1);
not not5078(N16407,R0);
not not5079(N16408,R1);
not not5080(N16419,R1);
not not5081(N16431,in0);
not not5082(N16432,R1);
not not5083(N16443,R1);
not not5084(N16455,in0);
not not5085(N16467,R0);
not not5086(N16468,R1);
not not5087(N16479,R3);
not not5088(N16491,R0);
not not5089(N16503,in0);
not not5090(N16504,R0);
not not5091(N16515,in2);
not not5092(N16516,R1);
not not5093(N16527,R1);
not not5094(N16528,R3);
not not5095(N16539,in0);
not not5096(N16540,R1);
not not5097(N16541,R2);
not not5098(N16551,R1);
not not5099(N16552,R2);
not not5100(N16563,in1);
not not5101(N16564,R1);
not not5102(N16575,in0);
not not5103(N16576,in1);
not not5104(N16587,in1);
not not5105(N16588,R1);
not not5106(N16589,R2);
not not5107(N16599,in2);
not not5108(N16600,R1);
not not5109(N16601,R2);
not not5110(N16611,in0);
not not5111(N16612,R1);
not not5112(N16613,R2);
not not5113(N16623,in0);
not not5114(N16624,in1);
not not5115(N16635,in0);
not not5116(N16636,in1);
not not5117(N16637,R0);
not not5118(N16647,R0);
not not5119(N16659,in0);
not not5120(N16660,R0);
not not5121(N16661,R3);
not not5122(N16671,in2);
not not5123(N16672,R0);
not not5124(N16683,in1);
not not5125(N16684,R0);
not not5126(N16695,in1);
not not5127(N16707,R1);
not not5128(N16719,R1);
not not5129(N16720,R2);
not not5130(N16721,R3);
not not5131(N16731,in2);
not not5132(N16732,R1);
not not5133(N16733,R3);
not not5134(N16743,in0);
not not5135(N16744,R2);
not not5136(N16755,R1);
not not5137(N16756,R2);
not not5138(N16767,R1);
not not5139(N16768,R2);
not not5140(N16779,in0);
not not5141(N16780,R1);
not not5142(N16791,in2);
not not5143(N16792,R1);
not not5144(N16803,R0);
not not5145(N16804,R1);
not not5146(N16815,R2);
not not5147(N16827,in2);
not not5148(N16839,R2);
not not5149(N16851,R0);
not not5150(N16852,R1);
not not5151(N16863,in1);
not not5152(N16864,R3);
not not5153(N16875,in2);
not not5154(N16876,R3);
not not5155(N16887,in0);
not not5156(N16888,in2);
not not5157(N16899,R0);
not not5158(N16900,R1);
not not5159(N16910,R0);
not not5160(N16921,in0);
not not5161(N16932,R1);
not not5162(N16943,in2);
not not5163(N16944,R1);
not not5164(N16964,R0);
not not5165(N16984,R2);
not not5166(N17004,in2);
not not5167(N17014,in0);
not not5168(N17033,in0);
not not5169(N17034,R0);
not not5170(N17035,R2);
not not5171(N17036,R3);
not not5172(N17037,R4);
not not5173(N17038,R5);
not not5174(N17049,in1);
not not5175(N17050,in2);
not not5176(N17051,R0);
not not5177(N17052,R2);
not not5178(N17053,R4);
not not5179(N17054,R5);
not not5180(N17065,in0);
not not5181(N17066,in2);
not not5182(N17067,R0);
not not5183(N17068,R3);
not not5184(N17069,R4);
not not5185(N17070,R5);
not not5186(N17080,in2);
not not5187(N17081,R1);
not not5188(N17082,R2);
not not5189(N17083,R3);
not not5190(N17084,R4);
not not5191(N17085,R5);
not not5192(N17095,in0);
not not5193(N17096,R0);
not not5194(N17097,R1);
not not5195(N17098,R2);
not not5196(N17099,R3);
not not5197(N17110,R0);
not not5198(N17111,R1);
not not5199(N17112,R3);
not not5200(N17113,R4);
not not5201(N17114,R5);
not not5202(N17125,in1);
not not5203(N17126,in2);
not not5204(N17127,R1);
not not5205(N17128,R2);
not not5206(N17129,R3);
not not5207(N17130,R4);
not not5208(N17140,in1);
not not5209(N17141,R1);
not not5210(N17142,R2);
not not5211(N17143,R4);
not not5212(N17144,R5);
not not5213(N17155,in0);
not not5214(N17156,in1);
not not5215(N17157,in2);
not not5216(N17158,R0);
not not5217(N17159,R3);
not not5218(N17160,R4);
not not5219(N17170,in0);
not not5220(N17171,in1);
not not5221(N17172,R2);
not not5222(N17173,R3);
not not5223(N17174,R4);
not not5224(N17175,R5);
not not5225(N17185,in0);
not not5226(N17186,in1);
not not5227(N17187,R0);
not not5228(N17188,R1);
not not5229(N17189,R2);
not not5230(N17190,R3);
not not5231(N17200,in1);
not not5232(N17201,in2);
not not5233(N17202,R0);
not not5234(N17203,R1);
not not5235(N17204,R2);
not not5236(N17205,R5);
not not5237(N17215,in0);
not not5238(N17216,in1);
not not5239(N17217,in2);
not not5240(N17218,R3);
not not5241(N17219,R5);
not not5242(N17230,in0);
not not5243(N17231,R2);
not not5244(N17232,R3);
not not5245(N17233,R4);
not not5246(N17234,R5);
not not5247(N17245,in0);
not not5248(N17246,in2);
not not5249(N17247,R2);
not not5250(N17248,R3);
not not5251(N17249,R4);
not not5252(N17250,R5);
not not5253(N17260,in0);
not not5254(N17261,in1);
not not5255(N17262,R0);
not not5256(N17263,R1);
not not5257(N17264,R3);
not not5258(N17265,R4);
not not5259(N17275,in0);
not not5260(N17276,in1);
not not5261(N17277,in2);
not not5262(N17278,R1);
not not5263(N17279,R3);
not not5264(N17280,R4);
not not5265(N17290,in1);
not not5266(N17291,in2);
not not5267(N17292,R1);
not not5268(N17293,R2);
not not5269(N17294,R4);
not not5270(N17295,R5);
not not5271(N17305,in2);
not not5272(N17306,R0);
not not5273(N17307,R2);
not not5274(N17308,R5);
not not5275(N17319,R1);
not not5276(N17320,R2);
not not5277(N17321,R3);
not not5278(N17322,R4);
not not5279(N17323,R5);
not not5280(N17333,in1);
not not5281(N17334,R1);
not not5282(N17335,R3);
not not5283(N17336,R5);
not not5284(N17347,R1);
not not5285(N17348,R2);
not not5286(N17349,R3);
not not5287(N17350,R4);
not not5288(N17361,in1);
not not5289(N17362,R0);
not not5290(N17363,R4);
not not5291(N17364,R5);
not not5292(N17375,in1);
not not5293(N17376,R1);
not not5294(N17377,R4);
not not5295(N17378,R5);
not not5296(N17389,in1);
not not5297(N17390,R0);
not not5298(N17391,R1);
not not5299(N17392,R4);
not not5300(N17393,R5);
not not5301(N17403,in2);
not not5302(N17404,R0);
not not5303(N17405,R1);
not not5304(N17406,R4);
not not5305(N17407,R5);
not not5306(N17417,in0);
not not5307(N17418,in1);
not not5308(N17419,in2);
not not5309(N17420,R0);
not not5310(N17421,R1);
not not5311(N17422,R2);
not not5312(N17431,in2);
not not5313(N17432,R1);
not not5314(N17433,R2);
not not5315(N17434,R4);
not not5316(N17445,in1);
not not5317(N17446,R0);
not not5318(N17447,R1);
not not5319(N17448,R4);
not not5320(N17459,in2);
not not5321(N17460,R0);
not not5322(N17461,R1);
not not5323(N17462,R2);
not not5324(N17463,R3);
not not5325(N17473,in0);
not not5326(N17474,in1);
not not5327(N17475,R1);
not not5328(N17476,R3);
not not5329(N17477,R4);
not not5330(N17478,R5);
not not5331(N17487,in1);
not not5332(N17488,R0);
not not5333(N17489,R1);
not not5334(N17490,R2);
not not5335(N17491,R4);
not not5336(N17492,R5);
not not5337(N17501,in0);
not not5338(N17502,R0);
not not5339(N17503,R1);
not not5340(N17504,R2);
not not5341(N17515,in0);
not not5342(N17516,in2);
not not5343(N17517,R1);
not not5344(N17518,R5);
not not5345(N17529,in0);
not not5346(N17530,in1);
not not5347(N17531,R0);
not not5348(N17532,R2);
not not5349(N17533,R4);
not not5350(N17543,in0);
not not5351(N17544,in1);
not not5352(N17545,in2);
not not5353(N17546,R1);
not not5354(N17547,R5);
not not5355(N17557,in0);
not not5356(N17558,in1);
not not5357(N17559,R3);
not not5358(N17560,R4);
not not5359(N17571,in1);
not not5360(N17572,R0);
not not5361(N17573,R1);
not not5362(N17574,R2);
not not5363(N17575,R4);
not not5364(N17585,in0);
not not5365(N17586,R0);
not not5366(N17587,R1);
not not5367(N17588,R2);
not not5368(N17589,R4);
not not5369(N17599,in0);
not not5370(N17600,in2);
not not5371(N17601,R0);
not not5372(N17602,R1);
not not5373(N17603,R2);
not not5374(N17613,in1);
not not5375(N17614,R0);
not not5376(N17615,R3);
not not5377(N17616,R5);
not not5378(N17627,in0);
not not5379(N17628,in1);
not not5380(N17629,R3);
not not5381(N17630,R4);
not not5382(N17631,R5);
not not5383(N17641,in2);
not not5384(N17642,R0);
not not5385(N17643,R1);
not not5386(N17644,R4);
not not5387(N17655,in0);
not not5388(N17656,in2);
not not5389(N17657,R1);
not not5390(N17658,R4);
not not5391(N17669,in0);
not not5392(N17670,R0);
not not5393(N17671,R1);
not not5394(N17672,R4);
not not5395(N17673,R5);
not not5396(N17683,in0);
not not5397(N17684,in2);
not not5398(N17685,R0);
not not5399(N17686,R3);
not not5400(N17687,R4);
not not5401(N17697,R1);
not not5402(N17698,R2);
not not5403(N17699,R3);
not not5404(N17700,R4);
not not5405(N17701,R5);
not not5406(N17711,R0);
not not5407(N17712,R1);
not not5408(N17713,R2);
not not5409(N17714,R3);
not not5410(N17725,in0);
not not5411(N17726,in1);
not not5412(N17727,in2);
not not5413(N17728,R1);
not not5414(N17739,in1);
not not5415(N17740,R0);
not not5416(N17741,R1);
not not5417(N17742,R2);
not not5418(N17743,R5);
not not5419(N17753,in2);
not not5420(N17754,R0);
not not5421(N17755,R3);
not not5422(N17756,R5);
not not5423(N17767,in1);
not not5424(N17768,R0);
not not5425(N17769,R1);
not not5426(N17770,R4);
not not5427(N17780,R2);
not not5428(N17781,R3);
not not5429(N17782,R4);
not not5430(N17783,R5);
not not5431(N17793,R0);
not not5432(N17794,R1);
not not5433(N17795,R4);
not not5434(N17796,R5);
not not5435(N17806,in1);
not not5436(N17807,R3);
not not5437(N17808,R4);
not not5438(N17819,in2);
not not5439(N17820,R1);
not not5440(N17821,R3);
not not5441(N17822,R4);
not not5442(N17832,in2);
not not5443(N17833,R1);
not not5444(N17834,R2);
not not5445(N17835,R3);
not not5446(N17845,R0);
not not5447(N17846,R3);
not not5448(N17847,R4);
not not5449(N17858,R0);
not not5450(N17859,R1);
not not5451(N17860,R3);
not not5452(N17861,R4);
not not5453(N17871,in2);
not not5454(N17872,R1);
not not5455(N17873,R4);
not not5456(N17884,in1);
not not5457(N17885,R1);
not not5458(N17886,R3);
not not5459(N17887,R4);
not not5460(N17897,R0);
not not5461(N17898,R4);
not not5462(N17899,R5);
not not5463(N17910,in0);
not not5464(N17911,in1);
not not5465(N17912,R0);
not not5466(N17913,R4);
not not5467(N17923,R1);
not not5468(N17924,R2);
not not5469(N17925,R3);
not not5470(N17926,R5);
not not5471(N17936,in2);
not not5472(N17937,R1);
not not5473(N17938,R2);
not not5474(N17939,R3);
not not5475(N17949,in2);
not not5476(N17950,R0);
not not5477(N17951,R3);
not not5478(N17952,R5);
not not5479(N17962,R0);
not not5480(N17963,R1);
not not5481(N17964,R4);
not not5482(N17965,R5);
not not5483(N17975,in0);
not not5484(N17976,in2);
not not5485(N17977,R1);
not not5486(N17978,R2);
not not5487(N17988,in1);
not not5488(N17989,R0);
not not5489(N17990,R1);
not not5490(N17991,R2);
not not5491(N17992,R4);
not not5492(N18001,in2);
not not5493(N18002,R0);
not not5494(N18003,R3);
not not5495(N18004,R4);
not not5496(N18005,R5);
not not5497(N18014,in0);
not not5498(N18015,in2);
not not5499(N18016,R1);
not not5500(N18017,R4);
not not5501(N18027,in1);
not not5502(N18028,in2);
not not5503(N18029,R1);
not not5504(N18040,in1);
not not5505(N18041,R1);
not not5506(N18042,R3);
not not5507(N18053,in0);
not not5508(N18054,R1);
not not5509(N18055,R3);
not not5510(N18066,in1);
not not5511(N18067,R1);
not not5512(N18068,R2);
not not5513(N18069,R3);
not not5514(N18070,R4);
not not5515(N18079,in0);
not not5516(N18080,in2);
not not5517(N18081,R1);
not not5518(N18082,R2);
not not5519(N18092,in0);
not not5520(N18093,in1);
not not5521(N18094,R1);
not not5522(N18095,R4);
not not5523(N18105,in2);
not not5524(N18106,R0);
not not5525(N18107,R1);
not not5526(N18118,in2);
not not5527(N18119,R1);
not not5528(N18120,R5);
not not5529(N18131,in2);
not not5530(N18132,R1);
not not5531(N18133,R3);
not not5532(N18144,in0);
not not5533(N18145,R1);
not not5534(N18146,R3);
not not5535(N18157,in0);
not not5536(N18158,in2);
not not5537(N18159,R1);
not not5538(N18160,R3);
not not5539(N18161,R4);
not not5540(N18170,in1);
not not5541(N18171,R2);
not not5542(N18172,R3);
not not5543(N18183,in1);
not not5544(N18184,R2);
not not5545(N18185,R4);
not not5546(N18186,R5);
not not5547(N18196,R0);
not not5548(N18197,R1);
not not5549(N18198,R2);
not not5550(N18199,R5);
not not5551(N18209,R0);
not not5552(N18210,R1);
not not5553(N18211,R2);
not not5554(N18212,R5);
not not5555(N18222,R0);
not not5556(N18223,R2);
not not5557(N18224,R4);
not not5558(N18235,in0);
not not5559(N18236,in2);
not not5560(N18237,R0);
not not5561(N18238,R4);
not not5562(N18248,in2);
not not5563(N18249,R0);
not not5564(N18250,R1);
not not5565(N18251,R2);
not not5566(N18261,in2);
not not5567(N18262,R0);
not not5568(N18263,R1);
not not5569(N18264,R4);
not not5570(N18274,in0);
not not5571(N18275,in1);
not not5572(N18276,in2);
not not5573(N18277,R2);
not not5574(N18287,in1);
not not5575(N18288,in2);
not not5576(N18289,R1);
not not5577(N18290,R4);
not not5578(N18300,in1);
not not5579(N18301,in2);
not not5580(N18302,R1);
not not5581(N18303,R4);
not not5582(N18313,in2);
not not5583(N18314,R1);
not not5584(N18315,R4);
not not5585(N18316,R5);
not not5586(N18326,in1);
not not5587(N18327,R1);
not not5588(N18328,R4);
not not5589(N18329,R5);
not not5590(N18339,in0);
not not5591(N18340,R2);
not not5592(N18341,R4);
not not5593(N18352,in1);
not not5594(N18353,R4);
not not5595(N18354,R5);
not not5596(N18365,in2);
not not5597(N18366,R2);
not not5598(N18367,R5);
not not5599(N18378,in0);
not not5600(N18379,in1);
not not5601(N18380,R0);
not not5602(N18381,R1);
not not5603(N18382,R4);
not not5604(N18391,in1);
not not5605(N18392,R1);
not not5606(N18393,R4);
not not5607(N18404,in0);
not not5608(N18405,in1);
not not5609(N18406,R0);
not not5610(N18407,R3);
not not5611(N18417,in2);
not not5612(N18418,R0);
not not5613(N18419,R1);
not not5614(N18420,R4);
not not5615(N18430,in0);
not not5616(N18431,in2);
not not5617(N18432,R4);
not not5618(N18443,in1);
not not5619(N18444,R0);
not not5620(N18445,R3);
not not5621(N18446,R4);
not not5622(N18456,R1);
not not5623(N18457,R2);
not not5624(N18458,R4);
not not5625(N18469,in0);
not not5626(N18470,R1);
not not5627(N18471,R4);
not not5628(N18482,R0);
not not5629(N18483,R2);
not not5630(N18484,R5);
not not5631(N18495,R0);
not not5632(N18496,R1);
not not5633(N18497,R2);
not not5634(N18498,R4);
not not5635(N18499,R5);
not not5636(N18508,in0);
not not5637(N18509,in1);
not not5638(N18510,R1);
not not5639(N18511,R2);
not not5640(N18521,in1);
not not5641(N18522,R1);
not not5642(N18523,R2);
not not5643(N18534,in0);
not not5644(N18535,in1);
not not5645(N18536,R0);
not not5646(N18537,R2);
not not5647(N18547,in1);
not not5648(N18548,R1);
not not5649(N18549,R3);
not not5650(N18550,R4);
not not5651(N18560,in2);
not not5652(N18561,R1);
not not5653(N18562,R3);
not not5654(N18563,R4);
not not5655(N18573,in1);
not not5656(N18574,in2);
not not5657(N18575,R1);
not not5658(N18576,R2);
not not5659(N18577,R4);
not not5660(N18586,in0);
not not5661(N18587,in1);
not not5662(N18588,in2);
not not5663(N18589,R1);
not not5664(N18599,in2);
not not5665(N18600,R3);
not not5666(N18611,in2);
not not5667(N18612,R4);
not not5668(N18613,R5);
not not5669(N18623,in2);
not not5670(N18624,R0);
not not5671(N18635,R3);
not not5672(N18636,R4);
not not5673(N18647,in1);
not not5674(N18648,R0);
not not5675(N18649,R4);
not not5676(N18659,in1);
not not5677(N18660,in2);
not not5678(N18661,R5);
not not5679(N18671,R0);
not not5680(N18672,R3);
not not5681(N18683,R2);
not not5682(N18684,R3);
not not5683(N18695,in0);
not not5684(N18696,R3);
not not5685(N18697,R4);
not not5686(N18707,in0);
not not5687(N18708,in1);
not not5688(N18709,R0);
not not5689(N18710,R2);
not not5690(N18719,in1);
not not5691(N18720,R3);
not not5692(N18721,R5);
not not5693(N18731,in2);
not not5694(N18732,R2);
not not5695(N18733,R4);
not not5696(N18743,in1);
not not5697(N18744,R4);
not not5698(N18745,R5);
not not5699(N18755,in1);
not not5700(N18756,R1);
not not5701(N18757,R3);
not not5702(N18767,in0);
not not5703(N18768,R2);
not not5704(N18779,R2);
not not5705(N18780,R3);
not not5706(N18781,R5);
not not5707(N18791,in1);
not not5708(N18792,R3);
not not5709(N18803,R1);
not not5710(N18804,R5);
not not5711(N18815,R1);
not not5712(N18816,R5);
not not5713(N18827,in1);
not not5714(N18828,in2);
not not5715(N18839,in2);
not not5716(N18840,R2);
not not5717(N18841,R4);
not not5718(N18851,in2);
not not5719(N18852,R0);
not not5720(N18853,R1);
not not5721(N18854,R2);
not not5722(N18863,in1);
not not5723(N18864,R0);
not not5724(N18865,R5);
not not5725(N18875,in2);
not not5726(N18876,R0);
not not5727(N18877,R5);
not not5728(N18887,in1);
not not5729(N18888,R1);
not not5730(N18889,R3);
not not5731(N18890,R4);
not not5732(N18899,R0);
not not5733(N18900,R1);
not not5734(N18901,R3);
not not5735(N18911,in2);
not not5736(N18912,R0);
not not5737(N18913,R2);
not not5738(N18923,R3);
not not5739(N18924,R4);
not not5740(N18925,R5);
not not5741(N18935,in1);
not not5742(N18936,in2);
not not5743(N18937,R3);
not not5744(N18947,R0);
not not5745(N18948,R1);
not not5746(N18949,R3);
not not5747(N18959,in1);
not not5748(N18960,R2);
not not5749(N18961,R4);
not not5750(N18971,in0);
not not5751(N18972,in1);
not not5752(N18973,R4);
not not5753(N18983,R0);
not not5754(N18984,R2);
not not5755(N18985,R4);
not not5756(N18995,in0);
not not5757(N18996,in2);
not not5758(N18997,R0);
not not5759(N18998,R5);
not not5760(N19007,R1);
not not5761(N19008,R2);
not not5762(N19009,R3);
not not5763(N19010,R4);
not not5764(N19019,in2);
not not5765(N19020,R4);
not not5766(N19031,in0);
not not5767(N19032,R0);
not not5768(N19033,R3);
not not5769(N19034,R5);
not not5770(N19043,R2);
not not5771(N19044,R3);
not not5772(N19055,in2);
not not5773(N19056,R3);
not not5774(N19057,R4);
not not5775(N19067,in1);
not not5776(N19068,R0);
not not5777(N19069,R1);
not not5778(N19070,R2);
not not5779(N19079,in0);
not not5780(N19080,in1);
not not5781(N19081,R3);
not not5782(N19091,in1);
not not5783(N19092,R1);
not not5784(N19093,R4);
not not5785(N19103,in2);
not not5786(N19104,R1);
not not5787(N19105,R4);
not not5788(N19115,R2);
not not5789(N19116,R5);
not not5790(N19127,R0);
not not5791(N19128,R1);
not not5792(N19129,R4);
not not5793(N19139,in2);
not not5794(N19140,R2);
not not5795(N19141,R4);
not not5796(N19151,in0);
not not5797(N19152,R2);
not not5798(N19163,R0);
not not5799(N19164,R4);
not not5800(N19174,in0);
not not5801(N19175,in2);
not not5802(N19185,in0);
not not5803(N19186,R1);
not not5804(N19187,R5);
not not5805(N19196,R3);
not not5806(N19197,R4);
not not5807(N19207,R1);
not not5808(N19208,R3);
not not5809(N19218,in1);
not not5810(N19219,R4);
not not5811(N19229,in1);
not not5812(N19230,R1);
not not5813(N19240,in1);
not not5814(N19241,R0);
not not5815(N19251,in0);
not not5816(N19252,in1);
not not5817(N19253,R3);
not not5818(N19262,in0);
not not5819(N19263,R0);
not not5820(N19264,R4);
not not5821(N19273,in0);
not not5822(N19274,in2);
not not5823(N19284,R2);
not not5824(N19285,R4);
not not5825(N19295,R1);
not not5826(N19296,R4);
not not5827(N19306,in0);
not not5828(N19317,R1);
not not5829(N19318,R4);
not not5830(N19328,in1);
not not5831(N19329,R3);
not not5832(N19330,R4);
not not5833(N19339,in2);
not not5834(N19340,R1);
not not5835(N19350,in0);
not not5836(N19351,R1);
not not5837(N19352,R2);
not not5838(N19361,R1);
not not5839(N19362,R3);
not not5840(N19372,in0);
not not5841(N19373,R3);
not not5842(N19374,R5);
not not5843(N19383,R0);
not not5844(N19384,R1);
not not5845(N19385,R5);
not not5846(N19394,in1);
not not5847(N19395,in2);
not not5848(N19405,in1);
not not5849(N19406,R3);
not not5850(N19407,R4);
not not5851(N19416,in1);
not not5852(N19417,in2);
not not5853(N19418,R0);
not not5854(N19427,in1);
not not5855(N19428,R0);
not not5856(N19438,in2);
not not5857(N19439,R2);
not not5858(N19449,in1);
not not5859(N19450,R1);
not not5860(N19460,R1);
not not5861(N19461,R4);
not not5862(N19471,in0);
not not5863(N19472,R2);
not not5864(N19482,R1);
not not5865(N19483,R3);
not not5866(N19493,R1);
not not5867(N19494,R3);
not not5868(N19504,in0);
not not5869(N19505,R0);
not not5870(N19515,in1);
not not5871(N19516,in2);
not not5872(N19517,R3);
not not5873(N19526,in2);
not not5874(N19527,R1);
not not5875(N19537,R0);
not not5876(N19538,R2);
not not5877(N19548,R3);
not not5878(N19549,R5);
not not5879(N19559,R0);
not not5880(N19560,R5);
not not5881(N19570,R4);
not not5882(N19581,in1);
not not5883(N19582,R2);
not not5884(N19591,in2);
not not5885(N19592,R5);
not not5886(N19601,R5);
not not5887(N19611,in1);
not not5888(N19612,R2);
not not5889(N19621,R2);
not not5890(N19622,R5);
not not5891(N19631,in1);
not not5892(N19632,R3);
not not5893(N19641,R2);
not not5894(N19642,R4);
not not5895(N19651,R0);
not not5896(N19652,R2);
not not5897(N19661,R3);
not not5898(N19671,R4);
not not5899(N19672,R5);
not not5900(N19681,in2);
not not5901(N19682,R5);
not not5902(N19691,R3);
not not5903(N19711,in0);
not not5904(N19712,R2);
not not5905(N19721,R0);
not not5906(N19731,R0);
not not5907(N19741,in1);
not not5908(N19751,in2);
not not5909(N19752,R5);
not not5910(N19761,R3);
not not5911(N19762,R4);
not not5912(N19771,in0);
not not5913(N19780,R5);
not not5914(N19789,R3);
not not5915(N19798,in1);
not not5916(N19807,in1);
not not5917(N19825,in1);
not not5918(N19834,R3);
not not5919(N19843,R2);
not not5920(N19859,in1);
not not5921(N19860,R2);
not not5922(N19861,R3);
not not5923(N19862,R4);
not not5924(N19863,R5);
not not5925(N19864,R6);
not not5926(N19865,R7);
not not5927(N19873,in1);
not not5928(N19874,R1);
not not5929(N19875,R2);
not not5930(N19876,R3);
not not5931(N19877,R4);
not not5932(N19878,R5);
not not5933(N19879,R7);
not not5934(N19887,R0);
not not5935(N19888,R2);
not not5936(N19889,R3);
not not5937(N19890,R4);
not not5938(N19891,R5);
not not5939(N19892,R6);
not not5940(N19893,R7);
not not5941(N19901,R0);
not not5942(N19902,R1);
not not5943(N19903,R2);
not not5944(N19904,R3);
not not5945(N19905,R4);
not not5946(N19906,R6);
not not5947(N19907,R7);
not not5948(N19915,in1);
not not5949(N19916,R0);
not not5950(N19917,R2);
not not5951(N19918,R3);
not not5952(N19919,R4);
not not5953(N19920,R5);
not not5954(N19921,R6);
not not5955(N19929,in1);
not not5956(N19930,R0);
not not5957(N19931,R1);
not not5958(N19932,R2);
not not5959(N19933,R6);
not not5960(N19934,R7);
not not5961(N19942,in2);
not not5962(N19943,R2);
not not5963(N19944,R3);
not not5964(N19945,R5);
not not5965(N19946,R6);
not not5966(N19947,R7);
not not5967(N19955,in0);
not not5968(N19956,in1);
not not5969(N19957,in2);
not not5970(N19958,R1);
not not5971(N19959,R6);
not not5972(N19960,R7);
not not5973(N19968,R2);
not not5974(N19969,R3);
not not5975(N19970,R4);
not not5976(N19971,R5);
not not5977(N19972,R6);
not not5978(N19980,in1);
not not5979(N19981,R1);
not not5980(N19982,R3);
not not5981(N19983,R4);
not not5982(N19984,R6);
not not5983(N19992,R0);
not not5984(N19993,R3);
not not5985(N19994,R4);
not not5986(N19995,R5);
not not5987(N19996,R6);
not not5988(N20004,in1);
not not5989(N20005,R0);
not not5990(N20006,R3);
not not5991(N20007,R6);
not not5992(N20008,R7);
not not5993(N20016,in2);
not not5994(N20017,R0);
not not5995(N20018,R2);
not not5996(N20019,R5);
not not5997(N20020,R6);
not not5998(N20028,in1);
not not5999(N20029,R0);
not not6000(N20030,R2);
not not6001(N20031,R4);
not not6002(N20032,R6);
not not6003(N20040,in2);
not not6004(N20041,R0);
not not6005(N20042,R2);
not not6006(N20043,R4);
not not6007(N20044,R6);
not not6008(N20052,in2);
not not6009(N20053,R0);
not not6010(N20054,R1);
not not6011(N20055,R3);
not not6012(N20056,R7);
not not6013(N20064,in2);
not not6014(N20065,R0);
not not6015(N20066,R3);
not not6016(N20067,R6);
not not6017(N20068,R7);
not not6018(N20076,R0);
not not6019(N20077,R1);
not not6020(N20078,R2);
not not6021(N20079,R6);
not not6022(N20080,R7);
not not6023(N20088,in1);
not not6024(N20089,R3);
not not6025(N20090,R4);
not not6026(N20091,R6);
not not6027(N20099,R1);
not not6028(N20100,R2);
not not6029(N20101,R3);
not not6030(N20102,R6);
not not6031(N20110,in1);
not not6032(N20111,R0);
not not6033(N20112,R4);
not not6034(N20113,R5);
not not6035(N20121,R1);
not not6036(N20122,R2);
not not6037(N20123,R5);
not not6038(N20124,R7);
not not6039(N20132,R1);
not not6040(N20133,R2);
not not6041(N20134,R5);
not not6042(N20135,R7);
not not6043(N20143,in1);
not not6044(N20144,R2);
not not6045(N20145,R3);
not not6046(N20146,R6);
not not6047(N20154,R1);
not not6048(N20155,R4);
not not6049(N20156,R5);
not not6050(N20157,R6);
not not6051(N20165,R1);
not not6052(N20166,R3);
not not6053(N20167,R4);
not not6054(N20168,R5);
not not6055(N20176,in1);
not not6056(N20177,in2);
not not6057(N20178,R0);
not not6058(N20179,R5);
not not6059(N20187,in2);
not not6060(N20188,R1);
not not6061(N20189,R2);
not not6062(N20190,R7);
not not6063(N20198,R3);
not not6064(N20199,R4);
not not6065(N20200,R6);
not not6066(N20201,R7);
not not6067(N20209,R0);
not not6068(N20210,R4);
not not6069(N20211,R5);
not not6070(N20212,R6);
not not6071(N20220,in1);
not not6072(N20221,R0);
not not6073(N20222,R1);
not not6074(N20223,R6);
not not6075(N20231,R0);
not not6076(N20232,R4);
not not6077(N20233,R7);
not not6078(N20241,R2);
not not6079(N20242,R5);
not not6080(N20243,R6);
not not6081(N20251,in1);
not not6082(N20252,R6);
not not6083(N20253,R7);
not not6084(N20261,R4);
not not6085(N20262,R6);
not not6086(N20263,R7);
not not6087(N20271,in1);
not not6088(N20272,R1);
not not6089(N20273,R5);
not not6090(N20281,R0);
not not6091(N20282,R1);
not not6092(N20283,R2);
not not6093(N20291,R2);
not not6094(N20292,R4);
not not6095(N20293,R5);
not not6096(N20301,in0);
not not6097(N20302,R1);
not not6098(N20303,R6);
not not6099(N20311,in2);
not not6100(N20312,R0);
not not6101(N20313,R1);
not not6102(N20321,in2);
not not6103(N20322,R1);
not not6104(N20323,R5);
not not6105(N20331,R1);
not not6106(N20332,R2);
not not6107(N20333,R7);
not not6108(N20341,R4);
not not6109(N20342,R5);
not not6110(N20350,R4);
not not6111(N20351,R7);
not not6112(N20359,R0);
not not6113(N20360,R7);
not not6114(N20368,R5);
not not6115(N20369,R6);
not not6116(N20377,R4);
not not6117(N20385,R7);
not not6118(N20393,R7);
not not6119(N20400,R6);
not not6120(N20401,R7);
not not6121(N15160,R4);
not not6122(N15161,R5);
not not6123(N15162,R6);
not not6124(N15163,R7);
not not6125(N15178,R5);
not not6126(N15179,R6);
not not6127(N15180,R7);
not not6128(N15195,R4);
not not6129(N15196,R5);
not not6130(N15197,R6);
not not6131(N15210,R4);
not not6132(N15211,R5);
not not6133(N15212,R6);
not not6134(N15213,R7);
not not6135(N15226,R4);
not not6136(N15227,R5);
not not6137(N15228,R6);
not not6138(N15229,R7);
not not6139(N15242,R4);
not not6140(N15243,R5);
not not6141(N15244,R6);
not not6142(N15245,R7);
not not6143(N15259,R3);
not not6144(N15260,R4);
not not6145(N15261,R7);
not not6146(N15275,R4);
not not6147(N15276,R5);
not not6148(N15277,R6);
not not6149(N15292,R3);
not not6150(N15293,R6);
not not6151(N15308,R3);
not not6152(N15309,R4);
not not6153(N15324,R4);
not not6154(N15325,R6);
not not6155(N15340,R4);
not not6156(N15341,R6);
not not6157(N15356,R6);
not not6158(N15368,R4);
not not6159(N15369,R5);
not not6160(N15370,R6);
not not6161(N15371,R7);
not not6162(N15385,R4);
not not6163(N15386,R6);
not not6164(N15401,R6);
not not6165(N15414,R5);
not not6166(N15415,R6);
not not6167(N15416,R7);
not not6168(N15430,R3);
not not6169(N15431,R6);
not not6170(N15444,R3);
not not6171(N15445,R4);
not not6172(N15446,R7);
not not6173(N15460,R5);
not not6174(N15461,R7);
not not6175(N15475,R6);
not not6176(N15476,R7);
not not6177(N15489,R5);
not not6178(N15490,R6);
not not6179(N15491,R7);
not not6180(N15504,R5);
not not6181(N15505,R6);
not not6182(N15506,R7);
not not6183(N15519,R4);
not not6184(N15520,R5);
not not6185(N15521,R7);
not not6186(N15534,R4);
not not6187(N15535,R5);
not not6188(N15536,R6);
not not6189(N15550,R3);
not not6190(N15551,R5);
not not6191(N15562,R4);
not not6192(N15563,R5);
not not6193(N15564,R6);
not not6194(N15565,R7);
not not6195(N15578,R6);
not not6196(N15579,R7);
not not6197(N15592,R4);
not not6198(N15593,R7);
not not6199(N15605,R3);
not not6200(N15606,R4);
not not6201(N15607,R7);
not not6202(N15621,R3);
not not6203(N15634,R4);
not not6204(N15635,R6);
not not6205(N15647,R4);
not not6206(N15648,R5);
not not6207(N15649,R6);
not not6208(N15662,R5);
not not6209(N15663,R6);
not not6210(N15676,R4);
not not6211(N15677,R7);
not not6212(N15690,R4);
not not6213(N15691,R7);
not not6214(N15704,R4);
not not6215(N15705,R7);
not not6216(N15731,R5);
not not6217(N15732,R6);
not not6218(N15733,R7);
not not6219(N15759,R3);
not not6220(N15760,R4);
not not6221(N15761,R6);
not not6222(N15774,R4);
not not6223(N15775,R6);
not not6224(N15787,R5);
not not6225(N15788,R6);
not not6226(N15789,R7);
not not6227(N15802,R4);
not not6228(N15803,R6);
not not6229(N15816,R4);
not not6230(N15817,R5);
not not6231(N15831,R4);
not not6232(N15844,R3);
not not6233(N15845,R4);
not not6234(N15858,R6);
not not6235(N15859,R7);
not not6236(N15885,R5);
not not6237(N15886,R6);
not not6238(N15887,R7);
not not6239(N15901,R7);
not not6240(N15913,R5);
not not6241(N15914,R6);
not not6242(N15915,R7);
not not6243(N15928,R3);
not not6244(N15929,R4);
not not6245(N15941,R4);
not not6246(N15942,R5);
not not6247(N15943,R7);
not not6248(N15957,R7);
not not6249(N15970,R3);
not not6250(N15971,R7);
not not6251(N15984,R3);
not not6252(N15985,R6);
not not6253(N15999,R5);
not not6254(N16013,R4);
not not6255(N16026,R5);
not not6256(N16027,R7);
not not6257(N16041,R4);
not not6258(N16055,R4);
not not6259(N16068,R4);
not not6260(N16069,R5);
not not6261(N16082,R4);
not not6262(N16083,R7);
not not6263(N16096,R4);
not not6264(N16097,R6);
not not6265(N16109,R6);
not not6266(N16110,R7);
not not6267(N16122,R6);
not not6268(N16123,R7);
not not6269(N16136,R5);
not not6270(N16149,R6);
not not6271(N16161,R4);
not not6272(N16162,R6);
not not6273(N16175,R4);
not not6274(N16187,R5);
not not6275(N16188,R7);
not not6276(N16201,R4);
not not6277(N16213,R4);
not not6278(N16214,R7);
not not6279(N16226,R4);
not not6280(N16227,R7);
not not6281(N16239,R6);
not not6282(N16240,R7);
not not6283(N16253,R5);
not not6284(N16265,R5);
not not6285(N16266,R7);
not not6286(N16279,R7);
not not6287(N16290,R5);
not not6288(N16291,R6);
not not6289(N16292,R7);
not not6290(N16305,R3);
not not6291(N16317,R3);
not not6292(N16318,R6);
not not6293(N16368,R4);
not not6294(N16369,R5);
not not6295(N16370,R7);
not not6296(N16383,R6);
not not6297(N16396,R7);
not not6298(N16409,R4);
not not6299(N16420,R6);
not not6300(N16421,R7);
not not6301(N16433,R6);
not not6302(N16444,R4);
not not6303(N16445,R6);
not not6304(N16456,R4);
not not6305(N16457,R6);
not not6306(N16469,R6);
not not6307(N16480,R4);
not not6308(N16481,R7);
not not6309(N16492,R4);
not not6310(N16493,R5);
not not6311(N16505,R5);
not not6312(N16517,R3);
not not6313(N16529,R4);
not not6314(N16553,R4);
not not6315(N16565,R4);
not not6316(N16577,R4);
not not6317(N16625,R6);
not not6318(N16648,R3);
not not6319(N16649,R5);
not not6320(N16673,R3);
not not6321(N16685,R4);
not not6322(N16696,R5);
not not6323(N16697,R7);
not not6324(N16708,R5);
not not6325(N16709,R7);
not not6326(N16745,R5);
not not6327(N16757,R5);
not not6328(N16769,R6);
not not6329(N16781,R6);
not not6330(N16793,R4);
not not6331(N16805,R3);
not not6332(N16816,R3);
not not6333(N16817,R6);
not not6334(N16828,R5);
not not6335(N16829,R6);
not not6336(N16840,R4);
not not6337(N16841,R6);
not not6338(N16853,R4);
not not6339(N16865,R7);
not not6340(N16877,R7);
not not6341(N16889,R4);
not not6342(N16911,R4);
not not6343(N16922,R4);
not not6344(N16933,R3);
not not6345(N16954,R6);
not not6346(N16974,R5);
not not6347(N16994,R6);
not not6348(N17024,R6);
not not6349(N17039,R6);
not not6350(N17040,R7);
not not6351(N17055,R6);
not not6352(N17056,R7);
not not6353(N17071,R6);
not not6354(N17086,R7);
not not6355(N17100,R6);
not not6356(N17101,R7);
not not6357(N17115,R6);
not not6358(N17116,R7);
not not6359(N17131,R6);
not not6360(N17145,R6);
not not6361(N17146,R7);
not not6362(N17161,R6);
not not6363(N17176,R6);
not not6364(N17191,R6);
not not6365(N17206,R6);
not not6366(N17220,R6);
not not6367(N17221,R7);
not not6368(N17235,R6);
not not6369(N17236,R7);
not not6370(N17251,R6);
not not6371(N17266,R6);
not not6372(N17281,R6);
not not6373(N17296,R7);
not not6374(N17309,R6);
not not6375(N17310,R7);
not not6376(N17324,R6);
not not6377(N17337,R6);
not not6378(N17338,R7);
not not6379(N17351,R6);
not not6380(N17352,R7);
not not6381(N17365,R6);
not not6382(N17366,R7);
not not6383(N17379,R6);
not not6384(N17380,R7);
not not6385(N17394,R7);
not not6386(N17408,R7);
not not6387(N17435,R6);
not not6388(N17436,R7);
not not6389(N17449,R5);
not not6390(N17450,R6);
not not6391(N17464,R6);
not not6392(N17505,R5);
not not6393(N17506,R6);
not not6394(N17519,R6);
not not6395(N17520,R7);
not not6396(N17534,R7);
not not6397(N17548,R7);
not not6398(N17561,R6);
not not6399(N17562,R7);
not not6400(N17576,R7);
not not6401(N17590,R7);
not not6402(N17604,R4);
not not6403(N17617,R6);
not not6404(N17618,R7);
not not6405(N17632,R7);
not not6406(N17645,R6);
not not6407(N17646,R7);
not not6408(N17659,R6);
not not6409(N17660,R7);
not not6410(N17674,R7);
not not6411(N17688,R6);
not not6412(N17702,R7);
not not6413(N17715,R6);
not not6414(N17716,R7);
not not6415(N17729,R5);
not not6416(N17730,R6);
not not6417(N17744,R6);
not not6418(N17757,R6);
not not6419(N17758,R7);
not not6420(N17771,R6);
not not6421(N17784,R6);
not not6422(N17797,R7);
not not6423(N17809,R5);
not not6424(N17810,R7);
not not6425(N17823,R6);
not not6426(N17836,R4);
not not6427(N17848,R5);
not not6428(N17849,R6);
not not6429(N17862,R7);
not not6430(N17874,R6);
not not6431(N17875,R7);
not not6432(N17888,R6);
not not6433(N17900,R6);
not not6434(N17901,R7);
not not6435(N17914,R6);
not not6436(N17927,R6);
not not6437(N17940,R6);
not not6438(N17953,R6);
not not6439(N17966,R6);
not not6440(N17979,R5);
not not6441(N18018,R7);
not not6442(N18030,R6);
not not6443(N18031,R7);
not not6444(N18043,R6);
not not6445(N18044,R7);
not not6446(N18056,R6);
not not6447(N18057,R7);
not not6448(N18083,R7);
not not6449(N18096,R5);
not not6450(N18108,R6);
not not6451(N18109,R7);
not not6452(N18121,R6);
not not6453(N18122,R7);
not not6454(N18134,R5);
not not6455(N18135,R7);
not not6456(N18147,R5);
not not6457(N18148,R7);
not not6458(N18173,R6);
not not6459(N18174,R7);
not not6460(N18187,R7);
not not6461(N18200,R7);
not not6462(N18213,R7);
not not6463(N18225,R6);
not not6464(N18226,R7);
not not6465(N18239,R5);
not not6466(N18252,R4);
not not6467(N18265,R6);
not not6468(N18278,R6);
not not6469(N18291,R7);
not not6470(N18304,R6);
not not6471(N18317,R7);
not not6472(N18330,R7);
not not6473(N18342,R5);
not not6474(N18343,R6);
not not6475(N18355,R6);
not not6476(N18356,R7);
not not6477(N18368,R6);
not not6478(N18369,R7);
not not6479(N18394,R6);
not not6480(N18395,R7);
not not6481(N18408,R5);
not not6482(N18421,R7);
not not6483(N18433,R6);
not not6484(N18434,R7);
not not6485(N18447,R7);
not not6486(N18459,R6);
not not6487(N18460,R7);
not not6488(N18472,R6);
not not6489(N18473,R7);
not not6490(N18485,R6);
not not6491(N18486,R7);
not not6492(N18512,R7);
not not6493(N18524,R6);
not not6494(N18525,R7);
not not6495(N18538,R6);
not not6496(N18551,R7);
not not6497(N18564,R7);
not not6498(N18590,R7);
not not6499(N18601,R5);
not not6500(N18602,R7);
not not6501(N18614,R6);
not not6502(N18625,R5);
not not6503(N18626,R6);
not not6504(N18637,R5);
not not6505(N18638,R7);
not not6506(N18650,R6);
not not6507(N18662,R7);
not not6508(N18673,R6);
not not6509(N18674,R7);
not not6510(N18685,R5);
not not6511(N18686,R6);
not not6512(N18698,R6);
not not6513(N18722,R7);
not not6514(N18734,R7);
not not6515(N18746,R7);
not not6516(N18758,R6);
not not6517(N18769,R6);
not not6518(N18770,R7);
not not6519(N18782,R6);
not not6520(N18793,R6);
not not6521(N18794,R7);
not not6522(N18805,R6);
not not6523(N18806,R7);
not not6524(N18817,R6);
not not6525(N18818,R7);
not not6526(N18829,R5);
not not6527(N18830,R6);
not not6528(N18842,R7);
not not6529(N18866,R7);
not not6530(N18878,R7);
not not6531(N18902,R7);
not not6532(N18914,R6);
not not6533(N18926,R7);
not not6534(N18938,R5);
not not6535(N18950,R6);
not not6536(N18962,R6);
not not6537(N18974,R6);
not not6538(N18986,R6);
not not6539(N19021,R5);
not not6540(N19022,R7);
not not6541(N19045,R6);
not not6542(N19046,R7);
not not6543(N19058,R6);
not not6544(N19082,R6);
not not6545(N19094,R6);
not not6546(N19106,R6);
not not6547(N19117,R6);
not not6548(N19118,R7);
not not6549(N19130,R7);
not not6550(N19142,R6);
not not6551(N19153,R4);
not not6552(N19154,R6);
not not6553(N19165,R6);
not not6554(N19176,R6);
not not6555(N19198,R6);
not not6556(N19209,R6);
not not6557(N19220,R5);
not not6558(N19231,R6);
not not6559(N19242,R5);
not not6560(N19275,R7);
not not6561(N19286,R7);
not not6562(N19297,R7);
not not6563(N19307,R5);
not not6564(N19308,R6);
not not6565(N19319,R7);
not not6566(N19341,R7);
not not6567(N19363,R5);
not not6568(N19396,R6);
not not6569(N19429,R6);
not not6570(N19440,R6);
not not6571(N19451,R7);
not not6572(N19462,R7);
not not6573(N19473,R7);
not not6574(N19484,R5);
not not6575(N19495,R5);
not not6576(N19506,R6);
not not6577(N19528,R6);
not not6578(N19539,R6);
not not6579(N19550,R6);
not not6580(N19561,R6);
not not6581(N19571,R6);
not not6582(N19572,R7);
not not6583(N19602,R7);
not not6584(N19662,R7);
not not6585(N19692,R7);
not not6586(N19701,R5);
not not6587(N19702,R6);
not not6588(N19722,R6);
not not6589(N19732,R7);
not not6590(N19742,R6);
not not6591(N19816,R7);
not not6592(N20645,in0);
not not6593(N20646,in1);
not not6594(N20660,in0);
not not6595(N20661,in1);
not not6596(N20662,in2);
not not6597(N20663,R1);
not not6598(N20664,R2);
not not6599(N20678,in0);
not not6600(N20679,in1);
not not6601(N20680,in2);
not not6602(N20681,R1);
not not6603(N20682,R2);
not not6604(N20683,R3);
not not6605(N20696,in0);
not not6606(N20697,R0);
not not6607(N20698,R1);
not not6608(N20699,R2);
not not6609(N20700,R3);
not not6610(N20713,in0);
not not6611(N20714,in1);
not not6612(N20715,R0);
not not6613(N20716,R1);
not not6614(N20717,R2);
not not6615(N20730,in0);
not not6616(N20731,in1);
not not6617(N20732,in2);
not not6618(N20733,R1);
not not6619(N20747,in0);
not not6620(N20748,in1);
not not6621(N20749,in2);
not not6622(N20750,R1);
not not6623(N20751,R2);
not not6624(N20764,in0);
not not6625(N20765,in1);
not not6626(N20766,in2);
not not6627(N20767,R0);
not not6628(N20768,R1);
not not6629(N20781,in0);
not not6630(N20782,in1);
not not6631(N20783,R1);
not not6632(N20784,R2);
not not6633(N20785,R3);
not not6634(N20798,in0);
not not6635(N20799,in1);
not not6636(N20800,R1);
not not6637(N20801,R2);
not not6638(N20802,R3);
not not6639(N20815,in0);
not not6640(N20816,in1);
not not6641(N20817,in2);
not not6642(N20818,R0);
not not6643(N20819,R1);
not not6644(N20820,R2);
not not6645(N20832,in0);
not not6646(N20833,in1);
not not6647(N20834,in2);
not not6648(N20835,R0);
not not6649(N20836,R1);
not not6650(N20837,R3);
not not6651(N20849,in0);
not not6652(N20850,in1);
not not6653(N20851,in2);
not not6654(N20852,R0);
not not6655(N20853,R1);
not not6656(N20854,R2);
not not6657(N20866,in0);
not not6658(N20867,in1);
not not6659(N20868,in2);
not not6660(N20869,R0);
not not6661(N20870,R1);
not not6662(N20871,R2);
not not6663(N20883,in0);
not not6664(N20884,in1);
not not6665(N20885,in2);
not not6666(N20886,R0);
not not6667(N20887,R1);
not not6668(N20888,R2);
not not6669(N20900,in0);
not not6670(N20901,in1);
not not6671(N20902,R0);
not not6672(N20903,R1);
not not6673(N20904,R2);
not not6674(N20917,in0);
not not6675(N20918,in1);
not not6676(N20919,R2);
not not6677(N20933,in0);
not not6678(N20934,in2);
not not6679(N20935,R2);
not not6680(N20949,in0);
not not6681(N20950,in2);
not not6682(N20951,R1);
not not6683(N20952,R2);
not not6684(N20965,in0);
not not6685(N20966,in1);
not not6686(N20967,R1);
not not6687(N20968,R2);
not not6688(N20981,in0);
not not6689(N20982,R1);
not not6690(N20983,R2);
not not6691(N20984,R3);
not not6692(N20997,in1);
not not6693(N20998,in2);
not not6694(N20999,R0);
not not6695(N21013,in0);
not not6696(N21014,in1);
not not6697(N21015,R0);
not not6698(N21016,R1);
not not6699(N21017,R3);
not not6700(N21029,in0);
not not6701(N21030,in2);
not not6702(N21031,R0);
not not6703(N21032,R1);
not not6704(N21045,in0);
not not6705(N21046,in1);
not not6706(N21047,R0);
not not6707(N21048,R2);
not not6708(N21049,R3);
not not6709(N21061,in0);
not not6710(N21062,in1);
not not6711(N21063,in2);
not not6712(N21064,R1);
not not6713(N21065,R2);
not not6714(N21077,in0);
not not6715(N21078,in1);
not not6716(N21079,R0);
not not6717(N21080,R1);
not not6718(N21081,R2);
not not6719(N21093,in0);
not not6720(N21094,in1);
not not6721(N21095,in2);
not not6722(N21096,R1);
not not6723(N21097,R2);
not not6724(N21109,in0);
not not6725(N21110,in1);
not not6726(N21111,R1);
not not6727(N21112,R2);
not not6728(N21113,R3);
not not6729(N21125,in0);
not not6730(N21126,in1);
not not6731(N21127,in2);
not not6732(N21128,R1);
not not6733(N21141,in0);
not not6734(N21142,in1);
not not6735(N21143,in2);
not not6736(N21144,R1);
not not6737(N21145,R3);
not not6738(N21157,in0);
not not6739(N21158,in1);
not not6740(N21159,in2);
not not6741(N21160,R1);
not not6742(N21161,R2);
not not6743(N21173,in0);
not not6744(N21174,in1);
not not6745(N21175,R0);
not not6746(N21176,R3);
not not6747(N21189,in0);
not not6748(N21190,in1);
not not6749(N21191,in2);
not not6750(N21192,R1);
not not6751(N21193,R2);
not not6752(N21205,in0);
not not6753(N21206,in1);
not not6754(N21207,in2);
not not6755(N21208,R3);
not not6756(N21221,in0);
not not6757(N21222,in1);
not not6758(N21223,in2);
not not6759(N21224,R2);
not not6760(N21237,in0);
not not6761(N21238,in1);
not not6762(N21239,in2);
not not6763(N21240,R0);
not not6764(N21253,in0);
not not6765(N21254,in1);
not not6766(N21255,R1);
not not6767(N21256,R2);
not not6768(N21269,in0);
not not6769(N21270,in2);
not not6770(N21271,R1);
not not6771(N21272,R2);
not not6772(N21273,R3);
not not6773(N21285,in0);
not not6774(N21286,in2);
not not6775(N21287,R0);
not not6776(N21288,R1);
not not6777(N21289,R2);
not not6778(N21301,in0);
not not6779(N21302,in2);
not not6780(N21303,R0);
not not6781(N21304,R2);
not not6782(N21317,in0);
not not6783(N21318,in2);
not not6784(N21319,R0);
not not6785(N21320,R1);
not not6786(N21332,in0);
not not6787(N21333,R0);
not not6788(N21347,in0);
not not6789(N21348,in1);
not not6790(N21349,in2);
not not6791(N21350,R1);
not not6792(N21362,in0);
not not6793(N21363,in1);
not not6794(N21364,R0);
not not6795(N21365,R1);
not not6796(N21366,R2);
not not6797(N21377,in0);
not not6798(N21378,in1);
not not6799(N21379,in2);
not not6800(N21380,R1);
not not6801(N21392,in0);
not not6802(N21393,in2);
not not6803(N21394,R3);
not not6804(N21407,in0);
not not6805(N21408,in1);
not not6806(N21409,R0);
not not6807(N21422,in0);
not not6808(N21423,in1);
not not6809(N21424,in2);
not not6810(N21425,R0);
not not6811(N21437,in0);
not not6812(N21438,in2);
not not6813(N21439,R1);
not not6814(N21440,R3);
not not6815(N21452,in0);
not not6816(N21453,in1);
not not6817(N21454,in2);
not not6818(N21455,R2);
not not6819(N21467,in0);
not not6820(N21468,in1);
not not6821(N21469,R3);
not not6822(N21482,in0);
not not6823(N21483,in1);
not not6824(N21484,R0);
not not6825(N21485,R1);
not not6826(N21497,in0);
not not6827(N21498,in2);
not not6828(N21499,R0);
not not6829(N21512,in1);
not not6830(N21513,R1);
not not6831(N21514,R3);
not not6832(N21527,in2);
not not6833(N21528,R1);
not not6834(N21529,R3);
not not6835(N21542,in0);
not not6836(N21543,in1);
not not6837(N21544,in2);
not not6838(N21545,R1);
not not6839(N21546,R2);
not not6840(N21557,in0);
not not6841(N21558,in2);
not not6842(N21559,R0);
not not6843(N21572,in0);
not not6844(N21573,in1);
not not6845(N21574,in2);
not not6846(N21575,R2);
not not6847(N21587,in0);
not not6848(N21588,R0);
not not6849(N21589,R1);
not not6850(N21602,in0);
not not6851(N21603,in2);
not not6852(N21617,in0);
not not6853(N21618,R0);
not not6854(N21619,R1);
not not6855(N21620,R2);
not not6856(N21632,in1);
not not6857(N21633,in2);
not not6858(N21634,R0);
not not6859(N21635,R1);
not not6860(N21647,in0);
not not6861(N21648,in1);
not not6862(N21649,R1);
not not6863(N21650,R2);
not not6864(N21651,R3);
not not6865(N21662,in0);
not not6866(N21663,R1);
not not6867(N21664,R2);
not not6868(N21665,R3);
not not6869(N21677,in0);
not not6870(N21678,in2);
not not6871(N21679,R0);
not not6872(N21680,R1);
not not6873(N21692,in0);
not not6874(N21693,R1);
not not6875(N21706,in0);
not not6876(N21707,in1);
not not6877(N21708,R1);
not not6878(N21709,R3);
not not6879(N21720,in0);
not not6880(N21721,R0);
not not6881(N21722,R1);
not not6882(N21723,R3);
not not6883(N21734,in0);
not not6884(N21735,R0);
not not6885(N21736,R3);
not not6886(N21748,R0);
not not6887(N21762,in2);
not not6888(N21763,R0);
not not6889(N21776,in0);
not not6890(N21777,in2);
not not6891(N21778,R0);
not not6892(N21790,in0);
not not6893(N21791,R1);
not not6894(N21792,R2);
not not6895(N21804,in0);
not not6896(N21805,in2);
not not6897(N21806,R2);
not not6898(N21818,in0);
not not6899(N21819,in1);
not not6900(N21820,R0);
not not6901(N21832,in0);
not not6902(N21833,R0);
not not6903(N21834,R3);
not not6904(N21846,in0);
not not6905(N21847,in2);
not not6906(N21848,R0);
not not6907(N21860,in0);
not not6908(N21861,in1);
not not6909(N21862,in2);
not not6910(N21874,in0);
not not6911(N21875,R1);
not not6912(N21888,in0);
not not6913(N21889,R2);
not not6914(N21890,R3);
not not6915(N21902,in0);
not not6916(N21903,in1);
not not6917(N21904,R2);
not not6918(N21916,in0);
not not6919(N21917,in1);
not not6920(N21918,in2);
not not6921(N21919,R0);
not not6922(N21930,in0);
not not6923(N21931,R1);
not not6924(N21932,R3);
not not6925(N21944,in0);
not not6926(N21945,in1);
not not6927(N21946,in2);
not not6928(N21958,in0);
not not6929(N21959,in2);
not not6930(N21960,R3);
not not6931(N21972,in0);
not not6932(N21973,R1);
not not6933(N21974,R2);
not not6934(N21986,in0);
not not6935(N21987,in1);
not not6936(N21988,R1);
not not6937(N22000,in0);
not not6938(N22001,R3);
not not6939(N22014,in0);
not not6940(N22015,R1);
not not6941(N22016,R2);
not not6942(N22028,in0);
not not6943(N22029,in1);
not not6944(N22042,in0);
not not6945(N22043,in1);
not not6946(N22044,R2);
not not6947(N22056,in0);
not not6948(N22057,R2);
not not6949(N22070,in0);
not not6950(N22071,in2);
not not6951(N22072,R1);
not not6952(N22084,in0);
not not6953(N22085,R1);
not not6954(N22086,R3);
not not6955(N22098,in0);
not not6956(N22099,R2);
not not6957(N22112,in0);
not not6958(N22113,in1);
not not6959(N22114,R0);
not not6960(N22126,in0);
not not6961(N22127,in1);
not not6962(N22128,R0);
not not6963(N22140,in0);
not not6964(N22141,in1);
not not6965(N22142,R0);
not not6966(N22143,R1);
not not6967(N22154,in0);
not not6968(N22155,in1);
not not6969(N22156,R1);
not not6970(N22157,R2);
not not6971(N22168,in0);
not not6972(N22169,R1);
not not6973(N22170,R2);
not not6974(N22182,in0);
not not6975(N22183,in1);
not not6976(N22184,R2);
not not6977(N22196,in0);
not not6978(N22197,in1);
not not6979(N22198,R0);
not not6980(N22199,R1);
not not6981(N22210,in0);
not not6982(N22211,in2);
not not6983(N22212,R0);
not not6984(N22223,in0);
not not6985(N22224,in1);
not not6986(N22225,in2);
not not6987(N22226,R2);
not not6988(N22236,in0);
not not6989(N22237,in2);
not not6990(N22238,R1);
not not6991(N22249,in0);
not not6992(N22250,R3);
not not6993(N22262,in0);
not not6994(N22263,R0);
not not6995(N22275,in2);
not not6996(N22276,R2);
not not6997(N22288,in0);
not not6998(N22289,R1);
not not6999(N22301,in0);
not not7000(N22314,in0);
not not7001(N22315,in2);
not not7002(N22316,R3);
not not7003(N22327,in0);
not not7004(N22328,in2);
not not7005(N22329,R1);
not not7006(N22330,R2);
not not7007(N22340,in0);
not not7008(N22341,in2);
not not7009(N22342,R2);
not not7010(N22353,in0);
not not7011(N22354,in1);
not not7012(N22355,R3);
not not7013(N22366,in0);
not not7014(N22367,in2);
not not7015(N22368,R0);
not not7016(N22379,in2);
not not7017(N22392,in0);
not not7018(N22393,in2);
not not7019(N22394,R1);
not not7020(N22395,R3);
not not7021(N22405,in0);
not not7022(N22406,R0);
not not7023(N22407,R2);
not not7024(N22418,R1);
not not7025(N22431,in0);
not not7026(N22432,in1);
not not7027(N22444,in0);
not not7028(N22445,in2);
not not7029(N22446,R2);
not not7030(N22457,in0);
not not7031(N22458,in1);
not not7032(N22459,R3);
not not7033(N22470,in0);
not not7034(N22471,in1);
not not7035(N22472,R3);
not not7036(N22483,in0);
not not7037(N22484,R0);
not not7038(N22485,R3);
not not7039(N22496,in0);
not not7040(N22497,in2);
not not7041(N22498,R0);
not not7042(N22509,in0);
not not7043(N22510,in2);
not not7044(N22511,R0);
not not7045(N22512,R1);
not not7046(N22522,in0);
not not7047(N22523,in1);
not not7048(N22535,R1);
not not7049(N22536,R2);
not not7050(N22548,in0);
not not7051(N22549,R1);
not not7052(N22561,R0);
not not7053(N22562,R1);
not not7054(N22574,in2);
not not7055(N22575,R0);
not not7056(N22576,R1);
not not7057(N22587,in0);
not not7058(N22588,R2);
not not7059(N22600,in1);
not not7060(N22601,in2);
not not7061(N22613,in0);
not not7062(N22614,R0);
not not7063(N22626,in0);
not not7064(N22627,in1);
not not7065(N22639,in0);
not not7066(N22640,R1);
not not7067(N22641,R2);
not not7068(N22652,in0);
not not7069(N22653,in2);
not not7070(N22654,R2);
not not7071(N22665,in0);
not not7072(N22666,R1);
not not7073(N22667,R2);
not not7074(N22678,R1);
not not7075(N22679,R2);
not not7076(N22691,in0);
not not7077(N22703,in0);
not not7078(N22704,in1);
not not7079(N22715,in0);
not not7080(N22716,in1);
not not7081(N22717,R0);
not not7082(N22727,in0);
not not7083(N22728,in1);
not not7084(N22729,R3);
not not7085(N22739,in0);
not not7086(N22740,R0);
not not7087(N22741,R1);
not not7088(N22751,in1);
not not7089(N22752,R0);
not not7090(N22763,in0);
not not7091(N22764,R1);
not not7092(N22775,in2);
not not7093(N22776,R0);
not not7094(N22787,in0);
not not7095(N22788,R0);
not not7096(N22799,in0);
not not7097(N22800,R0);
not not7098(N22801,R1);
not not7099(N22811,in0);
not not7100(N22812,in1);
not not7101(N22813,R2);
not not7102(N22823,in0);
not not7103(N22824,R0);
not not7104(N22825,R3);
not not7105(N22835,in0);
not not7106(N22836,in1);
not not7107(N22847,in0);
not not7108(N22848,R0);
not not7109(N22849,R1);
not not7110(N22859,in0);
not not7111(N22860,R1);
not not7112(N22871,R1);
not not7113(N22872,R3);
not not7114(N22883,in0);
not not7115(N22895,in1);
not not7116(N22907,R2);
not not7117(N22931,in0);
not not7118(N22942,in0);
not not7119(N22943,R0);
not not7120(N22953,in0);
not not7121(N22964,in0);
not not7122(N22997,in0);
not not7123(N22998,in2);
not not7124(N23008,R0);
not not7125(N23019,in0);
not not7126(N23038,in0);
not not7127(N23039,R0);
not not7128(N23040,R1);
not not7129(N23041,R2);
not not7130(N23042,R3);
not not7131(N23043,R5);
not not7132(N23054,in0);
not not7133(N23055,in2);
not not7134(N23056,R0);
not not7135(N23057,R2);
not not7136(N23058,R3);
not not7137(N23059,R4);
not not7138(N23070,in0);
not not7139(N23071,in2);
not not7140(N23072,R0);
not not7141(N23073,R2);
not not7142(N23074,R3);
not not7143(N23075,R4);
not not7144(N23076,R5);
not not7145(N23086,in0);
not not7146(N23087,in2);
not not7147(N23088,R0);
not not7148(N23089,R2);
not not7149(N23090,R5);
not not7150(N23101,R0);
not not7151(N23102,R1);
not not7152(N23103,R3);
not not7153(N23104,R4);
not not7154(N23105,R5);
not not7155(N23116,in0);
not not7156(N23117,in1);
not not7157(N23118,in2);
not not7158(N23119,R0);
not not7159(N23120,R3);
not not7160(N23131,in0);
not not7161(N23132,R0);
not not7162(N23133,R2);
not not7163(N23134,R4);
not not7164(N23145,in0);
not not7165(N23146,in1);
not not7166(N23147,R1);
not not7167(N23148,R3);
not not7168(N23159,in0);
not not7169(N23160,in2);
not not7170(N23161,R1);
not not7171(N23162,R4);
not not7172(N23163,R5);
not not7173(N23173,in0);
not not7174(N23174,R1);
not not7175(N23175,R2);
not not7176(N23176,R4);
not not7177(N23187,in0);
not not7178(N23188,in1);
not not7179(N23189,in2);
not not7180(N23190,R1);
not not7181(N23201,in0);
not not7182(N23202,in1);
not not7183(N23203,R1);
not not7184(N23204,R4);
not not7185(N23205,R5);
not not7186(N23215,in0);
not not7187(N23216,in2);
not not7188(N23217,R0);
not not7189(N23218,R1);
not not7190(N23219,R2);
not not7191(N23229,in0);
not not7192(N23230,R0);
not not7193(N23231,R1);
not not7194(N23232,R4);
not not7195(N23233,R5);
not not7196(N23243,in0);
not not7197(N23244,in2);
not not7198(N23245,R0);
not not7199(N23256,R1);
not not7200(N23257,R2);
not not7201(N23258,R3);
not not7202(N23259,R4);
not not7203(N23269,R3);
not not7204(N23270,R4);
not not7205(N23271,R5);
not not7206(N23282,R0);
not not7207(N23283,R1);
not not7208(N23284,R4);
not not7209(N23285,R5);
not not7210(N23295,R0);
not not7211(N23296,R1);
not not7212(N23297,R3);
not not7213(N23308,in0);
not not7214(N23309,in2);
not not7215(N23310,R0);
not not7216(N23311,R4);
not not7217(N23312,R5);
not not7218(N23321,in0);
not not7219(N23322,in1);
not not7220(N23323,in2);
not not7221(N23324,R1);
not not7222(N23325,R4);
not not7223(N23334,in0);
not not7224(N23335,in1);
not not7225(N23336,R1);
not not7226(N23337,R5);
not not7227(N23347,in0);
not not7228(N23348,in1);
not not7229(N23349,in2);
not not7230(N23350,R3);
not not7231(N23360,in0);
not not7232(N23361,in1);
not not7233(N23362,R0);
not not7234(N23363,R1);
not not7235(N23364,R3);
not not7236(N23373,in0);
not not7237(N23374,in1);
not not7238(N23375,R0);
not not7239(N23376,R1);
not not7240(N23377,R2);
not not7241(N23386,in0);
not not7242(N23387,R0);
not not7243(N23388,R1);
not not7244(N23389,R3);
not not7245(N23399,in1);
not not7246(N23400,R1);
not not7247(N23401,R2);
not not7248(N23402,R4);
not not7249(N23412,in2);
not not7250(N23413,R1);
not not7251(N23414,R2);
not not7252(N23415,R4);
not not7253(N23425,in0);
not not7254(N23426,R1);
not not7255(N23427,R3);
not not7256(N23428,R4);
not not7257(N23438,in2);
not not7258(N23439,R1);
not not7259(N23440,R2);
not not7260(N23441,R4);
not not7261(N23451,R2);
not not7262(N23452,R4);
not not7263(N23453,R5);
not not7264(N23463,R2);
not not7265(N23464,R5);
not not7266(N23475,in1);
not not7267(N23476,R0);
not not7268(N23487,in0);
not not7269(N23488,R3);
not not7270(N23489,R5);
not not7271(N23499,in0);
not not7272(N23500,in2);
not not7273(N23501,R1);
not not7274(N23511,in1);
not not7275(N23512,R2);
not not7276(N23513,R5);
not not7277(N23523,in0);
not not7278(N23524,in2);
not not7279(N23525,R3);
not not7280(N23535,R0);
not not7281(N23536,R1);
not not7282(N23537,R2);
not not7283(N23547,R2);
not not7284(N23548,R4);
not not7285(N23549,R5);
not not7286(N23559,in1);
not not7287(N23560,R1);
not not7288(N23561,R3);
not not7289(N23571,in1);
not not7290(N23572,R0);
not not7291(N23573,R1);
not not7292(N23574,R4);
not not7293(N23583,in1);
not not7294(N23584,R5);
not not7295(N23595,in2);
not not7296(N23596,R1);
not not7297(N23597,R3);
not not7298(N23607,in2);
not not7299(N23608,R0);
not not7300(N23609,R1);
not not7301(N23610,R4);
not not7302(N23619,R0);
not not7303(N23620,R2);
not not7304(N23621,R4);
not not7305(N23630,R3);
not not7306(N23631,R5);
not not7307(N23641,in0);
not not7308(N23642,R5);
not not7309(N23652,R3);
not not7310(N23653,R5);
not not7311(N23663,R3);
not not7312(N23664,R5);
not not7313(N23674,R1);
not not7314(N23675,R3);
not not7315(N23685,R1);
not not7316(N23686,R3);
not not7317(N23696,R0);
not not7318(N23697,R1);
not not7319(N23698,R4);
not not7320(N23707,R0);
not not7321(N23718,in0);
not not7322(N23719,R1);
not not7323(N23729,R4);
not not7324(N23747,R0);
not not7325(N23748,R1);
not not7326(N23749,R2);
not not7327(N23750,R4);
not not7328(N23751,R5);
not not7329(N23752,R6);
not not7330(N23760,R0);
not not7331(N23761,R1);
not not7332(N23762,R3);
not not7333(N23763,R4);
not not7334(N23764,R6);
not not7335(N23772,R0);
not not7336(N23773,R2);
not not7337(N23774,R6);
not not7338(N23775,R7);
not not7339(N23783,R1);
not not7340(N23784,R3);
not not7341(N23785,R4);
not not7342(N23786,R7);
not not7343(N23794,R0);
not not7344(N23795,R1);
not not7345(N23796,R5);
not not7346(N23804,R2);
not not7347(N23805,R4);
not not7348(N23806,R6);
not not7349(N23814,R1);
not not7350(N23822,R1);
not not7351(N20647,R3);
not not7352(N20648,R4);
not not7353(N20649,R5);
not not7354(N20650,R7);
not not7355(N20665,R3);
not not7356(N20666,R5);
not not7357(N20667,R6);
not not7358(N20668,R7);
not not7359(N20684,R4);
not not7360(N20685,R6);
not not7361(N20686,R7);
not not7362(N20701,R4);
not not7363(N20702,R5);
not not7364(N20703,R7);
not not7365(N20718,R5);
not not7366(N20719,R6);
not not7367(N20720,R7);
not not7368(N20734,R4);
not not7369(N20735,R5);
not not7370(N20736,R6);
not not7371(N20737,R7);
not not7372(N20752,R4);
not not7373(N20753,R6);
not not7374(N20754,R7);
not not7375(N20769,R3);
not not7376(N20770,R4);
not not7377(N20771,R6);
not not7378(N20786,R4);
not not7379(N20787,R5);
not not7380(N20788,R6);
not not7381(N20803,R4);
not not7382(N20804,R5);
not not7383(N20805,R7);
not not7384(N20821,R6);
not not7385(N20822,R7);
not not7386(N20838,R6);
not not7387(N20839,R7);
not not7388(N20855,R4);
not not7389(N20856,R7);
not not7390(N20872,R5);
not not7391(N20873,R6);
not not7392(N20889,R3);
not not7393(N20890,R6);
not not7394(N20905,R4);
not not7395(N20906,R5);
not not7396(N20907,R7);
not not7397(N20920,R3);
not not7398(N20921,R4);
not not7399(N20922,R5);
not not7400(N20923,R6);
not not7401(N20936,R3);
not not7402(N20937,R5);
not not7403(N20938,R6);
not not7404(N20939,R7);
not not7405(N20953,R5);
not not7406(N20954,R6);
not not7407(N20955,R7);
not not7408(N20969,R3);
not not7409(N20970,R5);
not not7410(N20971,R6);
not not7411(N20985,R4);
not not7412(N20986,R6);
not not7413(N20987,R7);
not not7414(N21000,R4);
not not7415(N21001,R5);
not not7416(N21002,R6);
not not7417(N21003,R7);
not not7418(N21018,R4);
not not7419(N21019,R7);
not not7420(N21033,R4);
not not7421(N21034,R5);
not not7422(N21035,R7);
not not7423(N21050,R4);
not not7424(N21051,R6);
not not7425(N21066,R5);
not not7426(N21067,R6);
not not7427(N21082,R4);
not not7428(N21083,R6);
not not7429(N21098,R3);
not not7430(N21099,R4);
not not7431(N21114,R6);
not not7432(N21115,R7);
not not7433(N21129,R5);
not not7434(N21130,R6);
not not7435(N21131,R7);
not not7436(N21146,R4);
not not7437(N21147,R5);
not not7438(N21162,R5);
not not7439(N21163,R7);
not not7440(N21177,R4);
not not7441(N21178,R6);
not not7442(N21179,R7);
not not7443(N21194,R3);
not not7444(N21195,R7);
not not7445(N21209,R4);
not not7446(N21210,R6);
not not7447(N21211,R7);
not not7448(N21225,R4);
not not7449(N21226,R5);
not not7450(N21227,R7);
not not7451(N21241,R4);
not not7452(N21242,R5);
not not7453(N21243,R6);
not not7454(N21257,R4);
not not7455(N21258,R6);
not not7456(N21259,R7);
not not7457(N21274,R4);
not not7458(N21275,R5);
not not7459(N21290,R5);
not not7460(N21291,R7);
not not7461(N21305,R4);
not not7462(N21306,R5);
not not7463(N21307,R6);
not not7464(N21321,R4);
not not7465(N21322,R6);
not not7466(N21334,R3);
not not7467(N21335,R4);
not not7468(N21336,R5);
not not7469(N21337,R6);
not not7470(N21351,R4);
not not7471(N21352,R6);
not not7472(N21367,R4);
not not7473(N21381,R3);
not not7474(N21382,R5);
not not7475(N21395,R4);
not not7476(N21396,R5);
not not7477(N21397,R6);
not not7478(N21410,R5);
not not7479(N21411,R6);
not not7480(N21412,R7);
not not7481(N21426,R4);
not not7482(N21427,R7);
not not7483(N21441,R4);
not not7484(N21442,R7);
not not7485(N21456,R3);
not not7486(N21457,R6);
not not7487(N21470,R5);
not not7488(N21471,R6);
not not7489(N21472,R7);
not not7490(N21486,R5);
not not7491(N21487,R6);
not not7492(N21500,R4);
not not7493(N21501,R6);
not not7494(N21502,R7);
not not7495(N21515,R5);
not not7496(N21516,R6);
not not7497(N21517,R7);
not not7498(N21530,R5);
not not7499(N21531,R6);
not not7500(N21532,R7);
not not7501(N21547,R4);
not not7502(N21560,R4);
not not7503(N21561,R5);
not not7504(N21562,R7);
not not7505(N21576,R4);
not not7506(N21577,R6);
not not7507(N21590,R3);
not not7508(N21591,R6);
not not7509(N21592,R7);
not not7510(N21604,R4);
not not7511(N21605,R5);
not not7512(N21606,R6);
not not7513(N21607,R7);
not not7514(N21621,R6);
not not7515(N21622,R7);
not not7516(N21636,R4);
not not7517(N21637,R7);
not not7518(N21652,R4);
not not7519(N21666,R5);
not not7520(N21667,R7);
not not7521(N21681,R3);
not not7522(N21682,R4);
not not7523(N21694,R4);
not not7524(N21695,R6);
not not7525(N21696,R7);
not not7526(N21710,R6);
not not7527(N21724,R6);
not not7528(N21737,R4);
not not7529(N21738,R5);
not not7530(N21749,R4);
not not7531(N21750,R5);
not not7532(N21751,R6);
not not7533(N21752,R7);
not not7534(N21764,R5);
not not7535(N21765,R6);
not not7536(N21766,R7);
not not7537(N21779,R5);
not not7538(N21780,R7);
not not7539(N21793,R6);
not not7540(N21794,R7);
not not7541(N21807,R6);
not not7542(N21808,R7);
not not7543(N21821,R4);
not not7544(N21822,R6);
not not7545(N21835,R4);
not not7546(N21836,R7);
not not7547(N21849,R4);
not not7548(N21850,R6);
not not7549(N21863,R5);
not not7550(N21864,R7);
not not7551(N21876,R4);
not not7552(N21877,R6);
not not7553(N21878,R7);
not not7554(N21891,R4);
not not7555(N21892,R6);
not not7556(N21905,R5);
not not7557(N21906,R6);
not not7558(N21920,R5);
not not7559(N21933,R4);
not not7560(N21934,R5);
not not7561(N21947,R5);
not not7562(N21948,R6);
not not7563(N21961,R4);
not not7564(N21962,R5);
not not7565(N21975,R4);
not not7566(N21976,R7);
not not7567(N21989,R4);
not not7568(N21990,R7);
not not7569(N22002,R4);
not not7570(N22003,R6);
not not7571(N22004,R7);
not not7572(N22017,R6);
not not7573(N22018,R7);
not not7574(N22030,R4);
not not7575(N22031,R5);
not not7576(N22032,R6);
not not7577(N22045,R6);
not not7578(N22046,R7);
not not7579(N22058,R4);
not not7580(N22059,R5);
not not7581(N22060,R7);
not not7582(N22073,R5);
not not7583(N22074,R6);
not not7584(N22087,R6);
not not7585(N22088,R7);
not not7586(N22100,R3);
not not7587(N22101,R6);
not not7588(N22102,R7);
not not7589(N22115,R5);
not not7590(N22116,R7);
not not7591(N22129,R4);
not not7592(N22130,R5);
not not7593(N22144,R3);
not not7594(N22158,R6);
not not7595(N22171,R4);
not not7596(N22172,R5);
not not7597(N22185,R5);
not not7598(N22186,R6);
not not7599(N22200,R7);
not not7600(N22213,R7);
not not7601(N22239,R6);
not not7602(N22251,R4);
not not7603(N22252,R7);
not not7604(N22264,R6);
not not7605(N22265,R7);
not not7606(N22277,R5);
not not7607(N22278,R6);
not not7608(N22290,R4);
not not7609(N22291,R5);
not not7610(N22302,R4);
not not7611(N22303,R6);
not not7612(N22304,R7);
not not7613(N22317,R6);
not not7614(N22343,R4);
not not7615(N22356,R5);
not not7616(N22369,R4);
not not7617(N22380,R5);
not not7618(N22381,R6);
not not7619(N22382,R7);
not not7620(N22408,R6);
not not7621(N22419,R3);
not not7622(N22420,R5);
not not7623(N22421,R6);
not not7624(N22433,R4);
not not7625(N22434,R5);
not not7626(N22447,R5);
not not7627(N22460,R6);
not not7628(N22473,R4);
not not7629(N22486,R6);
not not7630(N22499,R3);
not not7631(N22524,R5);
not not7632(N22525,R6);
not not7633(N22537,R4);
not not7634(N22538,R6);
not not7635(N22550,R4);
not not7636(N22551,R6);
not not7637(N22563,R4);
not not7638(N22564,R5);
not not7639(N22577,R4);
not not7640(N22589,R4);
not not7641(N22590,R7);
not not7642(N22602,R4);
not not7643(N22603,R5);
not not7644(N22615,R4);
not not7645(N22616,R7);
not not7646(N22628,R4);
not not7647(N22629,R6);
not not7648(N22642,R5);
not not7649(N22655,R7);
not not7650(N22668,R6);
not not7651(N22680,R4);
not not7652(N22681,R7);
not not7653(N22692,R6);
not not7654(N22693,R7);
not not7655(N22705,R7);
not not7656(N22753,R5);
not not7657(N22765,R4);
not not7658(N22777,R5);
not not7659(N22789,R6);
not not7660(N22837,R7);
not not7661(N22861,R7);
not not7662(N22873,R6);
not not7663(N22884,R3);
not not7664(N22885,R4);
not not7665(N22896,R4);
not not7666(N22897,R7);
not not7667(N22908,R5);
not not7668(N22909,R6);
not not7669(N22919,R5);
not not7670(N22920,R6);
not not7671(N22921,R7);
not not7672(N22932,R3);
not not7673(N22954,R5);
not not7674(N22965,R5);
not not7675(N22975,R4);
not not7676(N22976,R5);
not not7677(N22986,R4);
not not7678(N22987,R5);
not not7679(N23009,R5);
not not7680(N23029,R6);
not not7681(N23044,R6);
not not7682(N23045,R7);
not not7683(N23060,R5);
not not7684(N23061,R6);
not not7685(N23077,R6);
not not7686(N23091,R6);
not not7687(N23092,R7);
not not7688(N23106,R6);
not not7689(N23107,R7);
not not7690(N23121,R5);
not not7691(N23122,R6);
not not7692(N23135,R6);
not not7693(N23136,R7);
not not7694(N23149,R4);
not not7695(N23150,R6);
not not7696(N23164,R7);
not not7697(N23177,R5);
not not7698(N23178,R6);
not not7699(N23191,R6);
not not7700(N23192,R7);
not not7701(N23206,R6);
not not7702(N23220,R4);
not not7703(N23234,R6);
not not7704(N23246,R6);
not not7705(N23247,R7);
not not7706(N23260,R6);
not not7707(N23272,R6);
not not7708(N23273,R7);
not not7709(N23286,R7);
not not7710(N23298,R6);
not not7711(N23299,R7);
not not7712(N23338,R7);
not not7713(N23351,R5);
not not7714(N23390,R5);
not not7715(N23403,R7);
not not7716(N23416,R6);
not not7717(N23429,R6);
not not7718(N23442,R7);
not not7719(N23454,R7);
not not7720(N23465,R6);
not not7721(N23466,R7);
not not7722(N23477,R5);
not not7723(N23478,R6);
not not7724(N23490,R6);
not not7725(N23502,R7);
not not7726(N23514,R6);
not not7727(N23526,R6);
not not7728(N23538,R6);
not not7729(N23550,R6);
not not7730(N23562,R6);
not not7731(N23585,R6);
not not7732(N23586,R7);
not not7733(N23598,R6);
not not7734(N23632,R7);
not not7735(N23643,R7);
not not7736(N23654,R6);
not not7737(N23665,R6);
not not7738(N23676,R7);
not not7739(N23687,R7);
not not7740(N23708,R5);
not not7741(N23709,R6);
not not7742(N23720,R7);
not not7743(N23730,R7);
not not7744(N23739,R6);
not not7745(N24200,in0);
not not7746(N24201,in1);
not not7747(N24202,R0);
not not7748(N24203,R2);
not not7749(N24204,R3);
not not7750(N24218,in0);
not not7751(N24219,in1);
not not7752(N24220,R1);
not not7753(N24221,R2);
not not7754(N24222,R3);
not not7755(N24236,in1);
not not7756(N24237,in2);
not not7757(N24238,R0);
not not7758(N24239,R1);
not not7759(N24240,R2);
not not7760(N24241,R3);
not not7761(N24254,in0);
not not7762(N24255,in1);
not not7763(N24256,R0);
not not7764(N24257,R1);
not not7765(N24258,R2);
not not7766(N24259,R3);
not not7767(N24272,in1);
not not7768(N24273,R0);
not not7769(N24274,R1);
not not7770(N24275,R2);
not not7771(N24276,R3);
not not7772(N24290,in0);
not not7773(N24291,in2);
not not7774(N24292,R1);
not not7775(N24293,R2);
not not7776(N24294,R3);
not not7777(N24308,in1);
not not7778(N24309,in2);
not not7779(N24310,R0);
not not7780(N24311,R1);
not not7781(N24312,R2);
not not7782(N24326,in1);
not not7783(N24327,in2);
not not7784(N24328,R0);
not not7785(N24329,R2);
not not7786(N24330,R3);
not not7787(N24343,in1);
not not7788(N24344,in2);
not not7789(N24345,R1);
not not7790(N24346,R2);
not not7791(N24347,R3);
not not7792(N24360,in0);
not not7793(N24361,R0);
not not7794(N24362,R2);
not not7795(N24363,R3);
not not7796(N24377,in1);
not not7797(N24378,R0);
not not7798(N24379,R1);
not not7799(N24380,R3);
not not7800(N24394,in0);
not not7801(N24395,in1);
not not7802(N24396,in2);
not not7803(N24397,R0);
not not7804(N24398,R3);
not not7805(N24411,in0);
not not7806(N24412,R0);
not not7807(N24413,R1);
not not7808(N24414,R2);
not not7809(N24415,R3);
not not7810(N24428,in0);
not not7811(N24429,in1);
not not7812(N24430,in2);
not not7813(N24431,R0);
not not7814(N24432,R1);
not not7815(N24433,R2);
not not7816(N24445,in0);
not not7817(N24446,in1);
not not7818(N24447,in2);
not not7819(N24448,R0);
not not7820(N24449,R1);
not not7821(N24450,R2);
not not7822(N24462,in0);
not not7823(N24463,in1);
not not7824(N24464,in2);
not not7825(N24465,R0);
not not7826(N24466,R1);
not not7827(N24467,R2);
not not7828(N24479,in0);
not not7829(N24480,R0);
not not7830(N24481,R2);
not not7831(N24495,in0);
not not7832(N24496,in1);
not not7833(N24497,R0);
not not7834(N24511,R0);
not not7835(N24512,R1);
not not7836(N24513,R2);
not not7837(N24514,R3);
not not7838(N24527,in2);
not not7839(N24528,R1);
not not7840(N24529,R2);
not not7841(N24530,R3);
not not7842(N24543,R0);
not not7843(N24544,R1);
not not7844(N24545,R3);
not not7845(N24559,in0);
not not7846(N24560,R1);
not not7847(N24561,R3);
not not7848(N24575,R0);
not not7849(N24576,R1);
not not7850(N24577,R2);
not not7851(N24578,R3);
not not7852(N24591,in2);
not not7853(N24592,R1);
not not7854(N24593,R2);
not not7855(N24594,R3);
not not7856(N24607,R0);
not not7857(N24608,R1);
not not7858(N24609,R2);
not not7859(N24623,in2);
not not7860(N24624,R1);
not not7861(N24625,R2);
not not7862(N24639,in0);
not not7863(N24640,in1);
not not7864(N24641,R0);
not not7865(N24642,R1);
not not7866(N24643,R3);
not not7867(N24655,in0);
not not7868(N24656,in2);
not not7869(N24657,R3);
not not7870(N24671,in0);
not not7871(N24672,in1);
not not7872(N24673,R0);
not not7873(N24674,R1);
not not7874(N24687,in0);
not not7875(N24688,in2);
not not7876(N24689,R2);
not not7877(N24690,R3);
not not7878(N24703,in0);
not not7879(N24704,in1);
not not7880(N24705,in2);
not not7881(N24706,R1);
not not7882(N24719,in0);
not not7883(N24720,R0);
not not7884(N24721,R1);
not not7885(N24735,in0);
not not7886(N24736,in1);
not not7887(N24737,in2);
not not7888(N24738,R1);
not not7889(N24739,R2);
not not7890(N24751,in0);
not not7891(N24752,in2);
not not7892(N24753,R0);
not not7893(N24754,R1);
not not7894(N24767,in0);
not not7895(N24768,in1);
not not7896(N24769,in2);
not not7897(N24770,R0);
not not7898(N24783,in0);
not not7899(N24784,in2);
not not7900(N24785,R1);
not not7901(N24786,R2);
not not7902(N24787,R3);
not not7903(N24799,in1);
not not7904(N24800,in2);
not not7905(N24801,R0);
not not7906(N24802,R1);
not not7907(N24803,R3);
not not7908(N24815,in0);
not not7909(N24816,R1);
not not7910(N24817,R2);
not not7911(N24818,R3);
not not7912(N24831,in0);
not not7913(N24832,in1);
not not7914(N24833,in2);
not not7915(N24834,R1);
not not7916(N24835,R2);
not not7917(N24847,in1);
not not7918(N24848,in2);
not not7919(N24849,R0);
not not7920(N24850,R1);
not not7921(N24863,in1);
not not7922(N24864,in2);
not not7923(N24865,R1);
not not7924(N24866,R2);
not not7925(N24879,in0);
not not7926(N24880,in1);
not not7927(N24881,in2);
not not7928(N24882,R0);
not not7929(N24883,R2);
not not7930(N24895,in0);
not not7931(N24896,in1);
not not7932(N24897,R0);
not not7933(N24898,R1);
not not7934(N24899,R2);
not not7935(N24911,in0);
not not7936(N24912,in2);
not not7937(N24913,R0);
not not7938(N24914,R1);
not not7939(N24915,R2);
not not7940(N24927,in0);
not not7941(N24928,in2);
not not7942(N24929,R0);
not not7943(N24930,R1);
not not7944(N24931,R2);
not not7945(N24943,in0);
not not7946(N24944,in2);
not not7947(N24945,R1);
not not7948(N24946,R2);
not not7949(N24947,R3);
not not7950(N24959,in0);
not not7951(N24960,R1);
not not7952(N24974,in0);
not not7953(N24975,in1);
not not7954(N24976,in2);
not not7955(N24977,R1);
not not7956(N24989,in1);
not not7957(N24990,R2);
not not7958(N24991,R3);
not not7959(N25004,in2);
not not7960(N25005,R2);
not not7961(N25006,R3);
not not7962(N25019,R1);
not not7963(N25020,R2);
not not7964(N25021,R3);
not not7965(N25034,in2);
not not7966(N25035,R1);
not not7967(N25036,R2);
not not7968(N25049,in0);
not not7969(N25050,in1);
not not7970(N25051,R1);
not not7971(N25052,R2);
not not7972(N25064,in0);
not not7973(N25065,R0);
not not7974(N25066,R1);
not not7975(N25079,in0);
not not7976(N25080,in1);
not not7977(N25081,R0);
not not7978(N25082,R1);
not not7979(N25083,R2);
not not7980(N25094,in0);
not not7981(N25095,in2);
not not7982(N25096,R0);
not not7983(N25097,R3);
not not7984(N25109,in0);
not not7985(N25110,in1);
not not7986(N25111,in2);
not not7987(N25112,R0);
not not7988(N25124,in0);
not not7989(N25125,in1);
not not7990(N25126,R0);
not not7991(N25139,in1);
not not7992(N25140,in2);
not not7993(N25141,R3);
not not7994(N25154,in0);
not not7995(N25155,in1);
not not7996(N25156,R0);
not not7997(N25157,R2);
not not7998(N25169,in0);
not not7999(N25170,in2);
not not8000(N25171,R0);
not not8001(N25172,R2);
not not8002(N25184,in0);
not not8003(N25185,in2);
not not8004(N25186,R0);
not not8005(N25187,R3);
not not8006(N25199,in0);
not not8007(N25200,in1);
not not8008(N25201,R0);
not not8009(N25202,R2);
not not8010(N25214,in0);
not not8011(N25215,in1);
not not8012(N25216,in2);
not not8013(N25217,R1);
not not8014(N25218,R3);
not not8015(N25229,in0);
not not8016(N25230,in2);
not not8017(N25231,R1);
not not8018(N25232,R2);
not not8019(N25233,R3);
not not8020(N25244,in0);
not not8021(N25245,in1);
not not8022(N25246,R1);
not not8023(N25247,R2);
not not8024(N25259,in0);
not not8025(N25260,R0);
not not8026(N25261,R1);
not not8027(N25262,R2);
not not8028(N25274,in1);
not not8029(N25275,in2);
not not8030(N25276,R1);
not not8031(N25289,in0);
not not8032(N25290,in1);
not not8033(N25291,in2);
not not8034(N25304,in0);
not not8035(N25305,in1);
not not8036(N25306,R1);
not not8037(N25307,R3);
not not8038(N25319,in2);
not not8039(N25320,R1);
not not8040(N25321,R2);
not not8041(N25322,R3);
not not8042(N25334,R0);
not not8043(N25335,R2);
not not8044(N25336,R3);
not not8045(N25349,in0);
not not8046(N25350,in2);
not not8047(N25351,R1);
not not8048(N25352,R2);
not not8049(N25364,in0);
not not8050(N25365,in1);
not not8051(N25366,in2);
not not8052(N25367,R0);
not not8053(N25368,R1);
not not8054(N25379,in1);
not not8055(N25380,in2);
not not8056(N25381,R2);
not not8057(N25394,in0);
not not8058(N25395,in1);
not not8059(N25396,R2);
not not8060(N25409,in0);
not not8061(N25410,in2);
not not8062(N25411,R0);
not not8063(N25412,R2);
not not8064(N25424,in0);
not not8065(N25425,R0);
not not8066(N25426,R1);
not not8067(N25438,in0);
not not8068(N25439,R0);
not not8069(N25440,R1);
not not8070(N25441,R3);
not not8071(N25452,in0);
not not8072(N25453,R3);
not not8073(N25466,in0);
not not8074(N25467,in1);
not not8075(N25468,R0);
not not8076(N25480,in0);
not not8077(N25481,in2);
not not8078(N25482,R0);
not not8079(N25494,in0);
not not8080(N25495,in2);
not not8081(N25508,in0);
not not8082(N25509,in1);
not not8083(N25510,in2);
not not8084(N25511,R1);
not not8085(N25522,R0);
not not8086(N25523,R1);
not not8087(N25524,R2);
not not8088(N25525,R3);
not not8089(N25536,in0);
not not8090(N25537,in2);
not not8091(N25538,R2);
not not8092(N25550,in0);
not not8093(N25551,in1);
not not8094(N25552,R1);
not not8095(N25564,in0);
not not8096(N25565,R0);
not not8097(N25578,in0);
not not8098(N25579,in1);
not not8099(N25580,in2);
not not8100(N25581,R2);
not not8101(N25592,in0);
not not8102(N25593,R0);
not not8103(N25594,R1);
not not8104(N25595,R2);
not not8105(N25606,R1);
not not8106(N25607,R2);
not not8107(N25620,in0);
not not8108(N25621,R1);
not not8109(N25634,in0);
not not8110(N25635,R1);
not not8111(N25648,in0);
not not8112(N25649,R1);
not not8113(N25650,R3);
not not8114(N25662,in0);
not not8115(N25663,in2);
not not8116(N25664,R2);
not not8117(N25676,in0);
not not8118(N25677,in1);
not not8119(N25678,in2);
not not8120(N25679,R0);
not not8121(N25680,R1);
not not8122(N25690,R0);
not not8123(N25691,R1);
not not8124(N25692,R3);
not not8125(N25704,in1);
not not8126(N25705,R0);
not not8127(N25706,R1);
not not8128(N25718,R1);
not not8129(N25719,R2);
not not8130(N25732,in0);
not not8131(N25733,in1);
not not8132(N25734,in2);
not not8133(N25735,R0);
not not8134(N25746,in1);
not not8135(N25747,in2);
not not8136(N25760,in0);
not not8137(N25761,in1);
not not8138(N25762,in2);
not not8139(N25774,R1);
not not8140(N25775,R3);
not not8141(N25788,in0);
not not8142(N25789,in1);
not not8143(N25790,in2);
not not8144(N25802,in0);
not not8145(N25803,R1);
not not8146(N25804,R3);
not not8147(N25816,in2);
not not8148(N25817,R1);
not not8149(N25818,R2);
not not8150(N25830,in0);
not not8151(N25831,R1);
not not8152(N25832,R2);
not not8153(N25844,in0);
not not8154(N25845,in2);
not not8155(N25858,in0);
not not8156(N25859,in1);
not not8157(N25860,R1);
not not8158(N25872,in0);
not not8159(N25873,in1);
not not8160(N25886,R1);
not not8161(N25887,R2);
not not8162(N25900,in2);
not not8163(N25901,R2);
not not8164(N25914,R1);
not not8165(N25915,R3);
not not8166(N25928,in2);
not not8167(N25929,R1);
not not8168(N25942,in0);
not not8169(N25943,R3);
not not8170(N25956,in1);
not not8171(N25957,in2);
not not8172(N25970,in0);
not not8173(N25971,in2);
not not8174(N25972,R2);
not not8175(N25984,in0);
not not8176(N25985,in1);
not not8177(N25986,R2);
not not8178(N25998,in0);
not not8179(N25999,in1);
not not8180(N26000,R0);
not not8181(N26012,in0);
not not8182(N26013,R2);
not not8183(N26026,in0);
not not8184(N26027,in2);
not not8185(N26028,R0);
not not8186(N26040,in0);
not not8187(N26041,R0);
not not8188(N26042,R1);
not not8189(N26043,R3);
not not8190(N26054,in0);
not not8191(N26055,in1);
not not8192(N26056,R3);
not not8193(N26068,in0);
not not8194(N26069,in2);
not not8195(N26070,R0);
not not8196(N26071,R1);
not not8197(N26082,in1);
not not8198(N26083,R1);
not not8199(N26084,R2);
not not8200(N26096,in0);
not not8201(N26097,in1);
not not8202(N26098,R1);
not not8203(N26099,R2);
not not8204(N26110,in1);
not not8205(N26124,in1);
not not8206(N26125,R0);
not not8207(N26126,R1);
not not8208(N26138,in1);
not not8209(N26139,R1);
not not8210(N26140,R3);
not not8211(N26152,in1);
not not8212(N26153,in2);
not not8213(N26154,R1);
not not8214(N26155,R3);
not not8215(N26166,in0);
not not8216(N26167,in1);
not not8217(N26168,R2);
not not8218(N26180,in0);
not not8219(N26181,R1);
not not8220(N26182,R3);
not not8221(N26193,in0);
not not8222(N26194,in1);
not not8223(N26195,R0);
not not8224(N26206,in0);
not not8225(N26207,R1);
not not8226(N26219,R1);
not not8227(N26220,R3);
not not8228(N26232,in2);
not not8229(N26245,R1);
not not8230(N26258,R0);
not not8231(N26259,R2);
not not8232(N26271,in0);
not not8233(N26272,in1);
not not8234(N26273,in2);
not not8235(N26284,in0);
not not8236(N26285,R1);
not not8237(N26286,R2);
not not8238(N26297,in0);
not not8239(N26298,in1);
not not8240(N26299,R1);
not not8241(N26300,R2);
not not8242(N26310,R1);
not not8243(N26323,in0);
not not8244(N26324,in2);
not not8245(N26325,R1);
not not8246(N26326,R3);
not not8247(N26336,in0);
not not8248(N26349,in0);
not not8249(N26350,in1);
not not8250(N26351,R0);
not not8251(N26352,R2);
not not8252(N26362,R1);
not not8253(N26363,R2);
not not8254(N26364,R3);
not not8255(N26375,in2);
not not8256(N26376,R1);
not not8257(N26377,R3);
not not8258(N26388,in0);
not not8259(N26389,R0);
not not8260(N26390,R2);
not not8261(N26401,in1);
not not8262(N26402,R0);
not not8263(N26414,in2);
not not8264(N26415,R0);
not not8265(N26427,in1);
not not8266(N26428,R1);
not not8267(N26429,R3);
not not8268(N26440,in0);
not not8269(N26441,in1);
not not8270(N26442,R0);
not not8271(N26453,in0);
not not8272(N26454,in2);
not not8273(N26466,R1);
not not8274(N26467,R2);
not not8275(N26479,in2);
not not8276(N26480,R1);
not not8277(N26481,R2);
not not8278(N26492,in0);
not not8279(N26493,in2);
not not8280(N26494,R2);
not not8281(N26505,in0);
not not8282(N26506,R0);
not not8283(N26518,in2);
not not8284(N26519,R0);
not not8285(N26520,R1);
not not8286(N26531,in2);
not not8287(N26532,R2);
not not8288(N26544,in0);
not not8289(N26545,R1);
not not8290(N26557,R2);
not not8291(N26570,in2);
not not8292(N26571,R0);
not not8293(N26572,R1);
not not8294(N26583,in0);
not not8295(N26584,R0);
not not8296(N26596,in0);
not not8297(N26597,R2);
not not8298(N26609,in0);
not not8299(N26610,in1);
not not8300(N26611,R2);
not not8301(N26622,in0);
not not8302(N26634,in0);
not not8303(N26646,in1);
not not8304(N26647,R0);
not not8305(N26658,R0);
not not8306(N26670,in0);
not not8307(N26671,R0);
not not8308(N26682,R0);
not not8309(N26694,in0);
not not8310(N26695,R3);
not not8311(N26706,in0);
not not8312(N26707,in2);
not not8313(N26718,R2);
not not8314(N26730,in0);
not not8315(N26731,R0);
not not8316(N26742,R1);
not not8317(N26754,in1);
not not8318(N26766,in0);
not not8319(N26767,in1);
not not8320(N26768,R0);
not not8321(N26778,R0);
not not8322(N26779,R3);
not not8323(N26790,in1);
not not8324(N26791,R3);
not not8325(N26802,R0);
not not8326(N26803,R2);
not not8327(N26814,in0);
not not8328(N26826,in0);
not not8329(N26827,R0);
not not8330(N26838,in2);
not not8331(N26850,in2);
not not8332(N26851,R3);
not not8333(N26862,in0);
not not8334(N26874,R1);
not not8335(N26886,R1);
not not8336(N26887,R2);
not not8337(N26888,R3);
not not8338(N26898,in1);
not not8339(N26910,in1);
not not8340(N26911,in2);
not not8341(N26934,in1);
not not8342(N26935,R3);
not not8343(N26946,in1);
not not8344(N26947,R3);
not not8345(N26958,in2);
not not8346(N26959,R3);
not not8347(N26970,in1);
not not8348(N26971,in2);
not not8349(N26982,in0);
not not8350(N26983,R1);
not not8351(N26984,R2);
not not8352(N26994,R0);
not not8353(N26995,R1);
not not8354(N27006,R1);
not not8355(N27007,R3);
not not8356(N27018,in2);
not not8357(N27019,R1);
not not8358(N27030,R1);
not not8359(N27042,in1);
not not8360(N27054,in2);
not not8361(N27066,in0);
not not8362(N27067,R0);
not not8363(N27077,in0);
not not8364(N27088,in0);
not not8365(N27089,in1);
not not8366(N27099,R3);
not not8367(N27110,R1);
not not8368(N27130,in0);
not not8369(N27140,R2);
not not8370(N27160,in1);
not not8371(N27170,in0);
not not8372(N27209,in2);
not not8373(N27210,R0);
not not8374(N27211,R2);
not not8375(N27212,R3);
not not8376(N27213,R4);
not not8377(N27214,R5);
not not8378(N27225,in1);
not not8379(N27226,R0);
not not8380(N27227,R1);
not not8381(N27228,R2);
not not8382(N27229,R3);
not not8383(N27230,R4);
not not8384(N27241,in0);
not not8385(N27242,in1);
not not8386(N27243,in2);
not not8387(N27244,R1);
not not8388(N27245,R4);
not not8389(N27256,in0);
not not8390(N27257,in1);
not not8391(N27258,in2);
not not8392(N27259,R3);
not not8393(N27260,R4);
not not8394(N27271,in0);
not not8395(N27272,in1);
not not8396(N27273,in2);
not not8397(N27274,R0);
not not8398(N27275,R1);
not not8399(N27276,R4);
not not8400(N27286,in2);
not not8401(N27287,R0);
not not8402(N27288,R1);
not not8403(N27289,R3);
not not8404(N27300,R1);
not not8405(N27301,R2);
not not8406(N27302,R3);
not not8407(N27303,R5);
not not8408(N27314,in1);
not not8409(N27315,R0);
not not8410(N27316,R1);
not not8411(N27317,R3);
not not8412(N27318,R4);
not not8413(N27328,in1);
not not8414(N27329,R1);
not not8415(N27330,R2);
not not8416(N27331,R3);
not not8417(N27332,R4);
not not8418(N27342,in1);
not not8419(N27343,R3);
not not8420(N27344,R4);
not not8421(N27345,R5);
not not8422(N27356,in2);
not not8423(N27357,R3);
not not8424(N27358,R4);
not not8425(N27359,R5);
not not8426(N27370,in0);
not not8427(N27371,in2);
not not8428(N27372,R0);
not not8429(N27373,R1);
not not8430(N27374,R3);
not not8431(N27384,in0);
not not8432(N27385,R1);
not not8433(N27386,R2);
not not8434(N27387,R4);
not not8435(N27398,in0);
not not8436(N27399,R0);
not not8437(N27400,R1);
not not8438(N27401,R3);
not not8439(N27402,R4);
not not8440(N27412,in1);
not not8441(N27413,R1);
not not8442(N27414,R2);
not not8443(N27415,R3);
not not8444(N27416,R5);
not not8445(N27426,in0);
not not8446(N27427,in2);
not not8447(N27428,R0);
not not8448(N27429,R1);
not not8449(N27440,in1);
not not8450(N27441,R0);
not not8451(N27442,R1);
not not8452(N27443,R2);
not not8453(N27444,R3);
not not8454(N27454,in1);
not not8455(N27455,R0);
not not8456(N27456,R2);
not not8457(N27457,R4);
not not8458(N27468,in0);
not not8459(N27469,in1);
not not8460(N27470,R1);
not not8461(N27471,R3);
not not8462(N27482,in1);
not not8463(N27483,R0);
not not8464(N27484,R1);
not not8465(N27485,R2);
not not8466(N27486,R4);
not not8467(N27496,in0);
not not8468(N27497,in1);
not not8469(N27498,R1);
not not8470(N27499,R3);
not not8471(N27500,R5);
not not8472(N27510,in1);
not not8473(N27511,R0);
not not8474(N27512,R3);
not not8475(N27513,R5);
not not8476(N27524,in0);
not not8477(N27525,in1);
not not8478(N27526,R1);
not not8479(N27527,R3);
not not8480(N27538,in2);
not not8481(N27539,R0);
not not8482(N27540,R3);
not not8483(N27541,R5);
not not8484(N27552,in0);
not not8485(N27553,in1);
not not8486(N27554,in2);
not not8487(N27555,R3);
not not8488(N27556,R4);
not not8489(N27566,in0);
not not8490(N27567,in1);
not not8491(N27568,in2);
not not8492(N27569,R4);
not not8493(N27570,R5);
not not8494(N27580,R0);
not not8495(N27581,R1);
not not8496(N27582,R2);
not not8497(N27583,R4);
not not8498(N27594,in0);
not not8499(N27595,in1);
not not8500(N27596,R0);
not not8501(N27597,R1);
not not8502(N27608,R2);
not not8503(N27609,R3);
not not8504(N27610,R4);
not not8505(N27611,R5);
not not8506(N27621,R0);
not not8507(N27622,R4);
not not8508(N27623,R5);
not not8509(N27634,in2);
not not8510(N27635,R1);
not not8511(N27636,R4);
not not8512(N27637,R5);
not not8513(N27647,in2);
not not8514(N27648,R0);
not not8515(N27649,R2);
not not8516(N27650,R4);
not not8517(N27660,in0);
not not8518(N27661,in2);
not not8519(N27662,R0);
not not8520(N27663,R1);
not not8521(N27673,in1);
not not8522(N27674,R2);
not not8523(N27675,R5);
not not8524(N27686,in1);
not not8525(N27687,R1);
not not8526(N27688,R3);
not not8527(N27689,R4);
not not8528(N27699,in0);
not not8529(N27700,in1);
not not8530(N27701,R4);
not not8531(N27712,in0);
not not8532(N27713,in2);
not not8533(N27714,R1);
not not8534(N27715,R3);
not not8535(N27716,R4);
not not8536(N27725,R0);
not not8537(N27726,R1);
not not8538(N27727,R3);
not not8539(N27738,in0);
not not8540(N27739,R1);
not not8541(N27740,R2);
not not8542(N27751,in1);
not not8543(N27752,R1);
not not8544(N27753,R2);
not not8545(N27754,R3);
not not8546(N27755,R4);
not not8547(N27764,R0);
not not8548(N27765,R1);
not not8549(N27766,R2);
not not8550(N27767,R5);
not not8551(N27777,in0);
not not8552(N27778,R0);
not not8553(N27779,R3);
not not8554(N27780,R4);
not not8555(N27790,in0);
not not8556(N27791,in2);
not not8557(N27792,R3);
not not8558(N27793,R4);
not not8559(N27803,in1);
not not8560(N27804,in2);
not not8561(N27805,R2);
not not8562(N27806,R4);
not not8563(N27816,R0);
not not8564(N27817,R1);
not not8565(N27818,R4);
not not8566(N27819,R5);
not not8567(N27829,in2);
not not8568(N27830,R1);
not not8569(N27831,R2);
not not8570(N27832,R4);
not not8571(N27842,in0);
not not8572(N27843,R0);
not not8573(N27844,R1);
not not8574(N27855,in1);
not not8575(N27856,R3);
not not8576(N27857,R4);
not not8577(N27858,R5);
not not8578(N27868,in0);
not not8579(N27869,in1);
not not8580(N27870,R1);
not not8581(N27871,R5);
not not8582(N27881,in0);
not not8583(N27882,in2);
not not8584(N27883,R1);
not not8585(N27884,R2);
not not8586(N27885,R4);
not not8587(N27894,in0);
not not8588(N27895,in1);
not not8589(N27896,R2);
not not8590(N27897,R5);
not not8591(N27907,in0);
not not8592(N27908,R4);
not not8593(N27909,R5);
not not8594(N27920,in1);
not not8595(N27921,in2);
not not8596(N27922,R1);
not not8597(N27923,R3);
not not8598(N27933,in0);
not not8599(N27934,R0);
not not8600(N27935,R1);
not not8601(N27936,R5);
not not8602(N27946,R0);
not not8603(N27947,R1);
not not8604(N27948,R3);
not not8605(N27949,R4);
not not8606(N27959,R1);
not not8607(N27960,R2);
not not8608(N27961,R3);
not not8609(N27962,R4);
not not8610(N27972,R2);
not not8611(N27973,R3);
not not8612(N27974,R5);
not not8613(N27985,in2);
not not8614(N27986,R1);
not not8615(N27987,R3);
not not8616(N27988,R4);
not not8617(N27998,R0);
not not8618(N27999,R1);
not not8619(N28000,R3);
not not8620(N28011,in2);
not not8621(N28012,R1);
not not8622(N28013,R3);
not not8623(N28024,in2);
not not8624(N28025,R0);
not not8625(N28026,R4);
not not8626(N28037,in0);
not not8627(N28038,in1);
not not8628(N28039,R1);
not not8629(N28040,R3);
not not8630(N28050,in0);
not not8631(N28051,in1);
not not8632(N28052,R1);
not not8633(N28053,R5);
not not8634(N28063,R0);
not not8635(N28064,R1);
not not8636(N28065,R2);
not not8637(N28066,R4);
not not8638(N28076,R0);
not not8639(N28077,R3);
not not8640(N28078,R5);
not not8641(N28089,in2);
not not8642(N28090,R4);
not not8643(N28091,R5);
not not8644(N28102,in0);
not not8645(N28103,in1);
not not8646(N28104,R1);
not not8647(N28114,in0);
not not8648(N28115,R3);
not not8649(N28126,R1);
not not8650(N28127,R2);
not not8651(N28138,in0);
not not8652(N28139,R2);
not not8653(N28140,R5);
not not8654(N28150,R0);
not not8655(N28151,R3);
not not8656(N28152,R4);
not not8657(N28162,R0);
not not8658(N28163,R3);
not not8659(N28164,R4);
not not8660(N28174,in1);
not not8661(N28175,R0);
not not8662(N28176,R2);
not not8663(N28177,R4);
not not8664(N28186,in1);
not not8665(N28187,in2);
not not8666(N28188,R1);
not not8667(N28198,in0);
not not8668(N28199,in1);
not not8669(N28210,in0);
not not8670(N28211,in1);
not not8671(N28212,R3);
not not8672(N28222,in1);
not not8673(N28223,R1);
not not8674(N28224,R2);
not not8675(N28234,in2);
not not8676(N28235,R1);
not not8677(N28236,R2);
not not8678(N28237,R3);
not not8679(N28246,R3);
not not8680(N28247,R4);
not not8681(N28258,R1);
not not8682(N28259,R5);
not not8683(N28270,R1);
not not8684(N28271,R5);
not not8685(N28282,in1);
not not8686(N28283,R0);
not not8687(N28284,R4);
not not8688(N28294,in0);
not not8689(N28295,in2);
not not8690(N28296,R2);
not not8691(N28297,R5);
not not8692(N28306,R2);
not not8693(N28307,R3);
not not8694(N28318,in1);
not not8695(N28319,R0);
not not8696(N28320,R1);
not not8697(N28330,in0);
not not8698(N28331,in1);
not not8699(N28332,in2);
not not8700(N28333,R3);
not not8701(N28342,in1);
not not8702(N28343,R1);
not not8703(N28344,R3);
not not8704(N28345,R4);
not not8705(N28354,R2);
not not8706(N28355,R4);
not not8707(N28356,R5);
not not8708(N28366,R1);
not not8709(N28367,R2);
not not8710(N28368,R4);
not not8711(N28378,in2);
not not8712(N28379,R0);
not not8713(N28380,R4);
not not8714(N28381,R5);
not not8715(N28390,R0);
not not8716(N28391,R2);
not not8717(N28392,R5);
not not8718(N28402,R0);
not not8719(N28403,R1);
not not8720(N28404,R3);
not not8721(N28414,in1);
not not8722(N28415,R0);
not not8723(N28416,R1);
not not8724(N28417,R4);
not not8725(N28426,R2);
not not8726(N28427,R4);
not not8727(N28438,in1);
not not8728(N28439,in2);
not not8729(N28440,R1);
not not8730(N28441,R3);
not not8731(N28450,in0);
not not8732(N28451,R0);
not not8733(N28452,R1);
not not8734(N28462,R3);
not not8735(N28463,R5);
not not8736(N28473,in1);
not not8737(N28474,R5);
not not8738(N28484,in0);
not not8739(N28485,in2);
not not8740(N28495,in2);
not not8741(N28496,R0);
not not8742(N28497,R5);
not not8743(N28506,R3);
not not8744(N28507,R5);
not not8745(N28517,R5);
not not8746(N28528,in0);
not not8747(N28529,in2);
not not8748(N28539,R0);
not not8749(N28550,R2);
not not8750(N28551,R5);
not not8751(N28561,R0);
not not8752(N28562,R1);
not not8753(N28572,in0);
not not8754(N28573,R0);
not not8755(N28583,in0);
not not8756(N28584,R0);
not not8757(N28585,R1);
not not8758(N28594,R2);
not not8759(N28595,R4);
not not8760(N28605,in2);
not not8761(N28606,R3);
not not8762(N28616,in2);
not not8763(N28617,R5);
not not8764(N28627,in1);
not not8765(N28628,R1);
not not8766(N28638,in2);
not not8767(N28639,R1);
not not8768(N28649,R1);
not not8769(N28650,R2);
not not8770(N28660,R0);
not not8771(N28661,R4);
not not8772(N28671,R1);
not not8773(N28672,R3);
not not8774(N28673,R4);
not not8775(N28682,in0);
not not8776(N28683,R3);
not not8777(N28693,in2);
not not8778(N28694,R1);
not not8779(N28703,R1);
not not8780(N28704,R3);
not not8781(N28713,R1);
not not8782(N28714,R3);
not not8783(N28723,in2);
not not8784(N28724,R4);
not not8785(N28733,R1);
not not8786(N28734,R2);
not not8787(N28743,R1);
not not8788(N28744,R4);
not not8789(N28753,R2);
not not8790(N28754,R5);
not not8791(N28763,R1);
not not8792(N28773,in1);
not not8793(N28774,R2);
not not8794(N28783,in2);
not not8795(N28784,R2);
not not8796(N28793,R0);
not not8797(N28794,R3);
not not8798(N28803,in2);
not not8799(N28804,R2);
not not8800(N28813,in1);
not not8801(N28814,R2);
not not8802(N28823,R5);
not not8803(N28833,R0);
not not8804(N28843,in1);
not not8805(N28867,in2);
not not8806(N28868,R2);
not not8807(N28869,R3);
not not8808(N28870,R5);
not not8809(N28871,R6);
not not8810(N28872,R7);
not not8811(N28880,R3);
not not8812(N28881,R4);
not not8813(N28882,R5);
not not8814(N28883,R6);
not not8815(N28884,R7);
not not8816(N28892,in1);
not not8817(N28893,R1);
not not8818(N28894,R2);
not not8819(N28895,R4);
not not8820(N28896,R5);
not not8821(N28904,in1);
not not8822(N28905,R1);
not not8823(N28906,R3);
not not8824(N28907,R6);
not not8825(N28908,R7);
not not8826(N28916,R0);
not not8827(N28917,R1);
not not8828(N28918,R4);
not not8829(N28919,R5);
not not8830(N28920,R7);
not not8831(N28928,R2);
not not8832(N28929,R4);
not not8833(N28930,R5);
not not8834(N28931,R7);
not not8835(N28939,R0);
not not8836(N28940,R1);
not not8837(N28941,R3);
not not8838(N28942,R7);
not not8839(N28950,R3);
not not8840(N28951,R4);
not not8841(N28952,R5);
not not8842(N28953,R7);
not not8843(N28961,R0);
not not8844(N28962,R4);
not not8845(N28963,R5);
not not8846(N28964,R6);
not not8847(N28972,R0);
not not8848(N28973,R5);
not not8849(N28974,R6);
not not8850(N28982,R1);
not not8851(N28983,R4);
not not8852(N28984,R7);
not not8853(N28992,R0);
not not8854(N28993,R6);
not not8855(N28994,R7);
not not8856(N29002,R2);
not not8857(N29003,R5);
not not8858(N29004,R6);
not not8859(N29012,R0);
not not8860(N29013,R1);
not not8861(N29014,R5);
not not8862(N29022,R0);
not not8863(N29023,R2);
not not8864(N29024,R6);
not not8865(N29032,R1);
not not8866(N29033,R2);
not not8867(N29034,R6);
not not8868(N29042,R1);
not not8869(N29043,R5);
not not8870(N24205,R4);
not not8871(N24206,R5);
not not8872(N24207,R6);
not not8873(N24208,R7);
not not8874(N24223,R4);
not not8875(N24224,R5);
not not8876(N24225,R6);
not not8877(N24226,R7);
not not8878(N24242,R4);
not not8879(N24243,R5);
not not8880(N24244,R7);
not not8881(N24260,R5);
not not8882(N24261,R6);
not not8883(N24262,R7);
not not8884(N24277,R4);
not not8885(N24278,R5);
not not8886(N24279,R6);
not not8887(N24280,R7);
not not8888(N24295,R4);
not not8889(N24296,R5);
not not8890(N24297,R6);
not not8891(N24298,R7);
not not8892(N24313,R4);
not not8893(N24314,R5);
not not8894(N24315,R6);
not not8895(N24316,R7);
not not8896(N24331,R4);
not not8897(N24332,R5);
not not8898(N24333,R6);
not not8899(N24348,R4);
not not8900(N24349,R5);
not not8901(N24350,R6);
not not8902(N24364,R4);
not not8903(N24365,R5);
not not8904(N24366,R6);
not not8905(N24367,R7);
not not8906(N24381,R4);
not not8907(N24382,R5);
not not8908(N24383,R6);
not not8909(N24384,R7);
not not8910(N24399,R4);
not not8911(N24400,R5);
not not8912(N24401,R6);
not not8913(N24416,R4);
not not8914(N24417,R5);
not not8915(N24418,R6);
not not8916(N24434,R3);
not not8917(N24435,R6);
not not8918(N24451,R5);
not not8919(N24452,R6);
not not8920(N24468,R4);
not not8921(N24469,R7);
not not8922(N24482,R4);
not not8923(N24483,R5);
not not8924(N24484,R6);
not not8925(N24485,R7);
not not8926(N24498,R4);
not not8927(N24499,R5);
not not8928(N24500,R6);
not not8929(N24501,R7);
not not8930(N24515,R4);
not not8931(N24516,R5);
not not8932(N24517,R7);
not not8933(N24531,R4);
not not8934(N24532,R5);
not not8935(N24533,R7);
not not8936(N24546,R4);
not not8937(N24547,R5);
not not8938(N24548,R6);
not not8939(N24549,R7);
not not8940(N24562,R4);
not not8941(N24563,R5);
not not8942(N24564,R6);
not not8943(N24565,R7);
not not8944(N24579,R4);
not not8945(N24580,R6);
not not8946(N24581,R7);
not not8947(N24595,R4);
not not8948(N24596,R6);
not not8949(N24597,R7);
not not8950(N24610,R4);
not not8951(N24611,R5);
not not8952(N24612,R6);
not not8953(N24613,R7);
not not8954(N24626,R4);
not not8955(N24627,R5);
not not8956(N24628,R6);
not not8957(N24629,R7);
not not8958(N24644,R4);
not not8959(N24645,R7);
not not8960(N24658,R4);
not not8961(N24659,R5);
not not8962(N24660,R6);
not not8963(N24661,R7);
not not8964(N24675,R3);
not not8965(N24676,R4);
not not8966(N24677,R5);
not not8967(N24691,R4);
not not8968(N24692,R5);
not not8969(N24693,R6);
not not8970(N24707,R4);
not not8971(N24708,R6);
not not8972(N24709,R7);
not not8973(N24722,R4);
not not8974(N24723,R5);
not not8975(N24724,R6);
not not8976(N24725,R7);
not not8977(N24740,R3);
not not8978(N24741,R6);
not not8979(N24755,R3);
not not8980(N24756,R6);
not not8981(N24757,R7);
not not8982(N24771,R5);
not not8983(N24772,R6);
not not8984(N24773,R7);
not not8985(N24788,R4);
not not8986(N24789,R6);
not not8987(N24804,R4);
not not8988(N24805,R5);
not not8989(N24819,R4);
not not8990(N24820,R5);
not not8991(N24821,R7);
not not8992(N24836,R5);
not not8993(N24837,R7);
not not8994(N24851,R5);
not not8995(N24852,R6);
not not8996(N24853,R7);
not not8997(N24867,R5);
not not8998(N24868,R6);
not not8999(N24869,R7);
not not9000(N24884,R4);
not not9001(N24885,R7);
not not9002(N24900,R5);
not not9003(N24901,R7);
not not9004(N24916,R5);
not not9005(N24917,R7);
not not9006(N24932,R4);
not not9007(N24933,R6);
not not9008(N24948,R5);
not not9009(N24949,R6);
not not9010(N24961,R4);
not not9011(N24962,R5);
not not9012(N24963,R6);
not not9013(N24964,R7);
not not9014(N24978,R4);
not not9015(N24979,R6);
not not9016(N24992,R4);
not not9017(N24993,R5);
not not9018(N24994,R6);
not not9019(N25007,R4);
not not9020(N25008,R5);
not not9021(N25009,R6);
not not9022(N25022,R4);
not not9023(N25023,R5);
not not9024(N25024,R6);
not not9025(N25037,R3);
not not9026(N25038,R4);
not not9027(N25039,R6);
not not9028(N25053,R3);
not not9029(N25054,R6);
not not9030(N25067,R4);
not not9031(N25068,R5);
not not9032(N25069,R6);
not not9033(N25084,R4);
not not9034(N25098,R4);
not not9035(N25099,R6);
not not9036(N25113,R4);
not not9037(N25114,R7);
not not9038(N25127,R3);
not not9039(N25128,R4);
not not9040(N25129,R7);
not not9041(N25142,R4);
not not9042(N25143,R5);
not not9043(N25144,R6);
not not9044(N25158,R4);
not not9045(N25159,R6);
not not9046(N25173,R5);
not not9047(N25174,R6);
not not9048(N25188,R5);
not not9049(N25189,R6);
not not9050(N25203,R4);
not not9051(N25204,R6);
not not9052(N25219,R4);
not not9053(N25234,R7);
not not9054(N25248,R5);
not not9055(N25249,R6);
not not9056(N25263,R6);
not not9057(N25264,R7);
not not9058(N25277,R5);
not not9059(N25278,R6);
not not9060(N25279,R7);
not not9061(N25292,R4);
not not9062(N25293,R6);
not not9063(N25294,R7);
not not9064(N25308,R4);
not not9065(N25309,R5);
not not9066(N25323,R4);
not not9067(N25324,R5);
not not9068(N25337,R4);
not not9069(N25338,R6);
not not9070(N25339,R7);
not not9071(N25353,R6);
not not9072(N25354,R7);
not not9073(N25369,R3);
not not9074(N25382,R5);
not not9075(N25383,R6);
not not9076(N25384,R7);
not not9077(N25397,R4);
not not9078(N25398,R5);
not not9079(N25399,R6);
not not9080(N25413,R4);
not not9081(N25414,R6);
not not9082(N25427,R4);
not not9083(N25428,R6);
not not9084(N25442,R6);
not not9085(N25454,R4);
not not9086(N25455,R5);
not not9087(N25456,R6);
not not9088(N25469,R4);
not not9089(N25470,R5);
not not9090(N25483,R3);
not not9091(N25484,R5);
not not9092(N25496,R3);
not not9093(N25497,R4);
not not9094(N25498,R7);
not not9095(N25512,R5);
not not9096(N25526,R6);
not not9097(N25539,R5);
not not9098(N25540,R7);
not not9099(N25553,R4);
not not9100(N25554,R5);
not not9101(N25566,R4);
not not9102(N25567,R5);
not not9103(N25568,R7);
not not9104(N25582,R7);
not not9105(N25596,R4);
not not9106(N25608,R4);
not not9107(N25609,R5);
not not9108(N25610,R6);
not not9109(N25622,R3);
not not9110(N25623,R4);
not not9111(N25624,R6);
not not9112(N25636,R4);
not not9113(N25637,R6);
not not9114(N25638,R7);
not not9115(N25651,R6);
not not9116(N25652,R7);
not not9117(N25665,R6);
not not9118(N25666,R7);
not not9119(N25693,R4);
not not9120(N25694,R5);
not not9121(N25707,R3);
not not9122(N25708,R5);
not not9123(N25720,R3);
not not9124(N25721,R5);
not not9125(N25722,R7);
not not9126(N25736,R7);
not not9127(N25748,R4);
not not9128(N25749,R5);
not not9129(N25750,R7);
not not9130(N25763,R5);
not not9131(N25764,R6);
not not9132(N25776,R4);
not not9133(N25777,R6);
not not9134(N25778,R7);
not not9135(N25791,R3);
not not9136(N25792,R4);
not not9137(N25805,R5);
not not9138(N25806,R7);
not not9139(N25819,R3);
not not9140(N25820,R7);
not not9141(N25833,R4);
not not9142(N25834,R5);
not not9143(N25846,R4);
not not9144(N25847,R5);
not not9145(N25848,R7);
not not9146(N25861,R4);
not not9147(N25862,R7);
not not9148(N25874,R3);
not not9149(N25875,R5);
not not9150(N25876,R7);
not not9151(N25888,R5);
not not9152(N25889,R6);
not not9153(N25890,R7);
not not9154(N25902,R5);
not not9155(N25903,R6);
not not9156(N25904,R7);
not not9157(N25916,R5);
not not9158(N25917,R6);
not not9159(N25918,R7);
not not9160(N25930,R3);
not not9161(N25931,R5);
not not9162(N25932,R6);
not not9163(N25944,R5);
not not9164(N25945,R6);
not not9165(N25946,R7);
not not9166(N25958,R4);
not not9167(N25959,R5);
not not9168(N25960,R6);
not not9169(N25973,R3);
not not9170(N25974,R6);
not not9171(N25987,R3);
not not9172(N25988,R6);
not not9173(N26001,R5);
not not9174(N26002,R6);
not not9175(N26014,R4);
not not9176(N26015,R6);
not not9177(N26016,R7);
not not9178(N26029,R5);
not not9179(N26030,R6);
not not9180(N26044,R4);
not not9181(N26057,R4);
not not9182(N26058,R6);
not not9183(N26072,R7);
not not9184(N26085,R4);
not not9185(N26086,R7);
not not9186(N26100,R4);
not not9187(N26111,R4);
not not9188(N26112,R5);
not not9189(N26113,R6);
not not9190(N26114,R7);
not not9191(N26127,R4);
not not9192(N26128,R5);
not not9193(N26141,R5);
not not9194(N26142,R6);
not not9195(N26156,R7);
not not9196(N26169,R4);
not not9197(N26170,R5);
not not9198(N26183,R6);
not not9199(N26196,R7);
not not9200(N26208,R4);
not not9201(N26209,R6);
not not9202(N26221,R4);
not not9203(N26222,R5);
not not9204(N26233,R4);
not not9205(N26234,R5);
not not9206(N26235,R6);
not not9207(N26246,R4);
not not9208(N26247,R5);
not not9209(N26248,R6);
not not9210(N26260,R4);
not not9211(N26261,R7);
not not9212(N26274,R4);
not not9213(N26287,R5);
not not9214(N26311,R3);
not not9215(N26312,R5);
not not9216(N26313,R6);
not not9217(N26337,R4);
not not9218(N26338,R5);
not not9219(N26339,R6);
not not9220(N26365,R4);
not not9221(N26378,R4);
not not9222(N26391,R4);
not not9223(N26403,R5);
not not9224(N26404,R7);
not not9225(N26416,R5);
not not9226(N26417,R7);
not not9227(N26430,R6);
not not9228(N26443,R6);
not not9229(N26455,R4);
not not9230(N26456,R7);
not not9231(N26468,R4);
not not9232(N26469,R5);
not not9233(N26482,R7);
not not9234(N26495,R6);
not not9235(N26507,R4);
not not9236(N26508,R5);
not not9237(N26521,R4);
not not9238(N26533,R4);
not not9239(N26534,R6);
not not9240(N26546,R4);
not not9241(N26547,R7);
not not9242(N26558,R5);
not not9243(N26559,R6);
not not9244(N26560,R7);
not not9245(N26573,R7);
not not9246(N26585,R4);
not not9247(N26586,R7);
not not9248(N26598,R4);
not not9249(N26599,R7);
not not9250(N26612,R6);
not not9251(N26623,R6);
not not9252(N26624,R7);
not not9253(N26635,R3);
not not9254(N26636,R7);
not not9255(N26648,R5);
not not9256(N26659,R4);
not not9257(N26660,R5);
not not9258(N26672,R5);
not not9259(N26683,R4);
not not9260(N26684,R6);
not not9261(N26696,R7);
not not9262(N26708,R4);
not not9263(N26719,R5);
not not9264(N26720,R7);
not not9265(N26732,R4);
not not9266(N26743,R3);
not not9267(N26744,R6);
not not9268(N26755,R4);
not not9269(N26756,R6);
not not9270(N26780,R5);
not not9271(N26792,R5);
not not9272(N26804,R4);
not not9273(N26815,R3);
not not9274(N26816,R5);
not not9275(N26828,R7);
not not9276(N26839,R4);
not not9277(N26840,R7);
not not9278(N26852,R6);
not not9279(N26863,R3);
not not9280(N26864,R5);
not not9281(N26875,R5);
not not9282(N26876,R7);
not not9283(N26899,R4);
not not9284(N26900,R7);
not not9285(N26912,R6);
not not9286(N26922,R4);
not not9287(N26923,R5);
not not9288(N26924,R6);
not not9289(N26936,R6);
not not9290(N26948,R4);
not not9291(N26960,R4);
not not9292(N26972,R4);
not not9293(N26996,R4);
not not9294(N27008,R7);
not not9295(N27020,R3);
not not9296(N27031,R4);
not not9297(N27032,R7);
not not9298(N27043,R4);
not not9299(N27044,R5);
not not9300(N27055,R4);
not not9301(N27056,R5);
not not9302(N27078,R7);
not not9303(N27100,R5);
not not9304(N27120,R4);
not not9305(N27150,R4);
not not9306(N27180,R6);
not not9307(N27190,R4);
not not9308(N27200,R4);
not not9309(N27215,R6);
not not9310(N27216,R7);
not not9311(N27231,R6);
not not9312(N27232,R7);
not not9313(N27246,R5);
not not9314(N27247,R7);
not not9315(N27261,R6);
not not9316(N27262,R7);
not not9317(N27277,R6);
not not9318(N27290,R4);
not not9319(N27291,R6);
not not9320(N27304,R6);
not not9321(N27305,R7);
not not9322(N27319,R6);
not not9323(N27333,R6);
not not9324(N27346,R6);
not not9325(N27347,R7);
not not9326(N27360,R6);
not not9327(N27361,R7);
not not9328(N27375,R7);
not not9329(N27388,R6);
not not9330(N27389,R7);
not not9331(N27403,R6);
not not9332(N27417,R7);
not not9333(N27430,R6);
not not9334(N27431,R7);
not not9335(N27445,R6);
not not9336(N27458,R6);
not not9337(N27459,R7);
not not9338(N27472,R6);
not not9339(N27473,R7);
not not9340(N27487,R5);
not not9341(N27501,R7);
not not9342(N27514,R6);
not not9343(N27515,R7);
not not9344(N27528,R5);
not not9345(N27529,R7);
not not9346(N27542,R6);
not not9347(N27543,R7);
not not9348(N27557,R7);
not not9349(N27571,R6);
not not9350(N27584,R6);
not not9351(N27585,R7);
not not9352(N27598,R6);
not not9353(N27599,R7);
not not9354(N27612,R6);
not not9355(N27624,R6);
not not9356(N27625,R7);
not not9357(N27638,R6);
not not9358(N27651,R7);
not not9359(N27664,R6);
not not9360(N27676,R6);
not not9361(N27677,R7);
not not9362(N27690,R5);
not not9363(N27702,R6);
not not9364(N27703,R7);
not not9365(N27728,R6);
not not9366(N27729,R7);
not not9367(N27741,R6);
not not9368(N27742,R7);
not not9369(N27768,R7);
not not9370(N27781,R6);
not not9371(N27794,R6);
not not9372(N27807,R6);
not not9373(N27820,R7);
not not9374(N27833,R5);
not not9375(N27845,R5);
not not9376(N27846,R6);
not not9377(N27859,R7);
not not9378(N27872,R6);
not not9379(N27898,R7);
not not9380(N27910,R6);
not not9381(N27911,R7);
not not9382(N27924,R5);
not not9383(N27937,R6);
not not9384(N27950,R6);
not not9385(N27963,R6);
not not9386(N27975,R6);
not not9387(N27976,R7);
not not9388(N27989,R5);
not not9389(N28001,R6);
not not9390(N28002,R7);
not not9391(N28014,R6);
not not9392(N28015,R7);
not not9393(N28027,R6);
not not9394(N28028,R7);
not not9395(N28041,R5);
not not9396(N28054,R7);
not not9397(N28067,R5);
not not9398(N28079,R6);
not not9399(N28080,R7);
not not9400(N28092,R6);
not not9401(N28093,R7);
not not9402(N28105,R6);
not not9403(N28116,R6);
not not9404(N28117,R7);
not not9405(N28128,R6);
not not9406(N28129,R7);
not not9407(N28141,R6);
not not9408(N28153,R7);
not not9409(N28165,R7);
not not9410(N28189,R7);
not not9411(N28200,R6);
not not9412(N28201,R7);
not not9413(N28213,R6);
not not9414(N28225,R7);
not not9415(N28248,R6);
not not9416(N28249,R7);
not not9417(N28260,R6);
not not9418(N28261,R7);
not not9419(N28272,R6);
not not9420(N28273,R7);
not not9421(N28285,R6);
not not9422(N28308,R6);
not not9423(N28309,R7);
not not9424(N28321,R7);
not not9425(N28357,R6);
not not9426(N28369,R7);
not not9427(N28393,R6);
not not9428(N28405,R5);
not not9429(N28428,R6);
not not9430(N28429,R7);
not not9431(N28453,R6);
not not9432(N28464,R6);
not not9433(N28475,R7);
not not9434(N28486,R6);
not not9435(N28508,R7);
not not9436(N28518,R6);
not not9437(N28519,R7);
not not9438(N28530,R6);
not not9439(N28540,R6);
not not9440(N28541,R7);
not not9441(N28552,R6);
not not9442(N28563,R7);
not not9443(N28574,R6);
not not9444(N28596,R6);
not not9445(N28607,R5);
not not9446(N28618,R7);
not not9447(N28629,R7);
not not9448(N28640,R7);
not not9449(N28651,R7);
not not9450(N28662,R6);
not not9451(N28684,R6);
not not9452(N28764,R5);
not not9453(N28824,R7);
not not9454(N28834,R5);
not not9455(N29226,in0);
not not9456(N29227,in2);
not not9457(N29228,R0);
not not9458(N29244,in0);
not not9459(N29245,in1);
not not9460(N29246,in2);
not not9461(N29247,R0);
not not9462(N29248,R1);
not not9463(N29262,in0);
not not9464(N29263,in1);
not not9465(N29276,in0);
not not9466(N29277,in1);
not not9467(N29278,R0);
not not9468(N29279,R2);
not not9469(N29280,R3);
not not9470(N29294,in0);
not not9471(N29295,in2);
not not9472(N29296,R0);
not not9473(N29297,R1);
not not9474(N29298,R2);
not not9475(N29312,in0);
not not9476(N29313,in2);
not not9477(N29314,R0);
not not9478(N29315,R1);
not not9479(N29316,R3);
not not9480(N29330,in0);
not not9481(N29331,in2);
not not9482(N29332,R0);
not not9483(N29333,R1);
not not9484(N29334,R2);
not not9485(N29335,R3);
not not9486(N29348,in0);
not not9487(N29349,in1);
not not9488(N29350,R0);
not not9489(N29351,R1);
not not9490(N29352,R2);
not not9491(N29366,in0);
not not9492(N29367,in2);
not not9493(N29368,R0);
not not9494(N29369,R2);
not not9495(N29370,R3);
not not9496(N29383,in0);
not not9497(N29384,R0);
not not9498(N29385,R1);
not not9499(N29386,R2);
not not9500(N29387,R3);
not not9501(N29400,in0);
not not9502(N29401,in1);
not not9503(N29402,in2);
not not9504(N29403,R2);
not not9505(N29404,R3);
not not9506(N29417,in0);
not not9507(N29418,in1);
not not9508(N29419,R1);
not not9509(N29420,R2);
not not9510(N29434,in0);
not not9511(N29435,in1);
not not9512(N29436,in2);
not not9513(N29437,R0);
not not9514(N29451,in0);
not not9515(N29452,in1);
not not9516(N29453,in2);
not not9517(N29454,R0);
not not9518(N29455,R1);
not not9519(N29468,in0);
not not9520(N29469,in1);
not not9521(N29470,R1);
not not9522(N29471,R2);
not not9523(N29472,R3);
not not9524(N29485,in0);
not not9525(N29486,in1);
not not9526(N29487,in2);
not not9527(N29488,R0);
not not9528(N29489,R1);
not not9529(N29502,in0);
not not9530(N29503,in1);
not not9531(N29504,in2);
not not9532(N29505,R0);
not not9533(N29506,R1);
not not9534(N29507,R2);
not not9535(N29519,in0);
not not9536(N29520,in2);
not not9537(N29521,R0);
not not9538(N29522,R1);
not not9539(N29523,R2);
not not9540(N29536,in0);
not not9541(N29537,R2);
not not9542(N29538,R3);
not not9543(N29552,in0);
not not9544(N29553,R0);
not not9545(N29554,R1);
not not9546(N29555,R3);
not not9547(N29568,in0);
not not9548(N29569,in1);
not not9549(N29570,R3);
not not9550(N29584,in0);
not not9551(N29585,in2);
not not9552(N29586,R2);
not not9553(N29600,in0);
not not9554(N29601,in1);
not not9555(N29602,R2);
not not9556(N29603,R3);
not not9557(N29616,in0);
not not9558(N29617,in1);
not not9559(N29618,R0);
not not9560(N29619,R1);
not not9561(N29632,in0);
not not9562(N29633,in1);
not not9563(N29634,in2);
not not9564(N29635,R2);
not not9565(N29648,in0);
not not9566(N29649,in1);
not not9567(N29650,in2);
not not9568(N29651,R1);
not not9569(N29652,R2);
not not9570(N29664,in0);
not not9571(N29665,in1);
not not9572(N29666,R0);
not not9573(N29667,R1);
not not9574(N29680,in0);
not not9575(N29681,in2);
not not9576(N29682,R0);
not not9577(N29683,R1);
not not9578(N29684,R2);
not not9579(N29696,in0);
not not9580(N29697,R0);
not not9581(N29698,R2);
not not9582(N29699,R3);
not not9583(N29712,in0);
not not9584(N29713,in1);
not not9585(N29714,R0);
not not9586(N29715,R2);
not not9587(N29728,in0);
not not9588(N29729,in2);
not not9589(N29730,R0);
not not9590(N29731,R1);
not not9591(N29744,in0);
not not9592(N29745,in1);
not not9593(N29746,in2);
not not9594(N29747,R1);
not not9595(N29748,R2);
not not9596(N29760,in0);
not not9597(N29761,in1);
not not9598(N29762,in2);
not not9599(N29763,R0);
not not9600(N29764,R1);
not not9601(N29775,in0);
not not9602(N29776,in1);
not not9603(N29777,R0);
not not9604(N29778,R1);
not not9605(N29779,R3);
not not9606(N29790,in0);
not not9607(N29791,in1);
not not9608(N29792,R1);
not not9609(N29793,R2);
not not9610(N29805,in0);
not not9611(N29806,R3);
not not9612(N29820,in0);
not not9613(N29821,in2);
not not9614(N29822,R0);
not not9615(N29823,R1);
not not9616(N29835,in0);
not not9617(N29836,in1);
not not9618(N29837,R1);
not not9619(N29838,R2);
not not9620(N29850,in0);
not not9621(N29851,in1);
not not9622(N29852,in2);
not not9623(N29853,R0);
not not9624(N29854,R1);
not not9625(N29855,R2);
not not9626(N29865,in0);
not not9627(N29866,in1);
not not9628(N29867,in2);
not not9629(N29868,R0);
not not9630(N29880,in0);
not not9631(N29881,in2);
not not9632(N29882,R0);
not not9633(N29895,in0);
not not9634(N29896,in2);
not not9635(N29897,R1);
not not9636(N29910,in0);
not not9637(N29911,R1);
not not9638(N29912,R2);
not not9639(N29913,R3);
not not9640(N29925,in0);
not not9641(N29926,in1);
not not9642(N29927,R1);
not not9643(N29940,in0);
not not9644(N29941,in1);
not not9645(N29942,R1);
not not9646(N29955,in0);
not not9647(N29956,in1);
not not9648(N29957,R2);
not not9649(N29970,in0);
not not9650(N29971,R0);
not not9651(N29972,R1);
not not9652(N29973,R2);
not not9653(N29985,in0);
not not9654(N29986,in1);
not not9655(N29987,R3);
not not9656(N30000,in0);
not not9657(N30001,in1);
not not9658(N30002,in2);
not not9659(N30015,in0);
not not9660(N30016,in2);
not not9661(N30017,R1);
not not9662(N30018,R2);
not not9663(N30030,in0);
not not9664(N30031,in1);
not not9665(N30032,R2);
not not9666(N30045,in0);
not not9667(N30046,in2);
not not9668(N30047,R2);
not not9669(N30060,in0);
not not9670(N30061,in1);
not not9671(N30062,R0);
not not9672(N30063,R2);
not not9673(N30075,in0);
not not9674(N30076,R0);
not not9675(N30077,R1);
not not9676(N30089,in0);
not not9677(N30090,in1);
not not9678(N30091,R3);
not not9679(N30103,in0);
not not9680(N30104,in1);
not not9681(N30105,R0);
not not9682(N30117,in0);
not not9683(N30118,in2);
not not9684(N30119,R0);
not not9685(N30131,in0);
not not9686(N30132,R3);
not not9687(N30145,in0);
not not9688(N30146,in1);
not not9689(N30147,in2);
not not9690(N30148,R1);
not not9691(N30159,in0);
not not9692(N30160,in2);
not not9693(N30173,in0);
not not9694(N30174,in2);
not not9695(N30175,R0);
not not9696(N30187,in0);
not not9697(N30188,R0);
not not9698(N30201,in0);
not not9699(N30202,R1);
not not9700(N30215,in0);
not not9701(N30216,R1);
not not9702(N30217,R2);
not not9703(N30229,in0);
not not9704(N30230,R1);
not not9705(N30231,R3);
not not9706(N30243,in0);
not not9707(N30244,in1);
not not9708(N30245,in2);
not not9709(N30246,R1);
not not9710(N30257,in0);
not not9711(N30258,in1);
not not9712(N30259,R0);
not not9713(N30271,in0);
not not9714(N30272,in1);
not not9715(N30273,R2);
not not9716(N30285,in0);
not not9717(N30286,in1);
not not9718(N30287,in2);
not not9719(N30288,R2);
not not9720(N30299,in0);
not not9721(N30300,in1);
not not9722(N30301,R0);
not not9723(N30313,in0);
not not9724(N30314,R2);
not not9725(N30327,in0);
not not9726(N30328,in2);
not not9727(N30329,R0);
not not9728(N30341,in0);
not not9729(N30342,in2);
not not9730(N30343,R0);
not not9731(N30355,in0);
not not9732(N30356,in2);
not not9733(N30357,R1);
not not9734(N30369,in0);
not not9735(N30370,in1);
not not9736(N30371,in2);
not not9737(N30372,R0);
not not9738(N30383,in0);
not not9739(N30384,in1);
not not9740(N30397,in0);
not not9741(N30398,in2);
not not9742(N30399,R1);
not not9743(N30400,R3);
not not9744(N30411,in0);
not not9745(N30412,in1);
not not9746(N30413,in2);
not not9747(N30425,in0);
not not9748(N30426,in2);
not not9749(N30427,R1);
not not9750(N30428,R2);
not not9751(N30439,in0);
not not9752(N30440,in1);
not not9753(N30441,in2);
not not9754(N30442,R1);
not not9755(N30443,R3);
not not9756(N30453,in0);
not not9757(N30454,in1);
not not9758(N30455,in2);
not not9759(N30456,R0);
not not9760(N30457,R2);
not not9761(N30467,in0);
not not9762(N30468,R0);
not not9763(N30481,in0);
not not9764(N30482,R0);
not not9765(N30483,R1);
not not9766(N30495,in0);
not not9767(N30496,in1);
not not9768(N30497,R1);
not not9769(N30509,in0);
not not9770(N30510,in1);
not not9771(N30511,R0);
not not9772(N30512,R1);
not not9773(N30523,in0);
not not9774(N30524,R1);
not not9775(N30525,R2);
not not9776(N30537,in0);
not not9777(N30538,in2);
not not9778(N30539,R0);
not not9779(N30551,in0);
not not9780(N30552,in2);
not not9781(N30553,R0);
not not9782(N30554,R1);
not not9783(N30555,R2);
not not9784(N30565,in0);
not not9785(N30566,in1);
not not9786(N30567,R0);
not not9787(N30568,R1);
not not9788(N30579,in0);
not not9789(N30580,in1);
not not9790(N30581,R3);
not not9791(N30593,in0);
not not9792(N30594,in2);
not not9793(N30595,R1);
not not9794(N30607,in0);
not not9795(N30608,in1);
not not9796(N30609,R3);
not not9797(N30621,in0);
not not9798(N30622,in2);
not not9799(N30623,R1);
not not9800(N30635,in0);
not not9801(N30636,in2);
not not9802(N30637,R0);
not not9803(N30649,in0);
not not9804(N30650,R0);
not not9805(N30651,R1);
not not9806(N30663,in0);
not not9807(N30664,in1);
not not9808(N30677,in0);
not not9809(N30678,in1);
not not9810(N30679,in2);
not not9811(N30680,R2);
not not9812(N30691,in0);
not not9813(N30692,in1);
not not9814(N30705,in0);
not not9815(N30706,R2);
not not9816(N30719,in0);
not not9817(N30720,in2);
not not9818(N30732,in0);
not not9819(N30733,R0);
not not9820(N30734,R1);
not not9821(N30745,in0);
not not9822(N30746,R0);
not not9823(N30758,in0);
not not9824(N30759,in1);
not not9825(N30760,in2);
not not9826(N30771,in0);
not not9827(N30772,R1);
not not9828(N30784,in0);
not not9829(N30785,in2);
not not9830(N30786,R1);
not not9831(N30797,in0);
not not9832(N30798,in1);
not not9833(N30799,R0);
not not9834(N30800,R2);
not not9835(N30810,in0);
not not9836(N30811,in1);
not not9837(N30812,R1);
not not9838(N30823,in0);
not not9839(N30836,in0);
not not9840(N30837,in2);
not not9841(N30838,R1);
not not9842(N30849,in0);
not not9843(N30850,R1);
not not9844(N30851,R2);
not not9845(N30862,in0);
not not9846(N30863,R2);
not not9847(N30875,in0);
not not9848(N30876,in1);
not not9849(N30888,in0);
not not9850(N30889,R0);
not not9851(N30901,in0);
not not9852(N30902,in1);
not not9853(N30914,in0);
not not9854(N30915,R2);
not not9855(N30927,in0);
not not9856(N30940,in0);
not not9857(N30953,in0);
not not9858(N30954,R1);
not not9859(N30955,R3);
not not9860(N30966,in0);
not not9861(N30967,in2);
not not9862(N30979,in0);
not not9863(N30980,in1);
not not9864(N30981,in2);
not not9865(N30992,in0);
not not9866(N30993,in2);
not not9867(N31005,in0);
not not9868(N31006,in1);
not not9869(N31018,in0);
not not9870(N31019,R3);
not not9871(N31031,in0);
not not9872(N31032,R0);
not not9873(N31043,in0);
not not9874(N31044,R0);
not not9875(N31055,in0);
not not9876(N31056,in1);
not not9877(N31057,R1);
not not9878(N31067,in0);
not not9879(N31068,in1);
not not9880(N31069,R1);
not not9881(N31079,in0);
not not9882(N31080,R1);
not not9883(N31091,in0);
not not9884(N31092,in2);
not not9885(N31103,in0);
not not9886(N31104,in1);
not not9887(N31105,R1);
not not9888(N31115,in0);
not not9889(N31116,in1);
not not9890(N31127,in0);
not not9891(N31128,R1);
not not9892(N31139,in0);
not not9893(N31140,R0);
not not9894(N31141,R2);
not not9895(N31151,in0);
not not9896(N31152,R1);
not not9897(N31163,in0);
not not9898(N31164,in1);
not not9899(N31175,in0);
not not9900(N31176,in1);
not not9901(N31187,in0);
not not9902(N31188,R0);
not not9903(N31189,R1);
not not9904(N31199,in0);
not not9905(N31200,in1);
not not9906(N31201,R1);
not not9907(N31211,in0);
not not9908(N31212,R0);
not not9909(N31222,in0);
not not9910(N31233,in0);
not not9911(N31234,in1);
not not9912(N31243,in0);
not not9913(N31244,R1);
not not9914(N31245,R3);
not not9915(N31246,R4);
not not9916(N31247,R5);
not not9917(N31258,in0);
not not9918(N31259,in2);
not not9919(N31260,R1);
not not9920(N31261,R2);
not not9921(N31262,R4);
not not9922(N31273,in0);
not not9923(N31274,in2);
not not9924(N31275,R1);
not not9925(N31276,R2);
not not9926(N31277,R3);
not not9927(N31278,R4);
not not9928(N31288,in0);
not not9929(N31289,in1);
not not9930(N31290,R1);
not not9931(N31291,R3);
not not9932(N31292,R4);
not not9933(N31303,in0);
not not9934(N31304,R1);
not not9935(N31305,R3);
not not9936(N31306,R4);
not not9937(N31307,R5);
not not9938(N31317,in0);
not not9939(N31318,in1);
not not9940(N31319,R1);
not not9941(N31320,R2);
not not9942(N31321,R3);
not not9943(N31331,in0);
not not9944(N31332,in1);
not not9945(N31333,R2);
not not9946(N31334,R3);
not not9947(N31335,R4);
not not9948(N31345,in0);
not not9949(N31346,in2);
not not9950(N31347,R1);
not not9951(N31348,R2);
not not9952(N31349,R3);
not not9953(N31350,R4);
not not9954(N31359,in0);
not not9955(N31360,in2);
not not9956(N31361,R1);
not not9957(N31362,R2);
not not9958(N31363,R3);
not not9959(N31373,in0);
not not9960(N31374,in2);
not not9961(N31375,R1);
not not9962(N31376,R3);
not not9963(N31377,R4);
not not9964(N31378,R5);
not not9965(N31387,in0);
not not9966(N31388,in2);
not not9967(N31389,R3);
not not9968(N31390,R4);
not not9969(N31401,in0);
not not9970(N31402,in1);
not not9971(N31403,R3);
not not9972(N31414,in0);
not not9973(N31415,R1);
not not9974(N31416,R2);
not not9975(N31417,R4);
not not9976(N31427,in0);
not not9977(N31428,in2);
not not9978(N31429,R4);
not not9979(N31440,in0);
not not9980(N31441,in1);
not not9981(N31442,in2);
not not9982(N31443,R1);
not not9983(N31453,in0);
not not9984(N31454,in1);
not not9985(N31455,in2);
not not9986(N31456,R1);
not not9987(N31457,R3);
not not9988(N31466,in0);
not not9989(N31467,in1);
not not9990(N31468,R4);
not not9991(N31479,in0);
not not9992(N31480,in1);
not not9993(N31481,in2);
not not9994(N31482,R3);
not not9995(N31492,in0);
not not9996(N31493,R1);
not not9997(N31494,R3);
not not9998(N31495,R4);
not not9999(N31504,in0);
not not10000(N31505,R1);
not not10001(N31506,R3);
not not10002(N31507,R4);
not not10003(N31516,in0);
not not10004(N31517,in2);
not not10005(N31518,R2);
not not10006(N31519,R4);
not not10007(N31528,in0);
not not10008(N31529,R2);
not not10009(N31540,in0);
not not10010(N31541,R3);
not not10011(N31542,R4);
not not10012(N31551,in0);
not not10013(N31552,R0);
not not10014(N31562,in0);
not not10015(N31563,R4);
not not10016(N29229,R2);
not not10017(N29230,R4);
not not10018(N29231,R5);
not not10019(N29232,R6);
not not10020(N29233,R7);
not not10021(N29249,R3);
not not10022(N29250,R5);
not not10023(N29251,R7);
not not10024(N29264,R2);
not not10025(N29265,R5);
not not10026(N29266,R6);
not not10027(N29281,R4);
not not10028(N29282,R5);
not not10029(N29283,R6);
not not10030(N29284,R7);
not not10031(N29299,R3);
not not10032(N29300,R5);
not not10033(N29301,R6);
not not10034(N29302,R7);
not not10035(N29317,R4);
not not10036(N29318,R5);
not not10037(N29319,R6);
not not10038(N29320,R7);
not not10039(N29336,R4);
not not10040(N29337,R6);
not not10041(N29338,R7);
not not10042(N29353,R3);
not not10043(N29354,R4);
not not10044(N29355,R5);
not not10045(N29356,R7);
not not10046(N29371,R4);
not not10047(N29372,R5);
not not10048(N29373,R6);
not not10049(N29388,R5);
not not10050(N29389,R6);
not not10051(N29390,R7);
not not10052(N29405,R5);
not not10053(N29406,R6);
not not10054(N29407,R7);
not not10055(N29421,R4);
not not10056(N29422,R5);
not not10057(N29423,R6);
not not10058(N29424,R7);
not not10059(N29438,R4);
not not10060(N29439,R5);
not not10061(N29440,R6);
not not10062(N29441,R7);
not not10063(N29456,R3);
not not10064(N29457,R6);
not not10065(N29458,R7);
not not10066(N29473,R4);
not not10067(N29474,R5);
not not10068(N29475,R6);
not not10069(N29490,R4);
not not10070(N29491,R5);
not not10071(N29492,R6);
not not10072(N29508,R6);
not not10073(N29509,R7);
not not10074(N29524,R4);
not not10075(N29525,R5);
not not10076(N29526,R6);
not not10077(N29539,R4);
not not10078(N29540,R5);
not not10079(N29541,R6);
not not10080(N29542,R7);
not not10081(N29556,R4);
not not10082(N29557,R6);
not not10083(N29558,R7);
not not10084(N29571,R4);
not not10085(N29572,R5);
not not10086(N29573,R6);
not not10087(N29574,R7);
not not10088(N29587,R3);
not not10089(N29588,R4);
not not10090(N29589,R5);
not not10091(N29590,R6);
not not10092(N29604,R4);
not not10093(N29605,R5);
not not10094(N29606,R6);
not not10095(N29620,R3);
not not10096(N29621,R4);
not not10097(N29622,R7);
not not10098(N29636,R5);
not not10099(N29637,R6);
not not10100(N29638,R7);
not not10101(N29653,R4);
not not10102(N29654,R5);
not not10103(N29668,R5);
not not10104(N29669,R6);
not not10105(N29670,R7);
not not10106(N29685,R5);
not not10107(N29686,R7);
not not10108(N29700,R4);
not not10109(N29701,R6);
not not10110(N29702,R7);
not not10111(N29716,R4);
not not10112(N29717,R5);
not not10113(N29718,R6);
not not10114(N29732,R5);
not not10115(N29733,R6);
not not10116(N29734,R7);
not not10117(N29749,R4);
not not10118(N29750,R5);
not not10119(N29765,R4);
not not10120(N29780,R6);
not not10121(N29794,R6);
not not10122(N29795,R7);
not not10123(N29807,R4);
not not10124(N29808,R5);
not not10125(N29809,R6);
not not10126(N29810,R7);
not not10127(N29824,R5);
not not10128(N29825,R7);
not not10129(N29839,R6);
not not10130(N29840,R7);
not not10131(N29869,R4);
not not10132(N29870,R5);
not not10133(N29883,R3);
not not10134(N29884,R4);
not not10135(N29885,R7);
not not10136(N29898,R3);
not not10137(N29899,R6);
not not10138(N29900,R7);
not not10139(N29914,R5);
not not10140(N29915,R7);
not not10141(N29928,R5);
not not10142(N29929,R6);
not not10143(N29930,R7);
not not10144(N29943,R3);
not not10145(N29944,R6);
not not10146(N29945,R7);
not not10147(N29958,R3);
not not10148(N29959,R6);
not not10149(N29960,R7);
not not10150(N29974,R4);
not not10151(N29975,R5);
not not10152(N29988,R4);
not not10153(N29989,R5);
not not10154(N29990,R7);
not not10155(N30003,R4);
not not10156(N30004,R5);
not not10157(N30005,R6);
not not10158(N30019,R4);
not not10159(N30020,R6);
not not10160(N30033,R4);
not not10161(N30034,R6);
not not10162(N30035,R7);
not not10163(N30048,R5);
not not10164(N30049,R6);
not not10165(N30050,R7);
not not10166(N30064,R6);
not not10167(N30065,R7);
not not10168(N30078,R4);
not not10169(N30079,R6);
not not10170(N30092,R4);
not not10171(N30093,R7);
not not10172(N30106,R4);
not not10173(N30107,R5);
not not10174(N30120,R4);
not not10175(N30121,R5);
not not10176(N30133,R4);
not not10177(N30134,R5);
not not10178(N30135,R7);
not not10179(N30149,R3);
not not10180(N30161,R4);
not not10181(N30162,R5);
not not10182(N30163,R6);
not not10183(N30176,R5);
not not10184(N30177,R6);
not not10185(N30189,R4);
not not10186(N30190,R6);
not not10187(N30191,R7);
not not10188(N30203,R4);
not not10189(N30204,R5);
not not10190(N30205,R6);
not not10191(N30218,R5);
not not10192(N30219,R7);
not not10193(N30232,R5);
not not10194(N30233,R7);
not not10195(N30247,R5);
not not10196(N30260,R3);
not not10197(N30261,R6);
not not10198(N30274,R5);
not not10199(N30275,R7);
not not10200(N30289,R5);
not not10201(N30302,R4);
not not10202(N30303,R7);
not not10203(N30315,R3);
not not10204(N30316,R5);
not not10205(N30317,R6);
not not10206(N30330,R5);
not not10207(N30331,R6);
not not10208(N30344,R4);
not not10209(N30345,R7);
not not10210(N30358,R4);
not not10211(N30359,R7);
not not10212(N30373,R6);
not not10213(N30385,R5);
not not10214(N30386,R6);
not not10215(N30387,R7);
not not10216(N30401,R6);
not not10217(N30414,R3);
not not10218(N30415,R4);
not not10219(N30429,R7);
not not10220(N30469,R3);
not not10221(N30470,R6);
not not10222(N30471,R7);
not not10223(N30484,R5);
not not10224(N30485,R6);
not not10225(N30498,R4);
not not10226(N30499,R5);
not not10227(N30513,R6);
not not10228(N30526,R6);
not not10229(N30527,R7);
not not10230(N30540,R4);
not not10231(N30541,R5);
not not10232(N30569,R6);
not not10233(N30582,R5);
not not10234(N30583,R6);
not not10235(N30596,R4);
not not10236(N30597,R7);
not not10237(N30610,R5);
not not10238(N30611,R6);
not not10239(N30624,R3);
not not10240(N30625,R6);
not not10241(N30638,R5);
not not10242(N30639,R6);
not not10243(N30652,R5);
not not10244(N30653,R6);
not not10245(N30665,R4);
not not10246(N30666,R5);
not not10247(N30667,R6);
not not10248(N30681,R7);
not not10249(N30693,R4);
not not10250(N30694,R5);
not not10251(N30695,R7);
not not10252(N30707,R3);
not not10253(N30708,R6);
not not10254(N30709,R7);
not not10255(N30721,R6);
not not10256(N30722,R7);
not not10257(N30735,R5);
not not10258(N30747,R5);
not not10259(N30748,R6);
not not10260(N30761,R4);
not not10261(N30773,R4);
not not10262(N30774,R5);
not not10263(N30787,R4);
not not10264(N30813,R7);
not not10265(N30824,R4);
not not10266(N30825,R6);
not not10267(N30826,R7);
not not10268(N30839,R6);
not not10269(N30852,R4);
not not10270(N30864,R4);
not not10271(N30865,R6);
not not10272(N30877,R6);
not not10273(N30878,R7);
not not10274(N30890,R4);
not not10275(N30891,R6);
not not10276(N30903,R3);
not not10277(N30904,R7);
not not10278(N30916,R5);
not not10279(N30917,R7);
not not10280(N30928,R3);
not not10281(N30929,R5);
not not10282(N30930,R7);
not not10283(N30941,R5);
not not10284(N30942,R6);
not not10285(N30943,R7);
not not10286(N30956,R6);
not not10287(N30968,R4);
not not10288(N30969,R7);
not not10289(N30982,R6);
not not10290(N30994,R3);
not not10291(N30995,R6);
not not10292(N31007,R3);
not not10293(N31008,R6);
not not10294(N31020,R5);
not not10295(N31021,R6);
not not10296(N31033,R7);
not not10297(N31045,R7);
not not10298(N31081,R5);
not not10299(N31093,R5);
not not10300(N31117,R4);
not not10301(N31129,R5);
not not10302(N31153,R5);
not not10303(N31165,R5);
not not10304(N31177,R4);
not not10305(N31223,R5);
not not10306(N31248,R6);
not not10307(N31249,R7);
not not10308(N31263,R6);
not not10309(N31264,R7);
not not10310(N31279,R6);
not not10311(N31293,R6);
not not10312(N31294,R7);
not not10313(N31308,R6);
not not10314(N31322,R4);
not not10315(N31336,R6);
not not10316(N31364,R6);
not not10317(N31391,R6);
not not10318(N31392,R7);
not not10319(N31404,R6);
not not10320(N31405,R7);
not not10321(N31418,R7);
not not10322(N31430,R6);
not not10323(N31431,R7);
not not10324(N31444,R5);
not not10325(N31469,R6);
not not10326(N31470,R7);
not not10327(N31483,R6);
not not10328(N31530,R4);
not not10329(N31531,R5);
not not10330(N31553,R7);
not not10331(N31794,in0);
not not10332(N31795,R0);
not not10333(N31808,in0);
not not10334(N31809,in1);
not not10335(N31810,in2);
not not10336(N31811,R0);
not not10337(N31812,R2);
not not10338(N31826,in1);
not not10339(N31827,in2);
not not10340(N31828,R0);
not not10341(N31829,R1);
not not10342(N31830,R2);
not not10343(N31831,R3);
not not10344(N31844,in0);
not not10345(N31845,in2);
not not10346(N31846,R0);
not not10347(N31847,R1);
not not10348(N31848,R2);
not not10349(N31862,in0);
not not10350(N31863,in1);
not not10351(N31864,in2);
not not10352(N31865,R0);
not not10353(N31866,R1);
not not10354(N31880,in0);
not not10355(N31881,in2);
not not10356(N31882,R0);
not not10357(N31883,R1);
not not10358(N31884,R2);
not not10359(N31885,R3);
not not10360(N31898,in0);
not not10361(N31899,in2);
not not10362(N31900,R0);
not not10363(N31901,R1);
not not10364(N31902,R2);
not not10365(N31916,in0);
not not10366(N31917,in1);
not not10367(N31918,in2);
not not10368(N31919,R1);
not not10369(N31920,R2);
not not10370(N31921,R3);
not not10371(N31934,in0);
not not10372(N31935,R1);
not not10373(N31936,R2);
not not10374(N31937,R3);
not not10375(N31951,in0);
not not10376(N31952,in1);
not not10377(N31953,R0);
not not10378(N31954,R2);
not not10379(N31955,R3);
not not10380(N31968,in0);
not not10381(N31969,in1);
not not10382(N31970,in2);
not not10383(N31971,R0);
not not10384(N31972,R2);
not not10385(N31973,R3);
not not10386(N31985,in0);
not not10387(N31986,in1);
not not10388(N31987,R1);
not not10389(N31988,R2);
not not10390(N31989,R3);
not not10391(N32002,in0);
not not10392(N32003,in1);
not not10393(N32004,in2);
not not10394(N32005,R0);
not not10395(N32006,R1);
not not10396(N32007,R2);
not not10397(N32019,in0);
not not10398(N32020,in1);
not not10399(N32021,in2);
not not10400(N32022,R0);
not not10401(N32023,R1);
not not10402(N32024,R2);
not not10403(N32036,in0);
not not10404(N32037,R2);
not not10405(N32038,R3);
not not10406(N32052,R0);
not not10407(N32053,R1);
not not10408(N32054,R2);
not not10409(N32055,R3);
not not10410(N32068,R0);
not not10411(N32069,R1);
not not10412(N32070,R2);
not not10413(N32071,R3);
not not10414(N32084,in0);
not not10415(N32085,in1);
not not10416(N32086,R1);
not not10417(N32087,R2);
not not10418(N32100,in0);
not not10419(N32101,in1);
not not10420(N32102,R1);
not not10421(N32103,R2);
not not10422(N32116,in0);
not not10423(N32117,in2);
not not10424(N32118,R0);
not not10425(N32119,R2);
not not10426(N32132,in0);
not not10427(N32133,R0);
not not10428(N32134,R1);
not not10429(N32135,R3);
not not10430(N32148,in0);
not not10431(N32149,in1);
not not10432(N32150,in2);
not not10433(N32151,R0);
not not10434(N32164,in0);
not not10435(N32165,in1);
not not10436(N32166,R0);
not not10437(N32167,R1);
not not10438(N32168,R2);
not not10439(N32180,in0);
not not10440(N32181,in1);
not not10441(N32182,R2);
not not10442(N32183,R3);
not not10443(N32196,in0);
not not10444(N32197,in2);
not not10445(N32198,R1);
not not10446(N32199,R2);
not not10447(N32212,in0);
not not10448(N32213,in1);
not not10449(N32214,in2);
not not10450(N32215,R1);
not not10451(N32228,in0);
not not10452(N32229,R0);
not not10453(N32230,R1);
not not10454(N32244,in0);
not not10455(N32245,in1);
not not10456(N32246,R0);
not not10457(N32247,R1);
not not10458(N32260,in0);
not not10459(N32261,in2);
not not10460(N32262,R0);
not not10461(N32263,R1);
not not10462(N32276,in0);
not not10463(N32277,R0);
not not10464(N32278,R1);
not not10465(N32279,R3);
not not10466(N32292,in0);
not not10467(N32293,in2);
not not10468(N32294,R0);
not not10469(N32295,R1);
not not10470(N32296,R2);
not not10471(N32308,in0);
not not10472(N32309,in1);
not not10473(N32310,in2);
not not10474(N32311,R0);
not not10475(N32312,R1);
not not10476(N32324,in0);
not not10477(N32325,in2);
not not10478(N32326,R1);
not not10479(N32327,R2);
not not10480(N32340,in0);
not not10481(N32341,in1);
not not10482(N32342,in2);
not not10483(N32343,R1);
not not10484(N32344,R2);
not not10485(N32356,in0);
not not10486(N32357,in1);
not not10487(N32358,R0);
not not10488(N32359,R1);
not not10489(N32372,in0);
not not10490(N32373,in2);
not not10491(N32374,R1);
not not10492(N32375,R2);
not not10493(N32388,in0);
not not10494(N32389,in1);
not not10495(N32390,in2);
not not10496(N32391,R1);
not not10497(N32404,in0);
not not10498(N32405,in1);
not not10499(N32406,in2);
not not10500(N32407,R2);
not not10501(N32420,in0);
not not10502(N32421,in2);
not not10503(N32422,R0);
not not10504(N32423,R1);
not not10505(N32424,R2);
not not10506(N32436,in0);
not not10507(N32437,in2);
not not10508(N32438,R1);
not not10509(N32439,R2);
not not10510(N32440,R3);
not not10511(N32451,in0);
not not10512(N32452,in1);
not not10513(N32466,in0);
not not10514(N32467,R0);
not not10515(N32481,in0);
not not10516(N32482,R1);
not not10517(N32496,in0);
not not10518(N32497,in2);
not not10519(N32498,R2);
not not10520(N32511,in0);
not not10521(N32512,R1);
not not10522(N32513,R2);
not not10523(N32526,in0);
not not10524(N32527,R1);
not not10525(N32528,R2);
not not10526(N32529,R3);
not not10527(N32541,in0);
not not10528(N32542,in1);
not not10529(N32543,in2);
not not10530(N32544,R2);
not not10531(N32556,in0);
not not10532(N32557,in1);
not not10533(N32558,R2);
not not10534(N32571,in0);
not not10535(N32572,R0);
not not10536(N32573,R1);
not not10537(N32586,in0);
not not10538(N32587,R0);
not not10539(N32588,R1);
not not10540(N32589,R2);
not not10541(N32601,in0);
not not10542(N32602,R2);
not not10543(N32603,R3);
not not10544(N32616,in0);
not not10545(N32617,in1);
not not10546(N32618,in2);
not not10547(N32619,R0);
not not10548(N32631,in0);
not not10549(N32632,in2);
not not10550(N32633,R1);
not not10551(N32634,R3);
not not10552(N32646,in0);
not not10553(N32647,in1);
not not10554(N32648,R0);
not not10555(N32649,R1);
not not10556(N32661,in0);
not not10557(N32662,in1);
not not10558(N32663,in2);
not not10559(N32664,R0);
not not10560(N32665,R1);
not not10561(N32666,R2);
not not10562(N32676,in0);
not not10563(N32677,in2);
not not10564(N32678,R1);
not not10565(N32691,in0);
not not10566(N32692,in1);
not not10567(N32693,R1);
not not10568(N32694,R2);
not not10569(N32706,in0);
not not10570(N32707,in2);
not not10571(N32708,R2);
not not10572(N32721,in0);
not not10573(N32722,R2);
not not10574(N32736,in0);
not not10575(N32737,in1);
not not10576(N32738,in2);
not not10577(N32739,R0);
not not10578(N32740,R1);
not not10579(N32751,in0);
not not10580(N32752,in1);
not not10581(N32753,in2);
not not10582(N32754,R2);
not not10583(N32766,in0);
not not10584(N32767,in2);
not not10585(N32768,R2);
not not10586(N32781,in0);
not not10587(N32782,in1);
not not10588(N32783,R0);
not not10589(N32784,R1);
not not10590(N32796,in0);
not not10591(N32797,in1);
not not10592(N32798,in2);
not not10593(N32799,R1);
not not10594(N32811,in0);
not not10595(N32812,in2);
not not10596(N32826,in0);
not not10597(N32827,in2);
not not10598(N32828,R0);
not not10599(N32829,R1);
not not10600(N32840,in0);
not not10601(N32841,in2);
not not10602(N32842,R0);
not not10603(N32854,in0);
not not10604(N32855,in1);
not not10605(N32856,R0);
not not10606(N32868,in0);
not not10607(N32869,in1);
not not10608(N32870,in2);
not not10609(N32871,R0);
not not10610(N32882,in0);
not not10611(N32883,R0);
not not10612(N32896,in0);
not not10613(N32897,R1);
not not10614(N32898,R2);
not not10615(N32910,in0);
not not10616(N32911,R0);
not not10617(N32912,R1);
not not10618(N32924,in0);
not not10619(N32925,in2);
not not10620(N32926,R0);
not not10621(N32927,R1);
not not10622(N32928,R2);
not not10623(N32938,in0);
not not10624(N32939,R0);
not not10625(N32940,R3);
not not10626(N32952,in0);
not not10627(N32953,in1);
not not10628(N32954,R0);
not not10629(N32966,in0);
not not10630(N32967,in1);
not not10631(N32968,R2);
not not10632(N32980,in0);
not not10633(N32981,in1);
not not10634(N32982,R3);
not not10635(N32994,in0);
not not10636(N32995,R3);
not not10637(N33008,in0);
not not10638(N33009,in2);
not not10639(N33010,R0);
not not10640(N33011,R1);
not not10641(N33012,R3);
not not10642(N33022,in0);
not not10643(N33023,in1);
not not10644(N33036,in0);
not not10645(N33037,in2);
not not10646(N33038,R1);
not not10647(N33039,R2);
not not10648(N33050,in0);
not not10649(N33051,in1);
not not10650(N33052,R0);
not not10651(N33053,R3);
not not10652(N33064,in0);
not not10653(N33065,R0);
not not10654(N33066,R1);
not not10655(N33078,in0);
not not10656(N33079,in1);
not not10657(N33080,in2);
not not10658(N33081,R2);
not not10659(N33092,in0);
not not10660(N33093,in2);
not not10661(N33094,R2);
not not10662(N33106,in0);
not not10663(N33107,in1);
not not10664(N33108,R3);
not not10665(N33120,in0);
not not10666(N33121,R1);
not not10667(N33122,R2);
not not10668(N33134,in0);
not not10669(N33135,in2);
not not10670(N33136,R2);
not not10671(N33148,in0);
not not10672(N33149,R1);
not not10673(N33150,R2);
not not10674(N33151,R3);
not not10675(N33162,in0);
not not10676(N33163,in1);
not not10677(N33164,in2);
not not10678(N33165,R1);
not not10679(N33166,R2);
not not10680(N33176,in0);
not not10681(N33177,in2);
not not10682(N33178,R1);
not not10683(N33190,in0);
not not10684(N33191,in2);
not not10685(N33192,R0);
not not10686(N33204,in0);
not not10687(N33205,R1);
not not10688(N33206,R2);
not not10689(N33218,in0);
not not10690(N33219,in2);
not not10691(N33220,R2);
not not10692(N33232,in0);
not not10693(N33233,R1);
not not10694(N33234,R2);
not not10695(N33246,in0);
not not10696(N33247,in2);
not not10697(N33248,R0);
not not10698(N33249,R1);
not not10699(N33260,in0);
not not10700(N33261,R1);
not not10701(N33262,R2);
not not10702(N33274,in0);
not not10703(N33275,in1);
not not10704(N33276,in2);
not not10705(N33277,R2);
not not10706(N33288,in0);
not not10707(N33289,in1);
not not10708(N33290,R0);
not not10709(N33291,R1);
not not10710(N33302,in0);
not not10711(N33303,in2);
not not10712(N33304,R1);
not not10713(N33305,R2);
not not10714(N33316,in0);
not not10715(N33317,in2);
not not10716(N33318,R1);
not not10717(N33319,R2);
not not10718(N33330,in0);
not not10719(N33331,in2);
not not10720(N33332,R0);
not not10721(N33333,R1);
not not10722(N33344,in0);
not not10723(N33345,in2);
not not10724(N33346,R0);
not not10725(N33347,R1);
not not10726(N33358,in0);
not not10727(N33359,in1);
not not10728(N33360,R0);
not not10729(N33361,R1);
not not10730(N33372,in0);
not not10731(N33373,in2);
not not10732(N33374,R1);
not not10733(N33386,in0);
not not10734(N33387,in2);
not not10735(N33388,R2);
not not10736(N33400,in0);
not not10737(N33401,R1);
not not10738(N33402,R3);
not not10739(N33414,in1);
not not10740(N33415,in2);
not not10741(N33416,R1);
not not10742(N33427,in0);
not not10743(N33428,in1);
not not10744(N33429,R1);
not not10745(N33440,in0);
not not10746(N33441,in1);
not not10747(N33442,R0);
not not10748(N33453,in0);
not not10749(N33454,in1);
not not10750(N33455,in2);
not not10751(N33466,in0);
not not10752(N33467,in2);
not not10753(N33479,in0);
not not10754(N33480,R1);
not not10755(N33481,R2);
not not10756(N33492,in0);
not not10757(N33493,R0);
not not10758(N33505,in0);
not not10759(N33506,in1);
not not10760(N33518,in0);
not not10761(N33519,in1);
not not10762(N33520,in2);
not not10763(N33531,in0);
not not10764(N33532,R0);
not not10765(N33544,in0);
not not10766(N33545,in1);
not not10767(N33557,in0);
not not10768(N33558,in2);
not not10769(N33559,R1);
not not10770(N33570,in1);
not not10771(N33571,R1);
not not10772(N33583,in0);
not not10773(N33584,in1);
not not10774(N33585,R1);
not not10775(N33586,R3);
not not10776(N33596,in0);
not not10777(N33597,in1);
not not10778(N33598,R0);
not not10779(N33599,R2);
not not10780(N33609,R3);
not not10781(N33622,in0);
not not10782(N33623,R0);
not not10783(N33635,in1);
not not10784(N33636,in2);
not not10785(N33637,R3);
not not10786(N33648,in0);
not not10787(N33649,R1);
not not10788(N33650,R2);
not not10789(N33661,in0);
not not10790(N33662,R0);
not not10791(N33663,R1);
not not10792(N33674,in0);
not not10793(N33675,in2);
not not10794(N33676,R3);
not not10795(N33687,in0);
not not10796(N33688,R2);
not not10797(N33700,in0);
not not10798(N33701,in1);
not not10799(N33702,R0);
not not10800(N33703,R1);
not not10801(N33713,in0);
not not10802(N33714,in1);
not not10803(N33715,R2);
not not10804(N33726,in0);
not not10805(N33727,R0);
not not10806(N33738,in0);
not not10807(N33739,R1);
not not10808(N33750,in0);
not not10809(N33751,in2);
not not10810(N33762,in0);
not not10811(N33763,in1);
not not10812(N33774,in0);
not not10813(N33786,in0);
not not10814(N33787,R2);
not not10815(N33798,in0);
not not10816(N33799,R0);
not not10817(N33800,R3);
not not10818(N33810,in0);
not not10819(N33811,R0);
not not10820(N33812,R2);
not not10821(N33822,in0);
not not10822(N33834,in0);
not not10823(N33846,R1);
not not10824(N33858,in2);
not not10825(N33859,R1);
not not10826(N33870,in0);
not not10827(N33871,R2);
not not10828(N33882,in0);
not not10829(N33883,R0);
not not10830(N33894,in0);
not not10831(N33906,in0);
not not10832(N33907,R1);
not not10833(N33908,R2);
not not10834(N33918,in0);
not not10835(N33919,in2);
not not10836(N33930,in0);
not not10837(N33931,in1);
not not10838(N33942,in0);
not not10839(N33943,in2);
not not10840(N33954,in0);
not not10841(N33955,in1);
not not10842(N33956,in2);
not not10843(N33966,in0);
not not10844(N33967,in2);
not not10845(N33968,R1);
not not10846(N33978,R1);
not not10847(N33979,R3);
not not10848(N33989,R1);
not not10849(N34000,in0);
not not10850(N34011,in0);
not not10851(N34022,R3);
not not10852(N34033,R3);
not not10853(N34044,in0);
not not10854(N34053,in0);
not not10855(N34054,in1);
not not10856(N34055,R1);
not not10857(N34056,R2);
not not10858(N34057,R3);
not not10859(N34058,R5);
not not10860(N34069,in0);
not not10861(N34070,in1);
not not10862(N34071,in2);
not not10863(N34072,R2);
not not10864(N34073,R3);
not not10865(N34084,in0);
not not10866(N34085,in2);
not not10867(N34086,R1);
not not10868(N34087,R2);
not not10869(N34088,R3);
not not10870(N34089,R4);
not not10871(N34099,in0);
not not10872(N34100,in1);
not not10873(N34101,in2);
not not10874(N34102,R1);
not not10875(N34103,R3);
not not10876(N34104,R4);
not not10877(N34114,R0);
not not10878(N34115,R2);
not not10879(N34116,R3);
not not10880(N34117,R4);
not not10881(N34118,R5);
not not10882(N34128,in0);
not not10883(N34129,R1);
not not10884(N34130,R3);
not not10885(N34131,R5);
not not10886(N34142,in0);
not not10887(N34143,R0);
not not10888(N34144,R3);
not not10889(N34145,R4);
not not10890(N34156,in0);
not not10891(N34157,in1);
not not10892(N34158,R0);
not not10893(N34159,R1);
not not10894(N34170,in0);
not not10895(N34171,in1);
not not10896(N34172,R1);
not not10897(N34173,R4);
not not10898(N34184,in0);
not not10899(N34185,in2);
not not10900(N34186,R0);
not not10901(N34187,R3);
not not10902(N34188,R4);
not not10903(N34189,R5);
not not10904(N34198,in0);
not not10905(N34199,in1);
not not10906(N34200,R0);
not not10907(N34201,R2);
not not10908(N34212,R0);
not not10909(N34213,R1);
not not10910(N34214,R2);
not not10911(N34215,R3);
not not10912(N34226,in0);
not not10913(N34227,in1);
not not10914(N34228,in2);
not not10915(N34229,R1);
not not10916(N34230,R3);
not not10917(N34240,R0);
not not10918(N34241,R2);
not not10919(N34242,R3);
not not10920(N34243,R4);
not not10921(N34254,in0);
not not10922(N34255,in2);
not not10923(N34256,R3);
not not10924(N34257,R4);
not not10925(N34268,in0);
not not10926(N34269,in1);
not not10927(N34270,R0);
not not10928(N34271,R2);
not not10929(N34272,R4);
not not10930(N34282,in0);
not not10931(N34283,R0);
not not10932(N34284,R1);
not not10933(N34285,R4);
not not10934(N34296,in0);
not not10935(N34297,in1);
not not10936(N34298,in2);
not not10937(N34299,R0);
not not10938(N34300,R1);
not not10939(N34310,in0);
not not10940(N34311,in2);
not not10941(N34312,R0);
not not10942(N34313,R1);
not not10943(N34314,R3);
not not10944(N34324,R1);
not not10945(N34325,R2);
not not10946(N34326,R3);
not not10947(N34327,R5);
not not10948(N34337,in0);
not not10949(N34338,in2);
not not10950(N34339,R3);
not not10951(N34350,R0);
not not10952(N34351,R3);
not not10953(N34352,R5);
not not10954(N34363,in0);
not not10955(N34364,in2);
not not10956(N34365,R3);
not not10957(N34376,in0);
not not10958(N34377,in1);
not not10959(N34378,in2);
not not10960(N34379,R4);
not not10961(N34389,in0);
not not10962(N34390,in1);
not not10963(N34391,in2);
not not10964(N34392,R2);
not not10965(N34393,R5);
not not10966(N34402,R0);
not not10967(N34403,R2);
not not10968(N34404,R4);
not not10969(N34405,R5);
not not10970(N34415,in0);
not not10971(N34416,in1);
not not10972(N34417,in2);
not not10973(N34418,R2);
not not10974(N34428,in0);
not not10975(N34429,in1);
not not10976(N34430,R1);
not not10977(N34431,R3);
not not10978(N34441,in0);
not not10979(N34442,R1);
not not10980(N34453,in0);
not not10981(N34454,R1);
not not10982(N34455,R4);
not not10983(N34465,in0);
not not10984(N34466,R3);
not not10985(N34477,in0);
not not10986(N34478,in1);
not not10987(N34479,R1);
not not10988(N34480,R4);
not not10989(N34489,in0);
not not10990(N34490,R3);
not not10991(N34491,R4);
not not10992(N34501,in0);
not not10993(N34502,R0);
not not10994(N34513,in0);
not not10995(N34514,R3);
not not10996(N34515,R4);
not not10997(N34525,in0);
not not10998(N34526,in2);
not not10999(N34527,R0);
not not11000(N34537,in0);
not not11001(N34538,R1);
not not11002(N34539,R3);
not not11003(N34549,in0);
not not11004(N34550,in2);
not not11005(N34551,R1);
not not11006(N34561,in0);
not not11007(N34562,in1);
not not11008(N34563,R2);
not not11009(N34573,R3);
not not11010(N34574,R4);
not not11011(N34585,R0);
not not11012(N34586,R1);
not not11013(N34587,R3);
not not11014(N34597,R0);
not not11015(N34598,R1);
not not11016(N34599,R3);
not not11017(N34600,R5);
not not11018(N34609,R2);
not not11019(N34610,R3);
not not11020(N34621,in0);
not not11021(N34622,R3);
not not11022(N34623,R4);
not not11023(N34633,in0);
not not11024(N34634,R2);
not not11025(N34635,R4);
not not11026(N34645,in0);
not not11027(N34646,R0);
not not11028(N34647,R5);
not not11029(N34657,in0);
not not11030(N34658,in2);
not not11031(N34659,R3);
not not11032(N34669,in0);
not not11033(N34670,in1);
not not11034(N34671,R2);
not not11035(N34672,R5);
not not11036(N34681,in0);
not not11037(N34682,in1);
not not11038(N34683,R5);
not not11039(N34693,in0);
not not11040(N34694,in1);
not not11041(N34695,in2);
not not11042(N34696,R5);
not not11043(N34705,in0);
not not11044(N34706,R0);
not not11045(N34707,R2);
not not11046(N34716,R0);
not not11047(N34717,R2);
not not11048(N34727,in0);
not not11049(N34728,in1);
not not11050(N34729,R3);
not not11051(N34738,in0);
not not11052(N34739,in2);
not not11053(N34740,R0);
not not11054(N34749,in0);
not not11055(N34750,in1);
not not11056(N34751,R4);
not not11057(N34760,R1);
not not11058(N34761,R3);
not not11059(N34770,R3);
not not11060(N34771,R5);
not not11061(N34780,R3);
not not11062(N34790,R2);
not not11063(N34798,R1);
not not11064(N34799,R2);
not not11065(N34800,R4);
not not11066(N34801,R5);
not not11067(N34809,R1);
not not11068(N34810,R2);
not not11069(N34811,R4);
not not11070(N34812,R5);
not not11071(N34820,R0);
not not11072(N34821,R1);
not not11073(N34822,R2);
not not11074(N34823,R7);
not not11075(N31796,R2);
not not11076(N31797,R6);
not not11077(N31798,R7);
not not11078(N31813,R4);
not not11079(N31814,R5);
not not11080(N31815,R6);
not not11081(N31816,R7);
not not11082(N31832,R4);
not not11083(N31833,R5);
not not11084(N31834,R7);
not not11085(N31849,R3);
not not11086(N31850,R5);
not not11087(N31851,R6);
not not11088(N31852,R7);
not not11089(N31867,R3);
not not11090(N31868,R4);
not not11091(N31869,R6);
not not11092(N31870,R7);
not not11093(N31886,R4);
not not11094(N31887,R6);
not not11095(N31888,R7);
not not11096(N31903,R4);
not not11097(N31904,R5);
not not11098(N31905,R6);
not not11099(N31906,R7);
not not11100(N31922,R4);
not not11101(N31923,R5);
not not11102(N31924,R6);
not not11103(N31938,R4);
not not11104(N31939,R5);
not not11105(N31940,R6);
not not11106(N31941,R7);
not not11107(N31956,R4);
not not11108(N31957,R5);
not not11109(N31958,R6);
not not11110(N31974,R4);
not not11111(N31975,R6);
not not11112(N31990,R4);
not not11113(N31991,R5);
not not11114(N31992,R7);
not not11115(N32008,R5);
not not11116(N32009,R6);
not not11117(N32025,R6);
not not11118(N32026,R7);
not not11119(N32039,R4);
not not11120(N32040,R5);
not not11121(N32041,R6);
not not11122(N32042,R7);
not not11123(N32056,R4);
not not11124(N32057,R5);
not not11125(N32058,R7);
not not11126(N32072,R4);
not not11127(N32073,R5);
not not11128(N32074,R7);
not not11129(N32088,R3);
not not11130(N32089,R4);
not not11131(N32090,R6);
not not11132(N32104,R3);
not not11133(N32105,R4);
not not11134(N32106,R7);
not not11135(N32120,R4);
not not11136(N32121,R6);
not not11137(N32122,R7);
not not11138(N32136,R4);
not not11139(N32137,R5);
not not11140(N32138,R7);
not not11141(N32152,R3);
not not11142(N32153,R6);
not not11143(N32154,R7);
not not11144(N32169,R4);
not not11145(N32170,R7);
not not11146(N32184,R4);
not not11147(N32185,R5);
not not11148(N32186,R6);
not not11149(N32200,R4);
not not11150(N32201,R6);
not not11151(N32202,R7);
not not11152(N32216,R3);
not not11153(N32217,R4);
not not11154(N32218,R6);
not not11155(N32231,R4);
not not11156(N32232,R5);
not not11157(N32233,R6);
not not11158(N32234,R7);
not not11159(N32248,R3);
not not11160(N32249,R4);
not not11161(N32250,R6);
not not11162(N32264,R3);
not not11163(N32265,R4);
not not11164(N32266,R6);
not not11165(N32280,R4);
not not11166(N32281,R5);
not not11167(N32282,R6);
not not11168(N32297,R3);
not not11169(N32298,R6);
not not11170(N32313,R4);
not not11171(N32314,R6);
not not11172(N32328,R3);
not not11173(N32329,R5);
not not11174(N32330,R7);
not not11175(N32345,R5);
not not11176(N32346,R6);
not not11177(N32360,R4);
not not11178(N32361,R5);
not not11179(N32362,R7);
not not11180(N32376,R4);
not not11181(N32377,R5);
not not11182(N32378,R7);
not not11183(N32392,R4);
not not11184(N32393,R5);
not not11185(N32394,R7);
not not11186(N32408,R4);
not not11187(N32409,R5);
not not11188(N32410,R6);
not not11189(N32425,R4);
not not11190(N32426,R6);
not not11191(N32441,R6);
not not11192(N32453,R3);
not not11193(N32454,R4);
not not11194(N32455,R5);
not not11195(N32456,R7);
not not11196(N32468,R4);
not not11197(N32469,R5);
not not11198(N32470,R6);
not not11199(N32471,R7);
not not11200(N32483,R4);
not not11201(N32484,R5);
not not11202(N32485,R6);
not not11203(N32486,R7);
not not11204(N32499,R5);
not not11205(N32500,R6);
not not11206(N32501,R7);
not not11207(N32514,R5);
not not11208(N32515,R6);
not not11209(N32516,R7);
not not11210(N32530,R5);
not not11211(N32531,R6);
not not11212(N32545,R6);
not not11213(N32546,R7);
not not11214(N32559,R4);
not not11215(N32560,R5);
not not11216(N32561,R6);
not not11217(N32574,R5);
not not11218(N32575,R6);
not not11219(N32576,R7);
not not11220(N32590,R3);
not not11221(N32591,R6);
not not11222(N32604,R4);
not not11223(N32605,R6);
not not11224(N32606,R7);
not not11225(N32620,R4);
not not11226(N32621,R5);
not not11227(N32635,R5);
not not11228(N32636,R7);
not not11229(N32650,R5);
not not11230(N32651,R7);
not not11231(N32679,R3);
not not11232(N32680,R4);
not not11233(N32681,R5);
not not11234(N32695,R5);
not not11235(N32696,R7);
not not11236(N32709,R4);
not not11237(N32710,R5);
not not11238(N32711,R7);
not not11239(N32723,R4);
not not11240(N32724,R5);
not not11241(N32725,R6);
not not11242(N32726,R7);
not not11243(N32741,R5);
not not11244(N32755,R5);
not not11245(N32756,R6);
not not11246(N32769,R4);
not not11247(N32770,R5);
not not11248(N32771,R6);
not not11249(N32785,R5);
not not11250(N32786,R6);
not not11251(N32800,R4);
not not11252(N32801,R7);
not not11253(N32813,R4);
not not11254(N32814,R5);
not not11255(N32815,R6);
not not11256(N32816,R7);
not not11257(N32830,R6);
not not11258(N32843,R4);
not not11259(N32844,R6);
not not11260(N32857,R3);
not not11261(N32858,R5);
not not11262(N32872,R6);
not not11263(N32884,R4);
not not11264(N32885,R5);
not not11265(N32886,R7);
not not11266(N32899,R6);
not not11267(N32900,R7);
not not11268(N32913,R5);
not not11269(N32914,R6);
not not11270(N32941,R4);
not not11271(N32942,R6);
not not11272(N32955,R4);
not not11273(N32956,R7);
not not11274(N32969,R5);
not not11275(N32970,R7);
not not11276(N32983,R4);
not not11277(N32984,R7);
not not11278(N32996,R4);
not not11279(N32997,R5);
not not11280(N32998,R6);
not not11281(N33024,R4);
not not11282(N33025,R5);
not not11283(N33026,R6);
not not11284(N33040,R5);
not not11285(N33054,R5);
not not11286(N33067,R4);
not not11287(N33068,R5);
not not11288(N33082,R4);
not not11289(N33095,R4);
not not11290(N33096,R7);
not not11291(N33109,R4);
not not11292(N33110,R5);
not not11293(N33123,R3);
not not11294(N33124,R4);
not not11295(N33137,R3);
not not11296(N33138,R6);
not not11297(N33152,R7);
not not11298(N33179,R5);
not not11299(N33180,R7);
not not11300(N33193,R6);
not not11301(N33194,R7);
not not11302(N33207,R3);
not not11303(N33208,R4);
not not11304(N33221,R4);
not not11305(N33222,R5);
not not11306(N33235,R5);
not not11307(N33236,R7);
not not11308(N33250,R5);
not not11309(N33263,R6);
not not11310(N33264,R7);
not not11311(N33278,R6);
not not11312(N33292,R3);
not not11313(N33306,R6);
not not11314(N33320,R6);
not not11315(N33334,R4);
not not11316(N33348,R7);
not not11317(N33362,R4);
not not11318(N33375,R3);
not not11319(N33376,R4);
not not11320(N33389,R6);
not not11321(N33390,R7);
not not11322(N33403,R5);
not not11323(N33404,R6);
not not11324(N33417,R7);
not not11325(N33430,R5);
not not11326(N33443,R5);
not not11327(N33456,R3);
not not11328(N33468,R5);
not not11329(N33469,R7);
not not11330(N33482,R4);
not not11331(N33494,R3);
not not11332(N33495,R5);
not not11333(N33507,R5);
not not11334(N33508,R7);
not not11335(N33521,R7);
not not11336(N33533,R4);
not not11337(N33534,R7);
not not11338(N33546,R6);
not not11339(N33547,R7);
not not11340(N33560,R6);
not not11341(N33572,R5);
not not11342(N33573,R7);
not not11343(N33610,R4);
not not11344(N33611,R6);
not not11345(N33612,R7);
not not11346(N33624,R4);
not not11347(N33625,R6);
not not11348(N33638,R4);
not not11349(N33651,R6);
not not11350(N33664,R6);
not not11351(N33677,R7);
not not11352(N33689,R4);
not not11353(N33690,R7);
not not11354(N33716,R7);
not not11355(N33728,R4);
not not11356(N33740,R5);
not not11357(N33752,R6);
not not11358(N33764,R4);
not not11359(N33775,R5);
not not11360(N33776,R6);
not not11361(N33788,R4);
not not11362(N33823,R5);
not not11363(N33824,R7);
not not11364(N33835,R4);
not not11365(N33836,R5);
not not11366(N33847,R5);
not not11367(N33848,R7);
not not11368(N33860,R7);
not not11369(N33872,R4);
not not11370(N33884,R4);
not not11371(N33895,R6);
not not11372(N33896,R7);
not not11373(N33920,R7);
not not11374(N33932,R6);
not not11375(N33944,R5);
not not11376(N33990,R7);
not not11377(N34001,R3);
not not11378(N34012,R4);
not not11379(N34023,R4);
not not11380(N34034,R4);
not not11381(N34059,R6);
not not11382(N34060,R7);
not not11383(N34074,R6);
not not11384(N34075,R7);
not not11385(N34090,R6);
not not11386(N34105,R6);
not not11387(N34119,R6);
not not11388(N34132,R6);
not not11389(N34133,R7);
not not11390(N34146,R5);
not not11391(N34147,R6);
not not11392(N34160,R6);
not not11393(N34161,R7);
not not11394(N34174,R5);
not not11395(N34175,R6);
not not11396(N34202,R5);
not not11397(N34203,R6);
not not11398(N34216,R6);
not not11399(N34217,R7);
not not11400(N34231,R5);
not not11401(N34244,R6);
not not11402(N34245,R7);
not not11403(N34258,R6);
not not11404(N34259,R7);
not not11405(N34273,R6);
not not11406(N34286,R6);
not not11407(N34287,R7);
not not11408(N34301,R6);
not not11409(N34315,R6);
not not11410(N34328,R7);
not not11411(N34340,R6);
not not11412(N34341,R7);
not not11413(N34353,R6);
not not11414(N34354,R7);
not not11415(N34366,R6);
not not11416(N34367,R7);
not not11417(N34380,R7);
not not11418(N34406,R7);
not not11419(N34419,R6);
not not11420(N34432,R5);
not not11421(N34443,R6);
not not11422(N34444,R7);
not not11423(N34456,R6);
not not11424(N34467,R6);
not not11425(N34468,R7);
not not11426(N34492,R6);
not not11427(N34503,R5);
not not11428(N34504,R6);
not not11429(N34516,R7);
not not11430(N34528,R7);
not not11431(N34540,R7);
not not11432(N34552,R6);
not not11433(N34564,R6);
not not11434(N34575,R6);
not not11435(N34576,R7);
not not11436(N34588,R7);
not not11437(N34611,R6);
not not11438(N34612,R7);
not not11439(N34624,R7);
not not11440(N34636,R7);
not not11441(N34648,R6);
not not11442(N34660,R7);
not not11443(N34684,R6);
not not11444(N34718,R6);
not not11445(N34781,R6);
not not11446(N34895,R0);
not not11447(N34919,R0);
not not11448(N34931,R0);
not not11449(N34943,R1);
not not11450(N34954,R0);
not not11451(N34965,R0);
not not11452(N34976,R0);
not not11453(N34987,R0);
not not11454(N34998,R0);
not not11455(N35008,R0);
not not11456(N35018,R0);
not not11457(N35038,R0);
not not11458(N35058,R0);
not not11459(N35088,R0);
not not11460(N35137,R0);
not not11461(N35146,R0);
not not11462(N35155,R0);
not not11463(N35164,R0);
not not11464(N35182,R0);
not not11465(N35191,R0);
not not11466(N35209,R0);
not not11467(N35252,R0);
not not11468(N35268,R1);
not not11469(N35291,R0);
not not11470(N35319,R0);
not not11471(N35326,R0);
not not11472(N35332,R0);
not not11473(N35333,R1);
not not11474(N35342,R1);
not not11475(N35350,R1);
not not11476(N35358,R0);
not not11477(N34884,R1);
not not11478(N34885,R2);
not not11479(N34886,R4);
not not11480(N34887,R6);
not not11481(N34888,R7);
not not11482(N34896,R2);
not not11483(N34897,R4);
not not11484(N34898,R5);
not not11485(N34899,R6);
not not11486(N34900,R7);
not not11487(N34907,R1);
not not11488(N34908,R3);
not not11489(N34909,R4);
not not11490(N34910,R5);
not not11491(N34911,R6);
not not11492(N34912,R7);
not not11493(N34920,R1);
not not11494(N34921,R3);
not not11495(N34922,R4);
not not11496(N34923,R5);
not not11497(N34924,R7);
not not11498(N34932,R2);
not not11499(N34933,R3);
not not11500(N34934,R4);
not not11501(N34935,R5);
not not11502(N34936,R6);
not not11503(N34944,R4);
not not11504(N34945,R5);
not not11505(N34946,R6);
not not11506(N34947,R7);
not not11507(N34955,R1);
not not11508(N34956,R3);
not not11509(N34957,R4);
not not11510(N34958,R7);
not not11511(N34966,R1);
not not11512(N34967,R2);
not not11513(N34968,R3);
not not11514(N34969,R6);
not not11515(N34977,R2);
not not11516(N34978,R3);
not not11517(N34979,R4);
not not11518(N34980,R6);
not not11519(N34988,R2);
not not11520(N34989,R4);
not not11521(N34990,R5);
not not11522(N34991,R7);
not not11523(N34999,R3);
not not11524(N35000,R4);
not not11525(N35001,R5);
not not11526(N35009,R1);
not not11527(N35010,R4);
not not11528(N35011,R6);
not not11529(N35019,R1);
not not11530(N35020,R5);
not not11531(N35021,R6);
not not11532(N35028,R1);
not not11533(N35029,R2);
not not11534(N35030,R3);
not not11535(N35031,R6);
not not11536(N35039,R2);
not not11537(N35040,R6);
not not11538(N35041,R7);
not not11539(N35048,R1);
not not11540(N35049,R2);
not not11541(N35050,R4);
not not11542(N35051,R5);
not not11543(N35059,R1);
not not11544(N35060,R6);
not not11545(N35061,R7);
not not11546(N35068,R1);
not not11547(N35069,R2);
not not11548(N35070,R5);
not not11549(N35071,R7);
not not11550(N35078,R1);
not not11551(N35079,R2);
not not11552(N35080,R3);
not not11553(N35081,R4);
not not11554(N35089,R1);
not not11555(N35090,R2);
not not11556(N35091,R7);
not not11557(N35098,R1);
not not11558(N35099,R3);
not not11559(N35100,R6);
not not11560(N35101,R7);
not not11561(N35108,R3);
not not11562(N35109,R4);
not not11563(N35110,R6);
not not11564(N35111,R7);
not not11565(N35118,R2);
not not11566(N35119,R3);
not not11567(N35120,R5);
not not11568(N35121,R6);
not not11569(N35128,R1);
not not11570(N35129,R4);
not not11571(N35130,R6);
not not11572(N35138,R1);
not not11573(N35139,R6);
not not11574(N35147,R2);
not not11575(N35148,R6);
not not11576(N35156,R1);
not not11577(N35157,R2);
not not11578(N35165,R3);
not not11579(N35166,R6);
not not11580(N35173,R1);
not not11581(N35174,R4);
not not11582(N35175,R5);
not not11583(N35183,R1);
not not11584(N35184,R3);
not not11585(N35192,R4);
not not11586(N35193,R7);
not not11587(N35200,R4);
not not11588(N35201,R6);
not not11589(N35202,R7);
not not11590(N35210,R1);
not not11591(N35211,R3);
not not11592(N35218,R2);
not not11593(N35219,R6);
not not11594(N35220,R7);
not not11595(N35227,R4);
not not11596(N35228,R5);
not not11597(N35229,R6);
not not11598(N35236,R3);
not not11599(N35237,R4);
not not11600(N35244,R1);
not not11601(N35245,R6);
not not11602(N35253,R7);
not not11603(N35260,R3);
not not11604(N35261,R5);
not not11605(N35269,R3);
not not11606(N35276,R3);
not not11607(N35277,R6);
not not11608(N35284,R7);
not not11609(N35298,R7);
not not11610(N35305,R5);
not not11611(N35312,R2);
not not11612(N35334,R2);
not not11613(N35335,R6);
not not11614(N35336,R7);
not not11615(N35343,R2);
not not11616(N35344,R3);
not not11617(N35351,R5);
not not11618(N35352,R7);
not not11619(N35359,R3);
not not11620(N35360,R6);
not not11621(N35366,R3);
not not11622(N35367,R6);
not not11623(N35368,R7);
not not11624(N35374,R2);
not not11625(N35471,R0);
not not11626(N35483,R0);
not not11627(N35495,R0);
not not11628(N35516,R0);
not not11629(N35526,R0);
not not11630(N35546,R0);
not not11631(N35556,R1);
not not11632(N35624,R0);
not not11633(N35633,R0);
not not11634(N35642,R0);
not not11635(N35651,R0);
not not11636(N35736,R0);
not not11637(N35418,R3);
not not11638(N35419,R4);
not not11639(N35420,R5);
not not11640(N35421,R6);
not not11641(N35422,R7);
not not11642(N35430,R0);
not not11643(N35431,R1);
not not11644(N35432,R3);
not not11645(N35433,R6);
not not11646(N35434,R7);
not not11647(N35442,R0);
not not11648(N35443,R1);
not not11649(N35444,R2);
not not11650(N35445,R6);
not not11651(N35453,R3);
not not11652(N35454,R4);
not not11653(N35455,R6);
not not11654(N35463,R4);
not not11655(N35464,R5);
not not11656(N35472,R1);
not not11657(N35473,R3);
not not11658(N35474,R4);
not not11659(N35475,R5);
not not11660(N35476,R6);
not not11661(N35484,R1);
not not11662(N35485,R2);
not not11663(N35486,R4);
not not11664(N35487,R5);
not not11665(N35488,R6);
not not11666(N35496,R1);
not not11667(N35497,R3);
not not11668(N35498,R4);
not not11669(N35499,R6);
not not11670(N35506,R1);
not not11671(N35507,R2);
not not11672(N35508,R4);
not not11673(N35509,R6);
not not11674(N35517,R5);
not not11675(N35518,R6);
not not11676(N35519,R7);
not not11677(N35527,R4);
not not11678(N35528,R5);
not not11679(N35529,R7);
not not11680(N35536,R2);
not not11681(N35537,R4);
not not11682(N35538,R6);
not not11683(N35539,R7);
not not11684(N35547,R3);
not not11685(N35548,R4);
not not11686(N35549,R7);
not not11687(N35557,R2);
not not11688(N35558,R4);
not not11689(N35559,R7);
not not11690(N35566,R2);
not not11691(N35567,R5);
not not11692(N35568,R6);
not not11693(N35569,R7);
not not11694(N35576,R2);
not not11695(N35577,R4);
not not11696(N35578,R5);
not not11697(N35579,R6);
not not11698(N35586,R1);
not not11699(N35587,R4);
not not11700(N35588,R6);
not not11701(N35589,R7);
not not11702(N35596,R1);
not not11703(N35597,R3);
not not11704(N35598,R5);
not not11705(N35599,R6);
not not11706(N35606,R2);
not not11707(N35607,R5);
not not11708(N35608,R7);
not not11709(N35615,R1);
not not11710(N35616,R3);
not not11711(N35617,R7);
not not11712(N35625,R1);
not not11713(N35626,R5);
not not11714(N35634,R1);
not not11715(N35635,R4);
not not11716(N35643,R1);
not not11717(N35644,R4);
not not11718(N35652,R5);
not not11719(N35653,R6);
not not11720(N35660,R1);
not not11721(N35661,R2);
not not11722(N35662,R4);
not not11723(N35669,R5);
not not11724(N35670,R6);
not not11725(N35671,R7);
not not11726(N35678,R1);
not not11727(N35679,R3);
not not11728(N35680,R6);
not not11729(N35687,R3);
not not11730(N35688,R5);
not not11731(N35689,R6);
not not11732(N35696,R2);
not not11733(N35697,R6);
not not11734(N35704,R2);
not not11735(N35705,R6);
not not11736(N35712,R4);
not not11737(N35713,R7);
not not11738(N35720,R1);
not not11739(N35721,R5);
not not11740(N35728,R2);
not not11741(N35729,R6);
not not11742(N35737,R4);
not not11743(N35744,R3);
not not11744(N35751,R6);
not not11745(N35758,R1);
not not11746(N35911,R0);
not not11747(N35920,R0);
not not11748(N35779,R1);
not not11749(N35780,R2);
not not11750(N35781,R4);
not not11751(N35782,R5);
not not11752(N35783,R6);
not not11753(N35784,R7);
not not11754(N35792,R1);
not not11755(N35793,R2);
not not11756(N35794,R3);
not not11757(N35795,R4);
not not11758(N35796,R5);
not not11759(N35797,R7);
not not11760(N35805,R1);
not not11761(N35806,R3);
not not11762(N35807,R4);
not not11763(N35808,R5);
not not11764(N35809,R6);
not not11765(N35817,R0);
not not11766(N35818,R1);
not not11767(N35819,R4);
not not11768(N35820,R6);
not not11769(N35821,R7);
not not11770(N35829,R0);
not not11771(N35830,R1);
not not11772(N35831,R2);
not not11773(N35832,R4);
not not11774(N35833,R6);
not not11775(N35841,R0);
not not11776(N35842,R1);
not not11777(N35843,R3);
not not11778(N35844,R4);
not not11779(N35845,R5);
not not11780(N35853,R1);
not not11781(N35854,R2);
not not11782(N35855,R6);
not not11783(N35856,R7);
not not11784(N35864,R1);
not not11785(N35865,R2);
not not11786(N35866,R5);
not not11787(N35867,R6);
not not11788(N35875,R3);
not not11789(N35876,R5);
not not11790(N35877,R7);
not not11791(N35885,R1);
not not11792(N35886,R4);
not not11793(N35894,R5);
not not11794(N35895,R6);
not not11795(N35903,R2);
not not11796(N35904,R7);
not not11797(N35912,R2);
not not11798(N35913,R4);
not not11799(N35921,R3);
not not11800(N36039,R0);
not not11801(N36051,R1);
not not11802(N36063,R0);
not not11803(N36074,R0);
not not11804(N36095,R0);
not not11805(N36105,R0);
not not11806(N36115,R0);
not not11807(N36125,R1);
not not11808(N36165,R1);
not not11809(N36175,R0);
not not11810(N36205,R0);
not not11811(N36233,R0);
not not11812(N36242,R0);
not not11813(N36292,R0);
not not11814(N36300,R0);
not not11815(N36384,R2);
not not11816(N35973,R1);
not not11817(N35974,R2);
not not11818(N35975,R3);
not not11819(N35976,R4);
not not11820(N35977,R5);
not not11821(N35978,R7);
not not11822(N35986,R3);
not not11823(N35987,R4);
not not11824(N35988,R5);
not not11825(N35989,R6);
not not11826(N35990,R7);
not not11827(N35998,R0);
not not11828(N35999,R1);
not not11829(N36000,R3);
not not11830(N36001,R6);
not not11831(N36002,R7);
not not11832(N36010,R1);
not not11833(N36011,R2);
not not11834(N36012,R6);
not not11835(N36013,R7);
not not11836(N36021,R3);
not not11837(N36022,R4);
not not11838(N36023,R6);
not not11839(N36031,R4);
not not11840(N36032,R5);
not not11841(N36040,R1);
not not11842(N36041,R3);
not not11843(N36042,R4);
not not11844(N36043,R5);
not not11845(N36044,R6);
not not11846(N36052,R2);
not not11847(N36053,R4);
not not11848(N36054,R5);
not not11849(N36055,R6);
not not11850(N36056,R7);
not not11851(N36064,R1);
not not11852(N36065,R2);
not not11853(N36066,R4);
not not11854(N36067,R6);
not not11855(N36075,R1);
not not11856(N36076,R3);
not not11857(N36077,R4);
not not11858(N36078,R6);
not not11859(N36085,R1);
not not11860(N36086,R2);
not not11861(N36087,R4);
not not11862(N36088,R6);
not not11863(N36096,R5);
not not11864(N36097,R6);
not not11865(N36098,R7);
not not11866(N36106,R4);
not not11867(N36107,R5);
not not11868(N36108,R7);
not not11869(N36116,R3);
not not11870(N36117,R4);
not not11871(N36118,R7);
not not11872(N36126,R2);
not not11873(N36127,R4);
not not11874(N36128,R7);
not not11875(N36135,R2);
not not11876(N36136,R5);
not not11877(N36137,R6);
not not11878(N36138,R7);
not not11879(N36145,R2);
not not11880(N36146,R4);
not not11881(N36147,R5);
not not11882(N36148,R6);
not not11883(N36155,R1);
not not11884(N36156,R3);
not not11885(N36157,R5);
not not11886(N36158,R6);
not not11887(N36166,R4);
not not11888(N36167,R6);
not not11889(N36168,R7);
not not11890(N36176,R1);
not not11891(N36177,R4);
not not11892(N36178,R5);
not not11893(N36185,R1);
not not11894(N36186,R3);
not not11895(N36187,R4);
not not11896(N36188,R7);
not not11897(N36195,R1);
not not11898(N36196,R3);
not not11899(N36197,R5);
not not11900(N36198,R6);
not not11901(N36206,R1);
not not11902(N36207,R2);
not not11903(N36208,R6);
not not11904(N36215,R2);
not not11905(N36216,R5);
not not11906(N36217,R7);
not not11907(N36224,R2);
not not11908(N36225,R5);
not not11909(N36226,R6);
not not11910(N36234,R1);
not not11911(N36235,R5);
not not11912(N36243,R1);
not not11913(N36244,R4);
not not11914(N36251,R1);
not not11915(N36252,R3);
not not11916(N36253,R6);
not not11917(N36260,R5);
not not11918(N36261,R6);
not not11919(N36268,R2);
not not11920(N36269,R6);
not not11921(N36276,R1);
not not11922(N36277,R5);
not not11923(N36284,R1);
not not11924(N36285,R4);
not not11925(N36293,R3);
not not11926(N36301,R4);
not not11927(N36308,R3);
not not11928(N36309,R7);
not not11929(N36316,R5);
not not11930(N36317,R6);
not not11931(N36324,R5);
not not11932(N36325,R6);
not not11933(N36332,R3);
not not11934(N36333,R7);
not not11935(N36340,R2);
not not11936(N36341,R6);
not not11937(N36348,R2);
not not11938(N36349,R7);
not not11939(N36356,R4);
not not11940(N36357,R7);
not not11941(N36364,R3);
not not11942(N36371,R6);
not not11943(N36378,R1);
not not11944(N36385,R4);
not not11945(N36386,R7);
not not11946(N36575,R0);
not not11947(N36586,R1);
not not11948(N36607,R0);
not not11949(N36617,R0);
not not11950(N36415,R0);
not not11951(N36416,R1);
not not11952(N36417,R2);
not not11953(N36418,R3);
not not11954(N36419,R4);
not not11955(N36420,R5);
not not11956(N36421,R7);
not not11957(N36429,R0);
not not11958(N36430,R2);
not not11959(N36431,R3);
not not11960(N36432,R4);
not not11961(N36433,R5);
not not11962(N36434,R6);
not not11963(N36442,R0);
not not11964(N36443,R1);
not not11965(N36444,R2);
not not11966(N36445,R3);
not not11967(N36446,R6);
not not11968(N36447,R7);
not not11969(N36455,R0);
not not11970(N36456,R2);
not not11971(N36457,R3);
not not11972(N36458,R4);
not not11973(N36459,R6);
not not11974(N36460,R7);
not not11975(N36468,R1);
not not11976(N36469,R2);
not not11977(N36470,R4);
not not11978(N36471,R5);
not not11979(N36472,R6);
not not11980(N36480,R0);
not not11981(N36481,R2);
not not11982(N36482,R4);
not not11983(N36483,R5);
not not11984(N36484,R7);
not not11985(N36492,R2);
not not11986(N36493,R3);
not not11987(N36494,R5);
not not11988(N36495,R6);
not not11989(N36503,R3);
not not11990(N36504,R4);
not not11991(N36505,R6);
not not11992(N36506,R7);
not not11993(N36514,R0);
not not11994(N36515,R4);
not not11995(N36516,R6);
not not11996(N36517,R7);
not not11997(N36525,R4);
not not11998(N36526,R5);
not not11999(N36527,R6);
not not12000(N36528,R7);
not not12001(N36536,R0);
not not12002(N36537,R1);
not not12003(N36538,R3);
not not12004(N36539,R5);
not not12005(N36547,R2);
not not12006(N36548,R3);
not not12007(N36549,R6);
not not12008(N36550,R7);
not not12009(N36558,R1);
not not12010(N36559,R4);
not not12011(N36560,R6);
not not12012(N36568,R2);
not not12013(N36576,R1);
not not12014(N36577,R5);
not not12015(N36578,R6);
not not12016(N36579,R7);
not not12017(N36587,R2);
not not12018(N36588,R5);
not not12019(N36589,R6);
not not12020(N36590,R7);
not not12021(N36597,R3);
not not12022(N36598,R5);
not not12023(N36599,R6);
not not12024(N36600,R7);
not not12025(N36608,R1);
not not12026(N36609,R2);
not not12027(N36610,R7);
not not12028(N36618,R2);
not not12029(N36619,R6);
not not12030(N36626,R1);
not not12031(N36627,R2);
not not12032(N36628,R3);
not not12033(N36635,R1);
not not12034(N36636,R5);
not not12035(N36637,R7);
not not12036(N36644,R1);
not not12037(N36645,R7);
not not12038(N36758,R0);
not not12039(N36782,R0);
not not12040(N36794,R0);
not not12041(N36805,R1);
not not12042(N36816,R0);
not not12043(N36827,R0);
not not12044(N36838,R0);
not not12045(N36848,R0);
not not12046(N36858,R1);
not not12047(N36868,R0);
not not12048(N36878,R0);
not not12049(N36888,R0);
not not12050(N36958,R0);
not not12051(N36976,R0);
not not12052(N36985,R0);
not not12053(N36994,R0);
not not12054(N37003,R0);
not not12055(N37021,R0);
not not12056(N37061,R0);
not not12057(N37085,R1);
not not12058(N37093,R1);
not not12059(N37117,R0);
not not12060(N37124,R0);
not not12061(N37131,R0);
not not12062(N36700,R0);
not not12063(N36701,R1);
not not12064(N36702,R2);
not not12065(N36703,R3);
not not12066(N36704,R5);
not not12067(N36705,R6);
not not12068(N36706,R7);
not not12069(N36714,R1);
not not12070(N36715,R2);
not not12071(N36716,R4);
not not12072(N36717,R6);
not not12073(N36718,R7);
not not12074(N36726,R2);
not not12075(N36727,R3);
not not12076(N36728,R4);
not not12077(N36729,R6);
not not12078(N36730,R7);
not not12079(N36738,R1);
not not12080(N36739,R3);
not not12081(N36740,R4);
not not12082(N36741,R6);
not not12083(N36749,R4);
not not12084(N36750,R5);
not not12085(N36751,R6);
not not12086(N36759,R2);
not not12087(N36760,R4);
not not12088(N36761,R5);
not not12089(N36762,R6);
not not12090(N36763,R7);
not not12091(N36770,R1);
not not12092(N36771,R3);
not not12093(N36772,R4);
not not12094(N36773,R5);
not not12095(N36774,R6);
not not12096(N36775,R7);
not not12097(N36783,R1);
not not12098(N36784,R2);
not not12099(N36785,R3);
not not12100(N36786,R4);
not not12101(N36787,R6);
not not12102(N36795,R1);
not not12103(N36796,R3);
not not12104(N36797,R4);
not not12105(N36798,R7);
not not12106(N36806,R4);
not not12107(N36807,R5);
not not12108(N36808,R6);
not not12109(N36809,R7);
not not12110(N36817,R1);
not not12111(N36818,R3);
not not12112(N36819,R4);
not not12113(N36820,R7);
not not12114(N36828,R2);
not not12115(N36829,R5);
not not12116(N36830,R6);
not not12117(N36831,R7);
not not12118(N36839,R3);
not not12119(N36840,R4);
not not12120(N36841,R5);
not not12121(N36849,R1);
not not12122(N36850,R6);
not not12123(N36851,R7);
not not12124(N36859,R2);
not not12125(N36860,R3);
not not12126(N36861,R6);
not not12127(N36869,R1);
not not12128(N36870,R4);
not not12129(N36871,R6);
not not12130(N36879,R1);
not not12131(N36880,R5);
not not12132(N36881,R6);
not not12133(N36889,R2);
not not12134(N36890,R4);
not not12135(N36891,R6);
not not12136(N36898,R1);
not not12137(N36899,R2);
not not12138(N36900,R3);
not not12139(N36901,R6);
not not12140(N36908,R1);
not not12141(N36909,R2);
not not12142(N36910,R3);
not not12143(N36911,R4);
not not12144(N36918,R1);
not not12145(N36919,R2);
not not12146(N36920,R5);
not not12147(N36921,R7);
not not12148(N36928,R1);
not not12149(N36929,R2);
not not12150(N36930,R4);
not not12151(N36931,R5);
not not12152(N36938,R1);
not not12153(N36939,R3);
not not12154(N36940,R6);
not not12155(N36941,R7);
not not12156(N36948,R1);
not not12157(N36949,R3);
not not12158(N36950,R5);
not not12159(N36951,R7);
not not12160(N36959,R1);
not not12161(N36960,R6);
not not12162(N36967,R3);
not not12163(N36968,R6);
not not12164(N36969,R7);
not not12165(N36977,R1);
not not12166(N36978,R2);
not not12167(N36986,R3);
not not12168(N36987,R6);
not not12169(N36995,R3);
not not12170(N36996,R6);
not not12171(N37004,R1);
not not12172(N37005,R3);
not not12173(N37012,R1);
not not12174(N37013,R4);
not not12175(N37014,R5);
not not12176(N37022,R7);
not not12177(N37029,R3);
not not12178(N37030,R4);
not not12179(N37037,R6);
not not12180(N37038,R7);
not not12181(N37045,R1);
not not12182(N37046,R6);
not not12183(N37053,R6);
not not12184(N37054,R7);
not not12185(N37062,R5);
not not12186(N37069,R3);
not not12187(N37070,R5);
not not12188(N37077,R2);
not not12189(N37078,R5);
not not12190(N37086,R3);
not not12191(N37094,R2);
not not12192(N37101,R2);
not not12193(N37102,R4);
not not12194(N37109,R3);
not not12195(N37110,R6);
not not12196(N37138,R7);
not not12197(N37145,R5);

endmodule