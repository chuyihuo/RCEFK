//num of or = 2842
//num of and = 23701
//num of not = 12986
//num of wire = 39527
module c1126 (in0,in1,in2,O0,O1,O2,O3,O4,O5,clk,rst);

input in0,in1,in2,clk,rst;

output O0,O1,O2,O3,O4,O5;

wire in0,in1,in2,N0,N1,N2,N3,N4,N5,N6,N7,N8,
N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,
N19,N20,N21,N22,N23,N24,N25,N26,N27,N28,
N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,
N39,N40,N41,N42,N43,N44,N45,N46,N47,N48,
N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,
N59,N60,N61,N62,N63,N64,N65,N66,N67,N68,
N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,
N79,N80,N81,N82,N83,N84,N85,N86,N87,N88,
N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,
N99,N100,N101,N102,N103,N104,N105,N106,N107,N108,
N109,N110,N111,N112,N113,N114,N115,N116,N117,N118,
N119,N120,N121,N122,N123,N124,N125,N126,N127,N128,
N129,N130,N131,N132,N133,N134,N135,N136,N137,N138,
N139,N140,N141,N142,N143,N144,N145,N146,N147,N148,
N149,N150,N151,N152,N153,N154,N155,N156,N157,N158,
N159,N160,N161,N162,N163,N164,N165,N166,N167,N168,
N169,N170,N171,N172,N173,N174,N175,N176,N177,N178,
N179,N180,N181,N182,N183,N184,N185,N186,N187,N188,
N189,N190,N191,N192,N193,N194,N195,N196,N197,N198,
N199,N200,N201,N202,N203,N204,N205,N206,N207,N208,
N209,N210,N211,N212,N213,N214,N215,N216,N217,N218,
N219,N220,N221,N222,N223,N224,N225,N226,N227,N228,
N229,N230,N231,N232,N233,N234,N235,N236,N237,N238,
N239,N240,N241,N242,N243,N244,N245,N246,N247,N248,
N249,N250,N251,N252,N253,N254,N255,N256,N257,N258,
N259,N260,N261,N262,N263,N264,N265,N266,N267,N268,
N269,N270,N271,N272,N273,N274,N275,N276,N277,N278,
N279,N280,N281,N282,N283,N284,N285,N286,N287,N288,
N289,N290,N291,N292,N293,N294,N295,N296,N297,N298,
N299,N300,N301,N302,N303,N304,N305,N306,N307,N308,
N309,N310,N311,N312,N313,N314,N315,N316,N317,N318,
N319,N320,N321,N322,N323,N324,N325,N326,N327,N328,
N329,N330,N331,N332,N333,N334,N335,N336,N337,N338,
N339,N340,N341,N342,N343,N344,N345,N346,N347,N348,
N349,N350,N351,N352,N353,N354,N355,N356,N357,N358,
N359,N360,N361,N362,N363,N364,N365,N366,N367,N368,
N369,N370,N371,N372,N373,N374,N375,N376,N377,N378,
N379,N380,N381,N382,N383,N384,N385,N386,N387,N388,
N389,N390,N391,N392,N393,N394,N395,N396,N397,N398,
N399,N400,N401,N402,N403,N404,N405,N406,N407,N408,
N409,N410,N411,N412,N413,N414,N415,N416,N417,N418,
N419,N420,N421,N422,N423,N424,N425,N426,N427,N428,
N429,N430,N431,N432,N433,N434,N435,N436,N437,N438,
N439,N440,N441,N442,N443,N444,N445,N446,N447,N448,
N449,N450,N451,N452,N453,N454,N455,N456,N457,N458,
N459,N460,N461,N462,N463,N464,N465,N466,N467,N468,
N469,N470,N471,N472,N473,N474,N475,N476,N477,N478,
N479,N480,N481,N482,N483,N484,N485,N486,N487,N488,
N489,N490,N491,N492,N493,N494,N495,N496,N497,N498,
N499,N500,N501,N502,N503,N504,N505,N506,N507,N508,
N509,N510,N511,N512,N513,N514,N515,N516,N517,N518,
N519,N520,N521,N522,N523,N524,N525,N526,N527,N528,
N529,N530,N531,N532,N533,N534,N535,N536,N537,N538,
N539,N540,N541,N542,N543,N544,N545,N546,N547,N548,
N549,N550,N551,N552,N553,N554,N555,N556,N557,N558,
N559,N560,N561,N562,N563,N564,N565,N566,N567,N568,
N569,N570,N571,N572,N573,N574,N575,N576,N577,N578,
N579,N580,N581,N582,N583,N584,N585,N586,N587,N588,
N589,N590,N591,N592,N593,N594,N595,N596,N597,N598,
N599,N600,N601,N602,N603,N604,N605,N606,N607,N608,
N609,N610,N611,N612,N613,N614,N615,N616,N617,N618,
N619,N620,N621,N622,N623,N624,N625,N626,N627,N628,
N629,N630,N631,N632,N633,N634,N635,N636,N637,N638,
N639,N640,N641,N642,N643,N644,N645,N646,N647,N648,
N649,N650,N651,N652,N653,N654,N655,N656,N657,N658,
N659,N660,N661,N662,N663,N664,N665,N666,N667,N668,
N669,N670,N671,N672,N673,N674,N675,N676,N677,N678,
N679,N680,N681,N682,N683,N684,N685,N686,N687,N688,
N689,N690,N691,N692,N693,N694,N695,N696,N697,N698,
N699,N700,N701,N702,N703,N704,N705,N706,N707,N708,
N709,N710,N711,N712,N713,N714,N715,N716,N717,N718,
N719,N720,N721,N722,N723,N724,N725,N726,N727,N728,
N729,N730,N731,N732,N733,N734,N735,N736,N737,N738,
N739,N740,N741,N742,N743,N744,N745,N746,N747,N748,
N749,N750,N751,N752,N753,N754,N755,N756,N757,N758,
N759,N760,N761,N762,N763,N764,N765,N766,N767,N768,
N769,N770,N771,N772,N773,N774,N775,N776,N777,N778,
N779,N780,N781,N782,N783,N784,N785,N786,N787,N788,
N789,N790,N791,N792,N793,N794,N795,N796,N797,N798,
N799,N800,N801,N802,N803,N804,N805,N806,N807,N808,
N809,N810,N811,N812,N813,N814,N815,N816,N817,N818,
N819,N820,N821,N822,N823,N824,N825,N826,N827,N828,
N829,N830,N831,N832,N833,N834,N835,N836,N837,N838,
N839,N840,N841,N842,N843,N844,N845,N846,N847,N848,
N849,N850,N851,N852,N853,N854,N855,N856,N857,N858,
N859,N860,N861,N862,N863,N864,N865,N866,N867,N868,
N869,N870,N871,N872,N873,N874,N875,N876,N877,N878,
N879,N880,N881,N882,N883,N884,N885,N886,N887,N888,
N889,N890,N891,N892,N893,N894,N895,N896,N897,N898,
N899,N900,N901,N902,N903,N904,N905,N906,N907,N908,
N909,N910,N911,N912,N913,N914,N915,N916,N917,N918,
N919,N920,N921,N922,N923,N924,N925,N926,N927,N928,
N929,N930,N931,N932,N933,N934,N935,N936,N937,N938,
N939,N940,N941,N942,N943,N944,N945,N946,N947,N948,
N949,N950,N951,N952,N953,N954,N955,N956,N957,N958,
N959,N960,N961,N962,N963,N964,N965,N966,N967,N968,
N969,N970,N971,N972,N973,N974,N975,N976,N977,N978,
N979,N980,N981,N982,N983,N984,N985,N986,N987,N988,
N989,N990,N991,N992,N993,N994,N995,N996,N997,N998,
N999,N1000,N1001,N1002,N1003,N1004,N1005,N1006,N1007,N1008,
N1009,N1010,N1011,N1012,N1013,N1014,N1015,N1016,N1017,N1018,
N1019,N1020,N1021,N1022,N1023,N1024,N1025,N1026,N1027,N1028,
N1029,N1030,N1031,N1032,N1033,N1034,N1035,N1036,N1037,N1038,
N1039,N1040,N1041,N1042,N1043,N1044,N1045,N1046,N1047,N1048,
N1049,N1050,N1051,N1052,N1053,N1054,N1055,N1056,N1057,N1058,
N1059,N1060,N1061,N1062,N1063,N1064,N1065,N1066,N1067,N1068,
N1069,N1070,N1071,N1072,N1073,N1074,N1075,N1076,N1077,N1078,
N1079,N1080,N1081,N1082,N1083,N1084,N1085,N1086,N1087,N1088,
N1089,N1090,N1091,N1092,N1093,N1094,N1095,N1096,N1097,N1098,
N1099,N1100,N1101,N1102,N1103,N1104,N1105,N1106,N1107,N1108,
N1109,N1110,N1111,N1112,N1113,N1114,N1115,N1116,N1117,N1118,
N1119,N1120,N1121,N1122,N1123,N1124,N1125,N1126,N1127,N1128,
N1129,N1130,N1131,N1132,N1133,N1134,N1135,N1136,N1137,N1138,
N1139,N1140,N1141,N1142,N1143,N1144,N1145,N1146,N1147,N1148,
N1149,N1150,N1151,N1152,N1153,N1154,N1155,N1156,N1157,N1158,
N1159,N1160,N1161,N1162,N1163,N1164,N1165,N1166,N1167,N1168,
N1169,N1170,N1171,N1172,N1173,N1174,N1175,N1176,N1177,N1178,
N1179,N1180,N1181,N1182,N1183,N1184,N1185,N1186,N1187,N1188,
N1189,N1190,N1191,N1192,N1193,N1194,N1195,N1196,N1197,N1198,
N1199,N1200,N1201,N1202,N1203,N1204,N1205,N1206,N1207,N1208,
N1209,N1210,N1211,N1212,N1213,N1214,N1215,N1216,N1217,N1218,
N1219,N1220,N1221,N1222,N1223,N1224,N1225,N1226,N1227,N1228,
N1229,N1230,N1231,N1232,N1233,N1234,N1235,N1236,N1237,N1238,
N1239,N1240,N1241,N1242,N1243,N1244,N1245,N1246,N1247,N1248,
N1249,N1250,N1251,N1252,N1253,N1254,N1255,N1256,N1257,N1258,
N1259,N1260,N1261,N1262,N1263,N1264,N1265,N1266,N1267,N1268,
N1269,N1270,N1271,N1272,N1273,N1274,N1275,N1276,N1277,N1278,
N1279,N1280,N1281,N1282,N1283,N1284,N1285,N1286,N1287,N1288,
N1289,N1290,N1291,N1292,N1293,N1294,N1295,N1296,N1297,N1298,
N1299,N1300,N1301,N1302,N1303,N1304,N1305,N1306,N1307,N1308,
N1309,N1310,N1311,N1312,N1313,N1314,N1315,N1316,N1317,N1318,
N1319,N1320,N1321,N1322,N1323,N1324,N1325,N1326,N1327,N1328,
N1329,N1330,N1331,N1332,N1333,N1334,N1335,N1336,N1337,N1338,
N1339,N1340,N1341,N1342,N1343,N1344,N1345,N1346,N1347,N1348,
N1349,N1350,N1351,N1352,N1353,N1354,N1355,N1356,N1357,N1358,
N1359,N1360,N1361,N1362,N1363,N1364,N1365,N1366,N1367,N1368,
N1369,N1370,N1371,N1372,N1373,N1374,N1375,N1376,N1377,N1378,
N1379,N1380,N1381,N1382,N1383,N1384,N1385,N1386,N1387,N1388,
N1389,N1390,N1391,N1392,N1393,N1394,N1395,N1396,N1397,N1398,
N1399,N1400,N1401,N1402,N1403,N1404,N1405,N1406,N1407,N1408,
N1409,N1410,N1411,N1412,N1413,N1414,N1415,N1416,N1417,N1418,
N1419,N1420,N1421,N1422,N1423,N1424,N1425,N1426,N1427,N1428,
N1429,N1430,N1431,N1432,N1433,N1434,N1435,N1436,N1437,N1438,
N1439,N1440,N1441,N1442,N1443,N1444,N1445,N1446,N1447,N1448,
N1449,N1450,N1451,N1452,N1453,N1454,N1455,N1456,N1457,N1458,
N1459,N1460,N1461,N1462,N1463,N1464,N1465,N1466,N1467,N1468,
N1469,N1470,N1471,N1472,N1473,N1474,N1475,N1476,N1477,N1478,
N1479,N1480,N1481,N1482,N1483,N1484,N1485,N1486,N1487,N1488,
N1489,N1490,N1491,N1492,N1493,N1494,N1495,N1496,N1497,N1498,
N1499,N1500,N1501,N1502,N1503,N1504,N1505,N1506,N1507,N1508,
N1509,N1510,N1511,N1512,N1513,N1514,N1515,N1516,N1517,N1518,
N1519,N1520,N1521,N1522,N1523,N1524,N1525,N1526,N1527,N1528,
N1529,N1530,N1531,N1532,N1533,N1534,N1535,N1536,N1537,N1538,
N1539,N1540,N1541,N1542,N1543,N1544,N1545,N1546,N1547,N1548,
N1549,N1550,N1551,N1552,N1553,N1554,N1555,N1556,N1557,N1558,
N1559,N1560,N1561,N1562,N1563,N1564,N1565,N1566,N1567,N1568,
N1569,N1570,N1571,N1572,N1573,N1574,N1575,N1576,N1577,N1578,
N1579,N1580,N1581,N1582,N1583,N1584,N1585,N1586,N1587,N1588,
N1589,N1590,N1591,N1592,N1593,N1594,N1595,N1596,N1597,N1598,
N1599,N1600,N1601,N1602,N1603,N1604,N1605,N1606,N1607,N1608,
N1609,N1610,N1611,N1612,N1613,N1614,N1615,N1616,N1617,N1618,
N1619,N1620,N1621,N1622,N1623,N1624,N1625,N1626,N1627,N1628,
N1629,N1630,N1631,N1632,N1633,N1634,N1635,N1636,N1637,N1638,
N1639,N1640,N1641,N1642,N1643,N1644,N1645,N1646,N1647,N1648,
N1649,N1650,N1651,N1652,N1653,N1654,N1655,N1656,N1657,N1658,
N1659,N1660,N1661,N1662,N1663,N1664,N1665,N1666,N1667,N1668,
N1669,N1670,N1671,N1672,N1673,N1674,N1675,N1676,N1677,N1678,
N1679,N1680,N1681,N1682,N1683,N1684,N1685,N1686,N1687,N1688,
N1689,N1690,N1691,N1692,N1693,N1694,N1695,N1696,N1697,N1698,
N1699,N1700,N1701,N1702,N1703,N1704,N1705,N1706,N1707,N1708,
N1709,N1710,N1711,N1712,N1713,N1714,N1715,N1716,N1717,N1718,
N1719,N1720,N1721,N1722,N1723,N1724,N1725,N1726,N1727,N1728,
N1729,N1730,N1731,N1732,N1733,N1734,N1735,N1736,N1737,N1738,
N1739,N1740,N1741,N1742,N1743,N1744,N1745,N1746,N1747,N1748,
N1749,N1750,N1751,N1752,N1753,N1754,N1755,N1756,N1757,N1758,
N1759,N1760,N1761,N1762,N1763,N1764,N1765,N1766,N1767,N1768,
N1769,N1770,N1771,N1772,N1773,N1774,N1775,N1776,N1777,N1778,
N1779,N1780,N1781,N1782,N1783,N1784,N1785,N1786,N1787,N1788,
N1789,N1790,N1791,N1792,N1793,N1794,N1795,N1796,N1797,N1798,
N1799,N1800,N1801,N1802,N1803,N1804,N1805,N1806,N1807,N1808,
N1809,N1810,N1811,N1812,N1813,N1814,N1815,N1816,N1817,N1818,
N1819,N1820,N1821,N1822,N1823,N1824,N1825,N1826,N1827,N1828,
N1829,N1830,N1831,N1832,N1833,N1834,N1835,N1836,N1837,N1838,
N1839,N1840,N1841,N1842,N1843,N1844,N1845,N1846,N1847,N1848,
N1849,N1850,N1851,N1852,N1853,N1854,N1855,N1856,N1857,N1858,
N1859,N1860,N1861,N1862,N1863,N1864,N1865,N1866,N1867,N1868,
N1869,N1870,N1871,N1872,N1873,N1874,N1875,N1876,N1877,N1878,
N1879,N1880,N1881,N1882,N1883,N1884,N1885,N1886,N1887,N1888,
N1889,N1890,N1891,N1892,N1893,N1894,N1895,N1896,N1897,N1898,
N1899,N1900,N1901,N1902,N1903,N1904,N1905,N1906,N1907,N1908,
N1909,N1910,N1911,N1912,N1913,N1914,N1915,N1916,N1917,N1918,
N1919,N1920,N1921,N1922,N1923,N1924,N1925,N1926,N1927,N1928,
N1929,N1930,N1931,N1932,N1933,N1934,N1935,N1936,N1937,N1938,
N1939,N1940,N1941,N1942,N1943,N1944,N1945,N1946,N1947,N1948,
N1949,N1950,N1951,N1952,N1953,N1954,N1955,N1956,N1957,N1958,
N1959,N1960,N1961,N1962,N1963,N1964,N1965,N1966,N1967,N1968,
N1969,N1970,N1971,N1972,N1973,N1974,N1975,N1976,N1977,N1978,
N1979,N1980,N1981,N1982,N1983,N1984,N1985,N1986,N1987,N1988,
N1989,N1990,N1991,N1992,N1993,N1994,N1995,N1996,N1997,N1998,
N1999,N2000,N2001,N2002,N2003,N2004,N2005,N2006,N2007,N2008,
N2009,N2010,N2011,N2012,N2013,N2014,N2015,N2016,N2017,N2018,
N2019,N2020,N2021,N2022,N2023,N2024,N2025,N2026,N2027,N2028,
N2029,N2030,N2031,N2032,N2033,N2034,N2035,N2036,N2037,N2038,
N2039,N2040,N2041,N2042,N2043,N2044,N2045,N2046,N2047,N2048,
N2049,N2050,N2051,N2052,N2053,N2054,N2055,N2056,N2057,N2058,
N2059,N2060,N2061,N2062,N2063,N2064,N2065,N2066,N2067,N2068,
N2069,N2070,N2071,N2072,N2073,N2074,N2075,N2076,N2077,N2078,
N2079,N2080,N2081,N2082,N2083,N2084,N2085,N2086,N2087,N2088,
N2089,N2090,N2091,N2092,N2093,N2094,N2095,N2096,N2097,N2098,
N2099,N2100,N2101,N2102,N2103,N2104,N2105,N2106,N2107,N2108,
N2109,N2110,N2111,N2112,N2113,N2114,N2115,N2116,N2117,N2118,
N2119,N2120,N2121,N2122,N2123,N2124,N2125,N2126,N2127,N2128,
N2129,N2130,N2131,N2132,N2133,N2134,N2135,N2136,N2137,N2138,
N2139,N2140,N2141,N2142,N2143,N2144,N2145,N2146,N2147,N2148,
N2149,N2150,N2151,N2152,N2153,N2154,N2155,N2156,N2157,N2158,
N2159,N2160,N2161,N2162,N2163,N2164,N2165,N2166,N2167,N2168,
N2169,N2170,N2171,N2172,N2173,N2174,N2175,N2176,N2177,N2178,
N2179,N2180,N2181,N2182,N2183,N2184,N2185,N2186,N2187,N2188,
N2189,N2190,N2191,N2192,N2193,N2194,N2195,N2196,N2197,N2198,
N2199,N2200,N2201,N2202,N2203,N2204,N2205,N2206,N2207,N2208,
N2209,N2210,N2211,N2212,N2213,N2214,N2215,N2216,N2217,N2218,
N2219,N2220,N2221,N2222,N2223,N2224,N2225,N2226,N2227,N2228,
N2229,N2230,N2231,N2232,N2233,N2234,N2235,N2236,N2237,N2238,
N2239,N2240,N2241,N2242,N2243,N2244,N2245,N2246,N2247,N2248,
N2249,N2250,N2251,N2252,N2253,N2254,N2255,N2256,N2257,N2258,
N2259,N2260,N2261,N2262,N2263,N2264,N2265,N2266,N2267,N2268,
N2269,N2270,N2271,N2272,N2273,N2274,N2275,N2276,N2277,N2278,
N2279,N2280,N2281,N2282,N2283,N2284,N2285,N2286,N2287,N2288,
N2289,N2290,N2291,N2292,N2293,N2294,N2295,N2296,N2297,N2298,
N2299,N2300,N2301,N2302,N2303,N2304,N2305,N2306,N2307,N2308,
N2309,N2310,N2311,N2312,N2313,N2314,N2315,N2316,N2317,N2318,
N2319,N2320,N2321,N2322,N2323,N2324,N2325,N2326,N2327,N2328,
N2329,N2330,N2331,N2332,N2333,N2334,N2335,N2336,N2337,N2338,
N2339,N2340,N2341,N2342,N2343,N2344,N2345,N2346,N2347,N2348,
N2349,N2350,N2351,N2352,N2353,N2354,N2355,N2356,N2357,N2358,
N2359,N2360,N2361,N2362,N2363,N2364,N2365,N2366,N2367,N2368,
N2369,N2370,N2371,N2372,N2373,N2374,N2375,N2376,N2377,N2378,
N2379,N2380,N2381,N2382,N2383,N2384,N2385,N2386,N2387,N2388,
N2389,N2390,N2391,N2392,N2393,N2394,N2395,N2396,N2397,N2398,
N2399,N2400,N2401,N2402,N2403,N2404,N2405,N2406,N2407,N2408,
N2409,N2410,N2411,N2412,N2413,N2414,N2415,N2416,N2417,N2418,
N2419,N2420,N2421,N2422,N2423,N2424,N2425,N2426,N2427,N2428,
N2429,N2430,N2431,N2432,N2433,N2434,N2435,N2436,N2437,N2438,
N2439,N2440,N2441,N2442,N2443,N2444,N2445,N2446,N2447,N2448,
N2449,N2450,N2451,N2452,N2453,N2454,N2455,N2456,N2457,N2458,
N2459,N2460,N2461,N2462,N2463,N2464,N2465,N2466,N2467,N2468,
N2469,N2470,N2471,N2472,N2473,N2474,N2475,N2476,N2477,N2478,
N2479,N2480,N2481,N2482,N2483,N2484,N2485,N2486,N2487,N2488,
N2489,N2490,N2491,N2492,N2493,N2494,N2495,N2496,N2497,N2498,
N2499,N2500,N2501,N2502,N2503,N2504,N2505,N2506,N2507,N2508,
N2509,N2510,N2511,N2512,N2513,N2514,N2515,N2516,N2517,N2518,
N2519,N2520,N2521,N2522,N2523,N2524,N2525,N2526,N2527,N2528,
N2529,N2530,N2531,N2532,N2533,N2534,N2535,N2536,N2537,N2538,
N2539,N2540,N2541,N2542,N2543,N2544,N2545,N2546,N2547,N2548,
N2549,N2550,N2551,N2552,N2553,N2554,N2555,N2556,N2557,N2558,
N2559,N2560,N2561,N2562,N2563,N2564,N2565,N2566,N2567,N2568,
N2569,N2570,N2571,N2572,N2573,N2574,N2575,N2576,N2577,N2578,
N2579,N2580,N2581,N2582,N2583,N2584,N2585,N2586,N2587,N2588,
N2589,N2590,N2591,N2592,N2593,N2594,N2595,N2596,N2597,N2598,
N2599,N2600,N2601,N2602,N2603,N2604,N2605,N2606,N2607,N2608,
N2609,N2610,N2611,N2612,N2613,N2614,N2615,N2616,N2617,N2618,
N2619,N2620,N2621,N2622,N2623,N2624,N2625,N2626,N2627,N2628,
N2629,N2630,N2631,N2632,N2633,N2634,N2635,N2636,N2637,N2638,
N2639,N2640,N2641,N2642,N2643,N2644,N2645,N2646,N2647,N2648,
N2649,N2650,N2651,N2652,N2653,N2654,N2655,N2656,N2657,N2658,
N2659,N2660,N2661,N2662,N2663,N2664,N2665,N2666,N2667,N2668,
N2669,N2670,N2671,N2672,N2673,N2674,N2675,N2676,N2677,N2678,
N2679,N2680,N2681,N2682,N2683,N2684,N2685,N2686,N2687,N2688,
N2689,N2690,N2691,N2692,N2693,N2694,N2695,N2696,N2697,N2698,
N2699,N2700,N2701,N2702,N2703,N2704,N2705,N2706,N2707,N2708,
N2709,N2710,N2711,N2712,N2713,N2714,N2715,N2716,N2717,N2718,
N2719,N2720,N2721,N2722,N2723,N2724,N2725,N2726,N2727,N2728,
N2729,N2730,N2731,N2732,N2733,N2734,N2735,N2736,N2737,N2738,
N2739,N2740,N2741,N2742,N2743,N2744,N2745,N2746,N2747,N2748,
N2749,N2750,N2751,N2752,N2753,N2754,N2755,N2756,N2757,N2758,
N2759,N2760,N2761,N2762,N2763,N2764,N2765,N2766,N2767,N2768,
N2769,N2770,N2771,N2772,N2773,N2774,N2775,N2776,N2777,N2778,
N2779,N2780,N2781,N2782,N2783,N2784,N2785,N2786,N2787,N2788,
N2789,N2790,N2791,N2792,N2793,N2794,N2795,N2796,N2797,N2798,
N2799,N2800,N2801,N2802,N2803,N2804,N2805,N2806,N2807,N2808,
N2809,N2810,N2811,N2812,N2813,N2814,N2815,N2816,N2817,N2818,
N2819,N2820,N2821,N2822,N2823,N2824,N2825,N2826,N2827,N2828,
N2829,N2830,N2831,N2832,N2833,N2834,N2835,N2836,N2837,N2838,
N2839,N2840,N2841,N2842,N2843,N2844,N2845,N2846,N2847,N2848,
N2849,N2850,N2851,N2852,N2853,N2854,N2855,N2856,N2857,N2858,
N2859,N2860,N2861,N2862,N2863,N2864,N2865,N2866,N2867,N2868,
N2869,N2870,N2871,N2872,N2873,N2874,N2875,N2876,N2877,N2878,
N2879,N2880,N2881,N2882,N2883,N2884,N2885,N2886,N2887,N2888,
N2889,N2890,N2891,N2892,N2893,N2894,N2895,N2896,N2897,N2898,
N2899,N2900,N2901,N2902,N2903,N2904,N2905,N2906,N2907,N2908,
N2909,N2910,N2911,N2912,N2913,N2914,N2915,N2916,N2917,N2918,
N2919,N2920,N2921,N2922,N2923,N2924,N2925,N2926,N2927,N2928,
N2929,N2930,N2931,N2932,N2933,N2934,N2935,N2936,N2937,N2938,
N2939,N2940,N2941,N2942,N2943,N2944,N2945,N2946,N2947,N2948,
N2949,N2950,N2951,N2952,N2953,N2954,N2955,N2956,N2957,N2958,
N2959,N2960,N2961,N2962,N2963,N2964,N2965,N2966,N2967,N2968,
N2969,N2970,N2971,N2972,N2973,N2974,N2975,N2976,N2977,N2978,
N2979,N2980,N2981,N2982,N2983,N2984,N2985,N2986,N2987,N2988,
N2989,N2990,N2991,N2992,N2993,N2994,N2995,N2996,N2997,N2998,
N2999,N3000,N3001,N3002,N3003,N3004,N3005,N3006,N3007,N3008,
N3009,N3010,N3011,N3012,N3013,N3014,N3015,N3016,N3017,N3018,
N3019,N3020,N3021,N3022,N3023,N3024,N3025,N3026,N3027,N3028,
N3029,N3030,N3031,N3032,N3033,N3034,N3035,N3036,N3037,N3038,
N3039,N3040,N3041,N3042,N3043,N3044,N3045,N3046,N3047,N3048,
N3049,N3050,N3051,N3052,N3053,N3054,N3055,N3056,N3057,N3058,
N3059,N3060,N3061,N3062,N3063,N3064,N3065,N3066,N3067,N3068,
N3069,N3070,N3071,N3072,N3073,N3074,N3075,N3076,N3077,N3078,
N3079,N3080,N3081,N3082,N3083,N3084,N3085,N3086,N3087,N3088,
N3089,N3090,N3091,N3092,N3093,N3094,N3095,N3096,N3097,N3098,
N3099,N3100,N3101,N3102,N3103,N3104,N3105,N3106,N3107,N3108,
N3109,N3110,N3111,N3112,N3113,N3114,N3115,N3116,N3117,N3118,
N3119,N3120,N3121,N3122,N3123,N3124,N3125,N3126,N3127,N3128,
N3129,N3130,N3131,N3132,N3133,N3134,N3135,N3136,N3137,N3138,
N3139,N3140,N3141,N3142,N3143,N3144,N3145,N3146,N3147,N3148,
N3149,N3150,N3151,N3152,N3153,N3154,N3155,N3156,N3157,N3158,
N3159,N3160,N3161,N3162,N3163,N3164,N3165,N3166,N3167,N3168,
N3169,N3170,N3171,N3172,N3173,N3174,N3175,N3176,N3177,N3178,
N3179,N3180,N3181,N3182,N3183,N3184,N3185,N3186,N3187,N3188,
N3189,N3190,N3191,N3192,N3193,N3194,N3195,N3196,N3197,N3198,
N3199,N3200,N3201,N3202,N3203,N3204,N3205,N3206,N3207,N3208,
N3209,N3210,N3211,N3212,N3213,N3214,N3215,N3216,N3217,N3218,
N3219,N3220,N3221,N3222,N3223,N3224,N3225,N3226,N3227,N3228,
N3229,N3230,N3231,N3232,N3233,N3234,N3235,N3236,N3237,N3238,
N3239,N3240,N3241,N3242,N3243,N3244,N3245,N3246,N3247,N3248,
N3249,N3250,N3251,N3252,N3253,N3254,N3255,N3256,N3257,N3258,
N3259,N3260,N3261,N3262,N3263,N3264,N3265,N3266,N3267,N3268,
N3269,N3270,N3271,N3272,N3273,N3274,N3275,N3276,N3277,N3278,
N3279,N3280,N3281,N3282,N3283,N3284,N3285,N3286,N3287,N3288,
N3289,N3290,N3291,N3292,N3293,N3294,N3295,N3296,N3297,N3298,
N3299,N3300,N3301,N3302,N3303,N3304,N3305,N3306,N3307,N3308,
N3309,N3310,N3311,N3312,N3313,N3314,N3315,N3316,N3317,N3318,
N3319,N3320,N3321,N3322,N3323,N3324,N3325,N3326,N3327,N3328,
N3329,N3330,N3331,N3332,N3333,N3334,N3335,N3336,N3337,N3338,
N3339,N3340,N3341,N3342,N3343,N3344,N3345,N3346,N3347,N3348,
N3349,N3350,N3351,N3352,N3353,N3354,N3355,N3356,N3357,N3358,
N3359,N3360,N3361,N3362,N3363,N3364,N3365,N3366,N3367,N3368,
N3369,N3370,N3371,N3372,N3373,N3374,N3375,N3376,N3377,N3378,
N3379,N3380,N3381,N3382,N3383,N3384,N3385,N3386,N3387,N3388,
N3389,N3390,N3391,N3392,N3393,N3394,N3395,N3396,N3397,N3398,
N3399,N3400,N3401,N3402,N3403,N3404,N3405,N3406,N3407,N3408,
N3409,N3410,N3411,N3412,N3413,N3414,N3415,N3416,N3417,N3418,
N3419,N3420,N3421,N3422,N3423,N3424,N3425,N3426,N3427,N3428,
N3429,N3430,N3431,N3432,N3433,N3434,N3435,N3436,N3437,N3438,
N3439,N3440,N3441,N3442,N3443,N3444,N3445,N3446,N3447,N3448,
N3449,N3450,N3451,N3452,N3453,N3454,N3455,N3456,N3457,N3458,
N3459,N3460,N3461,N3462,N3463,N3464,N3465,N3466,N3467,N3468,
N3469,N3470,N3471,N3472,N3473,N3474,N3475,N3476,N3477,N3478,
N3479,N3480,N3481,N3482,N3483,N3484,N3485,N3486,N3487,N3488,
N3489,N3490,N3491,N3492,N3493,N3494,N3495,N3496,N3497,N3498,
N3499,N3500,N3501,N3502,N3503,N3504,N3505,N3506,N3507,N3508,
N3509,N3510,N3511,N3512,N3513,N3514,N3515,N3516,N3517,N3518,
N3519,N3520,N3521,N3522,N3523,N3524,N3525,N3526,N3527,N3528,
N3529,N3530,N3531,N3532,N3533,N3534,N3535,N3536,N3537,N3538,
N3539,N3540,N3541,N3542,N3543,N3544,N3545,N3546,N3547,N3548,
N3549,N3550,N3551,N3552,N3553,N3554,N3555,N3556,N3557,N3558,
N3559,N3560,N3561,N3562,N3563,N3564,N3565,N3566,N3567,N3568,
N3569,N3570,N3571,N3572,N3573,N3574,N3575,N3576,N3577,N3578,
N3579,N3580,N3581,N3582,N3583,N3584,N3585,N3586,N3587,N3588,
N3589,N3590,N3591,N3592,N3593,N3594,N3595,N3596,N3597,N3598,
N3599,N3600,N3601,N3602,N3603,N3604,N3605,N3606,N3607,N3608,
N3609,N3610,N3611,N3612,N3613,N3614,N3615,N3616,N3617,N3618,
N3619,N3620,N3621,N3622,N3623,N3624,N3625,N3626,N3627,N3628,
N3629,N3630,N3631,N3632,N3633,N3634,N3635,N3636,N3637,N3638,
N3639,N3640,N3641,N3642,N3643,N3644,N3645,N3646,N3647,N3648,
N3649,N3650,N3651,N3652,N3653,N3654,N3655,N3656,N3657,N3658,
N3659,N3660,N3661,N3662,N3663,N3664,N3665,N3666,N3667,N3668,
N3669,N3670,N3671,N3672,N3673,N3674,N3675,N3676,N3677,N3678,
N3679,N3680,N3681,N3682,N3683,N3684,N3685,N3686,N3687,N3688,
N3689,N3690,N3691,N3692,N3693,N3694,N3695,N3696,N3697,N3698,
N3699,N3700,N3701,N3702,N3703,N3704,N3705,N3706,N3707,N3708,
N3709,N3710,N3711,N3712,N3713,N3714,N3715,N3716,N3717,N3718,
N3719,N3720,N3721,N3722,N3723,N3724,N3725,N3726,N3727,N3728,
N3729,N3730,N3731,N3732,N3733,N3734,N3735,N3736,N3737,N3738,
N3739,N3740,N3741,N3742,N3743,N3744,N3745,N3746,N3747,N3748,
N3749,N3750,N3751,N3752,N3753,N3754,N3755,N3756,N3757,N3758,
N3759,N3760,N3761,N3762,N3763,N3764,N3765,N3766,N3767,N3768,
N3769,N3770,N3771,N3772,N3773,N3774,N3775,N3776,N3777,N3778,
N3779,N3780,N3781,N3782,N3783,N3784,N3785,N3786,N3787,N3788,
N3789,N3790,N3791,N3792,N3793,N3794,N3795,N3796,N3797,N3798,
N3799,N3800,N3801,N3802,N3803,N3804,N3805,N3806,N3807,N3808,
N3809,N3810,N3811,N3812,N3813,N3814,N3815,N3816,N3817,N3818,
N3819,N3820,N3821,N3822,N3823,N3824,N3825,N3826,N3827,N3828,
N3829,N3830,N3831,N3832,N3833,N3834,N3835,N3836,N3837,N3838,
N3839,N3840,N3841,N3842,N3843,N3844,N3845,N3846,N3847,N3848,
N3849,N3850,N3851,N3852,N3853,N3854,N3855,N3856,N3857,N3858,
N3859,N3860,N3861,N3862,N3863,N3864,N3865,N3866,N3867,N3868,
N3869,N3870,N3871,N3872,N3873,N3874,N3875,N3876,N3877,N3878,
N3879,N3880,N3881,N3882,N3883,N3884,N3885,N3886,N3887,N3888,
N3889,N3890,N3891,N3892,N3893,N3894,N3895,N3896,N3897,N3898,
N3899,N3900,N3901,N3902,N3903,N3904,N3905,N3906,N3907,N3908,
N3909,N3910,N3911,N3912,N3913,N3914,N3915,N3916,N3917,N3918,
N3919,N3920,N3921,N3922,N3923,N3924,N3925,N3926,N3927,N3928,
N3929,N3930,N3931,N3932,N3933,N3934,N3935,N3936,N3937,N3938,
N3939,N3940,N3941,N3942,N3943,N3944,N3945,N3946,N3947,N3948,
N3949,N3950,N3951,N3952,N3953,N3954,N3955,N3956,N3957,N3958,
N3959,N3960,N3961,N3962,N3963,N3964,N3965,N3966,N3967,N3968,
N3969,N3970,N3971,N3972,N3973,N3974,N3975,N3976,N3977,N3978,
N3979,N3980,N3981,N3982,N3983,N3984,N3985,N3986,N3987,N3988,
N3989,N3990,N3991,N3992,N3993,N3994,N3995,N3996,N3997,N3998,
N3999,N4000,N4001,N4002,N4003,N4004,N4005,N4006,N4007,N4008,
N4009,N4010,N4011,N4012,N4013,N4014,N4015,N4016,N4017,N4018,
N4019,N4020,N4021,N4022,N4023,N4024,N4025,N4026,N4027,N4028,
N4029,N4030,N4031,N4032,N4033,N4034,N4035,N4036,N4037,N4038,
N4039,N4040,N4041,N4042,N4043,N4044,N4045,N4046,N4047,N4048,
N4049,N4050,N4051,N4052,N4053,N4054,N4055,N4056,N4057,N4058,
N4059,N4060,N4061,N4062,N4063,N4064,N4065,N4066,N4067,N4068,
N4069,N4070,N4071,N4072,N4073,N4074,N4075,N4076,N4077,N4078,
N4079,N4080,N4081,N4082,N4083,N4084,N4085,N4086,N4087,N4088,
N4089,N4090,N4091,N4092,N4093,N4094,N4095,N4096,N4097,N4098,
N4099,N4100,N4101,N4102,N4103,N4104,N4105,N4106,N4107,N4108,
N4109,N4110,N4111,N4112,N4113,N4114,N4115,N4116,N4117,N4118,
N4119,N4120,N4121,N4122,N4123,N4124,N4125,N4126,N4127,N4128,
N4129,N4130,N4131,N4132,N4133,N4134,N4135,N4136,N4137,N4138,
N4139,N4140,N4141,N4142,N4143,N4144,N4145,N4146,N4147,N4148,
N4149,N4150,N4151,N4152,N4153,N4154,N4155,N4156,N4157,N4158,
N4159,N4160,N4161,N4162,N4163,N4164,N4165,N4166,N4167,N4168,
N4169,N4170,N4171,N4172,N4173,N4174,N4175,N4176,N4177,N4178,
N4179,N4180,N4181,N4182,N4183,N4184,N4185,N4186,N4187,N4188,
N4189,N4190,N4191,N4192,N4193,N4194,N4195,N4196,N4197,N4198,
N4199,N4200,N4201,N4202,N4203,N4204,N4205,N4206,N4207,N4208,
N4209,N4210,N4211,N4212,N4213,N4214,N4215,N4216,N4217,N4218,
N4219,N4220,N4221,N4222,N4223,N4224,N4225,N4226,N4227,N4228,
N4229,N4230,N4231,N4232,N4233,N4234,N4235,N4236,N4237,N4238,
N4239,N4240,N4241,N4242,N4243,N4244,N4245,N4246,N4247,N4248,
N4249,N4250,N4251,N4252,N4253,N4254,N4255,N4256,N4257,N4258,
N4259,N4260,N4261,N4262,N4263,N4264,N4265,N4266,N4267,N4268,
N4269,N4270,N4271,N4272,N4273,N4274,N4275,N4276,N4277,N4278,
N4279,N4280,N4281,N4282,N4283,N4284,N4285,N4286,N4287,N4288,
N4289,N4290,N4291,N4292,N4293,N4294,N4295,N4296,N4297,N4298,
N4299,N4300,N4301,N4302,N4303,N4304,N4305,N4306,N4307,N4308,
N4309,N4310,N4311,N4312,N4313,N4314,N4315,N4316,N4317,N4318,
N4319,N4320,N4321,N4322,N4323,N4324,N4325,N4326,N4327,N4328,
N4329,N4330,N4331,N4332,N4333,N4334,N4335,N4336,N4337,N4338,
N4339,N4340,N4341,N4342,N4343,N4344,N4345,N4346,N4347,N4348,
N4349,N4350,N4351,N4352,N4353,N4354,N4355,N4356,N4357,N4358,
N4359,N4360,N4361,N4362,N4363,N4364,N4365,N4366,N4367,N4368,
N4369,N4370,N4371,N4372,N4373,N4374,N4375,N4376,N4377,N4378,
N4379,N4380,N4381,N4382,N4383,N4384,N4385,N4386,N4387,N4388,
N4389,N4390,N4391,N4392,N4393,N4394,N4395,N4396,N4397,N4398,
N4399,N4400,N4401,N4402,N4403,N4404,N4405,N4406,N4407,N4408,
N4409,N4410,N4411,N4412,N4413,N4414,N4415,N4416,N4417,N4418,
N4419,N4420,N4421,N4422,N4423,N4424,N4425,N4426,N4427,N4428,
N4429,N4430,N4431,N4432,N4433,N4434,N4435,N4436,N4437,N4438,
N4439,N4440,N4441,N4442,N4443,N4444,N4445,N4446,N4447,N4448,
N4449,N4450,N4451,N4452,N4453,N4454,N4455,N4456,N4457,N4458,
N4459,N4460,N4461,N4462,N4463,N4464,N4465,N4466,N4467,N4468,
N4469,N4470,N4471,N4472,N4473,N4474,N4475,N4476,N4477,N4478,
N4479,N4480,N4481,N4482,N4483,N4484,N4485,N4486,N4487,N4488,
N4489,N4490,N4491,N4492,N4493,N4494,N4495,N4496,N4497,N4498,
N4499,N4500,N4501,N4502,N4503,N4504,N4505,N4506,N4507,N4508,
N4509,N4510,N4511,N4512,N4513,N4514,N4515,N4516,N4517,N4518,
N4519,N4520,N4521,N4522,N4523,N4524,N4525,N4526,N4527,N4528,
N4529,N4530,N4531,N4532,N4533,N4534,N4535,N4536,N4537,N4538,
N4539,N4540,N4541,N4542,N4543,N4544,N4545,N4546,N4547,N4548,
N4549,N4550,N4551,N4552,N4553,N4554,N4555,N4556,N4557,N4558,
N4559,N4560,N4561,N4562,N4563,N4564,N4565,N4566,N4567,N4568,
N4569,N4570,N4571,N4572,N4573,N4574,N4575,N4576,N4577,N4578,
N4579,N4580,N4581,N4582,N4583,N4584,N4585,N4586,N4587,N4588,
N4589,N4590,N4591,N4592,N4593,N4594,N4595,N4596,N4597,N4598,
N4599,N4600,N4601,N4602,N4603,N4604,N4605,N4606,N4607,N4608,
N4609,N4610,N4611,N4612,N4613,N4614,N4615,N4616,N4617,N4618,
N4619,N4620,N4621,N4622,N4623,N4624,N4625,N4626,N4627,N4628,
N4629,N4630,N4631,N4632,N4633,N4634,N4635,N4636,N4637,N4638,
N4639,N4640,N4641,N4642,N4643,N4644,N4645,N4646,N4647,N4648,
N4649,N4650,N4651,N4652,N4653,N4654,N4655,N4656,N4657,N4658,
N4659,N4660,N4661,N4662,N4663,N4664,N4665,N4666,N4667,N4668,
N4669,N4670,N4671,N4672,N4673,N4674,N4675,N4676,N4677,N4678,
N4679,N4680,N4681,N4682,N4683,N4684,N4685,N4686,N4687,N4688,
N4689,N4690,N4691,N4692,N4693,N4694,N4695,N4696,N4697,N4698,
N4699,N4700,N4701,N4702,N4703,N4704,N4705,N4706,N4707,N4708,
N4709,N4710,N4711,N4712,N4713,N4714,N4715,N4716,N4717,N4718,
N4719,N4720,N4721,N4722,N4723,N4724,N4725,N4726,N4727,N4728,
N4729,N4730,N4731,N4732,N4733,N4734,N4735,N4736,N4737,N4738,
N4739,N4740,N4741,N4742,N4743,N4744,N4745,N4746,N4747,N4748,
N4749,N4750,N4751,N4752,N4753,N4754,N4755,N4756,N4757,N4758,
N4759,N4760,N4761,N4762,N4763,N4764,N4765,N4766,N4767,N4768,
N4769,N4770,N4771,N4772,N4773,N4774,N4775,N4776,N4777,N4778,
N4779,N4780,N4781,N4782,N4783,N4784,N4785,N4786,N4787,N4788,
N4789,N4790,N4791,N4792,N4793,N4794,N4795,N4796,N4797,N4798,
N4799,N4800,N4801,N4802,N4803,N4804,N4805,N4806,N4807,N4808,
N4809,N4810,N4811,N4812,N4813,N4814,N4815,N4816,N4817,N4818,
N4819,N4820,N4821,N4822,N4823,N4824,N4825,N4826,N4827,N4828,
N4829,N4830,N4831,N4832,N4833,N4834,N4835,N4836,N4837,N4838,
N4839,N4840,N4841,N4842,N4843,N4844,N4845,N4846,N4847,N4848,
N4849,N4850,N4851,N4852,N4853,N4854,N4855,N4856,N4857,N4858,
N4859,N4860,N4861,N4862,N4863,N4864,N4865,N4866,N4867,N4868,
N4869,N4870,N4871,N4872,N4873,N4874,N4875,N4876,N4877,N4878,
N4879,N4880,N4881,N4882,N4883,N4884,N4885,N4886,N4887,N4888,
N4889,N4890,N4891,N4892,N4893,N4894,N4895,N4896,N4897,N4898,
N4899,N4900,N4901,N4902,N4903,N4904,N4905,N4906,N4907,N4908,
N4909,N4910,N4911,N4912,N4913,N4914,N4915,N4916,N4917,N4918,
N4919,N4920,N4921,N4922,N4923,N4924,N4925,N4926,N4927,N4928,
N4929,N4930,N4931,N4932,N4933,N4934,N4935,N4936,N4937,N4938,
N4939,N4940,N4941,N4942,N4943,N4944,N4945,N4946,N4947,N4948,
N4949,N4950,N4951,N4952,N4953,N4954,N4955,N4956,N4957,N4958,
N4959,N4960,N4961,N4962,N4963,N4964,N4965,N4966,N4967,N4968,
N4969,N4970,N4971,N4972,N4973,N4974,N4975,N4976,N4977,N4978,
N4979,N4980,N4981,N4982,N4983,N4984,N4985,N4986,N4987,N4988,
N4989,N4990,N4991,N4992,N4993,N4994,N4995,N4996,N4997,N4998,
N4999,N5000,N5001,N5002,N5003,N5004,N5005,N5006,N5007,N5008,
N5009,N5010,N5011,N5012,N5013,N5014,N5015,N5016,N5017,N5018,
N5019,N5020,N5021,N5022,N5023,N5024,N5025,N5026,N5027,N5028,
N5029,N5030,N5031,N5032,N5033,N5034,N5035,N5036,N5037,N5038,
N5039,N5040,N5041,N5042,N5043,N5044,N5045,N5046,N5047,N5048,
N5049,N5050,N5051,N5052,N5053,N5054,N5055,N5056,N5057,N5058,
N5059,N5060,N5061,N5062,N5063,N5064,N5065,N5066,N5067,N5068,
N5069,N5070,N5071,N5072,N5073,N5074,N5075,N5076,N5077,N5078,
N5079,N5080,N5081,N5082,N5083,N5084,N5085,N5086,N5087,N5088,
N5089,N5090,N5091,N5092,N5093,N5094,N5095,N5096,N5097,N5098,
N5099,N5100,N5101,N5102,N5103,N5104,N5105,N5106,N5107,N5108,
N5109,N5110,N5111,N5112,N5113,N5114,N5115,N5116,N5117,N5118,
N5119,N5120,N5121,N5122,N5123,N5124,N5125,N5126,N5127,N5128,
N5129,N5130,N5131,N5132,N5133,N5134,N5135,N5136,N5137,N5138,
N5139,N5140,N5141,N5142,N5143,N5144,N5145,N5146,N5147,N5148,
N5149,N5150,N5151,N5152,N5153,N5154,N5155,N5156,N5157,N5158,
N5159,N5160,N5161,N5162,N5163,N5164,N5165,N5166,N5167,N5168,
N5169,N5170,N5171,N5172,N5173,N5174,N5175,N5176,N5177,N5178,
N5179,N5180,N5181,N5182,N5183,N5184,N5185,N5186,N5187,N5188,
N5189,N5190,N5191,N5192,N5193,N5194,N5195,N5196,N5197,N5198,
N5199,N5200,N5201,N5202,N5203,N5204,N5205,N5206,N5207,N5208,
N5209,N5210,N5211,N5212,N5213,N5214,N5215,N5216,N5217,N5218,
N5219,N5220,N5221,N5222,N5223,N5224,N5225,N5226,N5227,N5228,
N5229,N5230,N5231,N5232,N5233,N5234,N5235,N5236,N5237,N5238,
N5239,N5240,N5241,N5242,N5243,N5244,N5245,N5246,N5247,N5248,
N5249,N5250,N5251,N5252,N5253,N5254,N5255,N5256,N5257,N5258,
N5259,N5260,N5261,N5262,N5263,N5264,N5265,N5266,N5267,N5268,
N5269,N5270,N5271,N5272,N5273,N5274,N5275,N5276,N5277,N5278,
N5279,N5280,N5281,N5282,N5283,N5284,N5285,N5286,N5287,N5288,
N5289,N5290,N5291,N5292,N5293,N5294,N5295,N5296,N5297,N5298,
N5299,N5300,N5301,N5302,N5303,N5304,N5305,N5306,N5307,N5308,
N5309,N5310,N5311,N5312,N5313,N5314,N5315,N5316,N5317,N5318,
N5319,N5320,N5321,N5322,N5323,N5324,N5325,N5326,N5327,N5328,
N5329,N5330,N5331,N5332,N5333,N5334,N5335,N5336,N5337,N5338,
N5339,N5340,N5341,N5342,N5343,N5344,N5345,N5346,N5347,N5348,
N5349,N5350,N5351,N5352,N5353,N5354,N5355,N5356,N5357,N5358,
N5359,N5360,N5361,N5362,N5363,N5364,N5365,N5366,N5367,N5368,
N5369,N5370,N5371,N5372,N5373,N5374,N5375,N5376,N5377,N5378,
N5379,N5380,N5381,N5382,N5383,N5384,N5385,N5386,N5387,N5388,
N5389,N5390,N5391,N5392,N5393,N5394,N5395,N5396,N5397,N5398,
N5399,N5400,N5401,N5402,N5403,N5404,N5405,N5406,N5407,N5408,
N5409,N5410,N5411,N5412,N5413,N5414,N5415,N5416,N5417,N5418,
N5419,N5420,N5421,N5422,N5423,N5424,N5425,N5426,N5427,N5428,
N5429,N5430,N5431,N5432,N5433,N5434,N5435,N5436,N5437,N5438,
N5439,N5440,N5441,N5442,N5443,N5444,N5445,N5446,N5447,N5448,
N5449,N5450,N5451,N5452,N5453,N5454,N5455,N5456,N5457,N5458,
N5459,N5460,N5461,N5462,N5463,N5464,N5465,N5466,N5467,N5468,
N5469,N5470,N5471,N5472,N5473,N5474,N5475,N5476,N5477,N5478,
N5479,N5480,N5481,N5482,N5483,N5484,N5485,N5486,N5487,N5488,
N5489,N5490,N5491,N5492,N5493,N5494,N5495,N5496,N5497,N5498,
N5499,N5500,N5501,N5502,N5503,N5504,N5505,N5506,N5507,N5508,
N5509,N5510,N5511,N5512,N5513,N5514,N5515,N5516,N5517,N5518,
N5519,N5520,N5521,N5522,N5523,N5524,N5525,N5526,N5527,N5528,
N5529,N5530,N5531,N5532,N5533,N5534,N5535,N5536,N5537,N5538,
N5539,N5540,N5541,N5542,N5543,N5544,N5545,N5546,N5547,N5548,
N5549,N5550,N5551,N5552,N5553,N5554,N5555,N5556,N5557,N5558,
N5559,N5560,N5561,N5562,N5563,N5564,N5565,N5566,N5567,N5568,
N5569,N5570,N5571,N5572,N5573,N5574,N5575,N5576,N5577,N5578,
N5579,N5580,N5581,N5582,N5583,N5584,N5585,N5586,N5587,N5588,
N5589,N5590,N5591,N5592,N5593,N5594,N5595,N5596,N5597,N5598,
N5599,N5600,N5601,N5602,N5603,N5604,N5605,N5606,N5607,N5608,
N5609,N5610,N5611,N5612,N5613,N5614,N5615,N5616,N5617,N5618,
N5619,N5620,N5621,N5622,N5623,N5624,N5625,N5626,N5627,N5628,
N5629,N5630,N5631,N5632,N5633,N5634,N5635,N5636,N5637,N5638,
N5639,N5640,N5641,N5642,N5643,N5644,N5645,N5646,N5647,N5648,
N5649,N5650,N5651,N5652,N5653,N5654,N5655,N5656,N5657,N5658,
N5659,N5660,N5661,N5662,N5663,N5664,N5665,N5666,N5667,N5668,
N5669,N5670,N5671,N5672,N5673,N5674,N5675,N5676,N5677,N5678,
N5679,N5680,N5681,N5682,N5683,N5684,N5685,N5686,N5687,N5688,
N5689,N5690,N5691,N5692,N5693,N5694,N5695,N5696,N5697,N5698,
N5699,N5700,N5701,N5702,N5703,N5704,N5705,N5706,N5707,N5708,
N5709,N5710,N5711,N5712,N5713,N5714,N5715,N5716,N5717,N5718,
N5719,N5720,N5721,N5722,N5723,N5724,N5725,N5726,N5727,N5728,
N5729,N5730,N5731,N5732,N5733,N5734,N5735,N5736,N5737,N5738,
N5739,N5740,N5741,N5742,N5743,N5744,N5745,N5746,N5747,N5748,
N5749,N5750,N5751,N5752,N5753,N5754,N5755,N5756,N5757,N5758,
N5759,N5760,N5761,N5762,N5763,N5764,N5765,N5766,N5767,N5768,
N5769,N5770,N5771,N5772,N5773,N5774,N5775,N5776,N5777,N5778,
N5779,N5780,N5781,N5782,N5783,N5784,N5785,N5786,N5787,N5788,
N5789,N5790,N5791,N5792,N5793,N5794,N5795,N5796,N5797,N5798,
N5799,N5800,N5801,N5802,N5803,N5804,N5805,N5806,N5807,N5808,
N5809,N5810,N5811,N5812,N5813,N5814,N5815,N5816,N5817,N5818,
N5819,N5820,N5821,N5822,N5823,N5824,N5825,N5826,N5827,N5828,
N5829,N5830,N5831,N5832,N5833,N5834,N5835,N5836,N5837,N5838,
N5839,N5840,N5841,N5842,N5843,N5844,N5845,N5846,N5847,N5848,
N5849,N5850,N5851,N5852,N5853,N5854,N5855,N5856,N5857,N5858,
N5859,N5860,N5861,N5862,N5863,N5864,N5865,N5866,N5867,N5868,
N5869,N5870,N5871,N5872,N5873,N5874,N5875,N5876,N5877,N5878,
N5879,N5880,N5881,N5882,N5883,N5884,N5885,N5886,N5887,N5888,
N5889,N5890,N5891,N5892,N5893,N5894,N5895,N5896,N5897,N5898,
N5899,N5900,N5901,N5902,N5903,N5904,N5905,N5906,N5907,N5908,
N5909,N5910,N5911,N5912,N5913,N5914,N5915,N5916,N5917,N5918,
N5919,N5920,N5921,N5922,N5923,N5924,N5925,N5926,N5927,N5928,
N5929,N5930,N5931,N5932,N5933,N5934,N5935,N5936,N5937,N5938,
N5939,N5940,N5941,N5942,N5943,N5944,N5945,N5946,N5947,N5948,
N5949,N5950,N5951,N5952,N5953,N5954,N5955,N5956,N5957,N5958,
N5959,N5960,N5961,N5962,N5963,N5964,N5965,N5966,N5967,N5968,
N5969,N5970,N5971,N5972,N5973,N5974,N5975,N5976,N5977,N5978,
N5979,N5980,N5981,N5982,N5983,N5984,N5985,N5986,N5987,N5988,
N5989,N5990,N5991,N5992,N5993,N5994,N5995,N5996,N5997,N5998,
N5999,N6000,N6001,N6002,N6003,N6004,N6005,N6006,N6007,N6008,
N6009,N6010,N6011,N6012,N6013,N6014,N6015,N6016,N6017,N6018,
N6019,N6020,N6021,N6022,N6023,N6024,N6025,N6026,N6027,N6028,
N6029,N6030,N6031,N6032,N6033,N6034,N6035,N6036,N6037,N6038,
N6039,N6040,N6041,N6042,N6043,N6044,N6045,N6046,N6047,N6048,
N6049,N6050,N6051,N6052,N6053,N6054,N6055,N6056,N6057,N6058,
N6059,N6060,N6061,N6062,N6063,N6064,N6065,N6066,N6067,N6068,
N6069,N6070,N6071,N6072,N6073,N6074,N6075,N6076,N6077,N6078,
N6079,N6080,N6081,N6082,N6083,N6084,N6085,N6086,N6087,N6088,
N6089,N6090,N6091,N6092,N6093,N6094,N6095,N6096,N6097,N6098,
N6099,N6100,N6101,N6102,N6103,N6104,N6105,N6106,N6107,N6108,
N6109,N6110,N6111,N6112,N6113,N6114,N6115,N6116,N6117,N6118,
N6119,N6120,N6121,N6122,N6123,N6124,N6125,N6126,N6127,N6128,
N6129,N6130,N6131,N6132,N6133,N6134,N6135,N6136,N6137,N6138,
N6139,N6140,N6141,N6142,N6143,N6144,N6145,N6146,N6147,N6148,
N6149,N6150,N6151,N6152,N6153,N6154,N6155,N6156,N6157,N6158,
N6159,N6160,N6161,N6162,N6163,N6164,N6165,N6166,N6167,N6168,
N6169,N6170,N6171,N6172,N6173,N6174,N6175,N6176,N6177,N6178,
N6179,N6180,N6181,N6182,N6183,N6184,N6185,N6186,N6187,N6188,
N6189,N6190,N6191,N6192,N6193,N6194,N6195,N6196,N6197,N6198,
N6199,N6200,N6201,N6202,N6203,N6204,N6205,N6206,N6207,N6208,
N6209,N6210,N6211,N6212,N6213,N6214,N6215,N6216,N6217,N6218,
N6219,N6220,N6221,N6222,N6223,N6224,N6225,N6226,N6227,N6228,
N6229,N6230,N6231,N6232,N6233,N6234,N6235,N6236,N6237,N6238,
N6239,N6240,N6241,N6242,N6243,N6244,N6245,N6246,N6247,N6248,
N6249,N6250,N6251,N6252,N6253,N6254,N6255,N6256,N6257,N6258,
N6259,N6260,N6261,N6262,N6263,N6264,N6265,N6266,N6267,N6268,
N6269,N6270,N6271,N6272,N6273,N6274,N6275,N6276,N6277,N6278,
N6279,N6280,N6281,N6282,N6283,N6284,N6285,N6286,N6287,N6288,
N6289,N6290,N6291,N6292,N6293,N6294,N6295,N6296,N6297,N6298,
N6299,N6300,N6301,N6302,N6303,N6304,N6305,N6306,N6307,N6308,
N6309,N6310,N6311,N6312,N6313,N6314,N6315,N6316,N6317,N6318,
N6319,N6320,N6321,N6322,N6323,N6324,N6325,N6326,N6327,N6328,
N6329,N6330,N6331,N6332,N6333,N6334,N6335,N6336,N6337,N6338,
N6339,N6340,N6341,N6342,N6343,N6344,N6345,N6346,N6347,N6348,
N6349,N6350,N6351,N6352,N6353,N6354,N6355,N6356,N6357,N6358,
N6359,N6360,N6361,N6362,N6363,N6364,N6365,N6366,N6367,N6368,
N6369,N6370,N6371,N6372,N6373,N6374,N6375,N6376,N6377,N6378,
N6379,N6380,N6381,N6382,N6383,N6384,N6385,N6386,N6387,N6388,
N6389,N6390,N6391,N6392,N6393,N6394,N6395,N6396,N6397,N6398,
N6399,N6400,N6401,N6402,N6403,N6404,N6405,N6406,N6407,N6408,
N6409,N6410,N6411,N6412,N6413,N6414,N6415,N6416,N6417,N6418,
N6419,N6420,N6421,N6422,N6423,N6424,N6425,N6426,N6427,N6428,
N6429,N6430,N6431,N6432,N6433,N6434,N6435,N6436,N6437,N6438,
N6439,N6440,N6441,N6442,N6443,N6444,N6445,N6446,N6447,N6448,
N6449,N6450,N6451,N6452,N6453,N6454,N6455,N6456,N6457,N6458,
N6459,N6460,N6461,N6462,N6463,N6464,N6465,N6466,N6467,N6468,
N6469,N6470,N6471,N6472,N6473,N6474,N6475,N6476,N6477,N6478,
N6479,N6480,N6481,N6482,N6483,N6484,N6485,N6486,N6487,N6488,
N6489,N6490,N6491,N6492,N6493,N6494,N6495,N6496,N6497,N6498,
N6499,N6500,N6501,N6502,N6503,N6504,N6505,N6506,N6507,N6508,
N6509,N6510,N6511,N6512,N6513,N6514,N6515,N6516,N6517,N6518,
N6519,N6520,N6521,N6522,N6523,N6524,N6525,N6526,N6527,N6528,
N6529,N6530,N6531,N6532,N6533,N6534,N6535,N6536,N6537,N6538,
N6539,N6540,N6541,N6542,N6543,N6544,N6545,N6546,N6547,N6548,
N6549,N6550,N6551,N6552,N6553,N6554,N6555,N6556,N6557,N6558,
N6559,N6560,N6561,N6562,N6563,N6564,N6565,N6566,N6567,N6568,
N6569,N6570,N6571,N6572,N6573,N6574,N6575,N6576,N6577,N6578,
N6579,N6580,N6581,N6582,N6583,N6584,N6585,N6586,N6587,N6588,
N6589,N6590,N6591,N6592,N6593,N6594,N6595,N6596,N6597,N6598,
N6599,N6600,N6601,N6602,N6603,N6604,N6605,N6606,N6607,N6608,
N6609,N6610,N6611,N6612,N6613,N6614,N6615,N6616,N6617,N6618,
N6619,N6620,N6621,N6622,N6623,N6624,N6625,N6626,N6627,N6628,
N6629,N6630,N6631,N6632,N6633,N6634,N6635,N6636,N6637,N6638,
N6639,N6640,N6641,N6642,N6643,N6644,N6645,N6646,N6647,N6648,
N6649,N6650,N6651,N6652,N6653,N6654,N6655,N6656,N6657,N6658,
N6659,N6660,N6661,N6662,N6663,N6664,N6665,N6666,N6667,N6668,
N6669,N6670,N6671,N6672,N6673,N6674,N6675,N6676,N6677,N6678,
N6679,N6680,N6681,N6682,N6683,N6684,N6685,N6686,N6687,N6688,
N6689,N6690,N6691,N6692,N6693,N6694,N6695,N6696,N6697,N6698,
N6699,N6700,N6701,N6702,N6703,N6704,N6705,N6706,N6707,N6708,
N6709,N6710,N6711,N6712,N6713,N6714,N6715,N6716,N6717,N6718,
N6719,N6720,N6721,N6722,N6723,N6724,N6725,N6726,N6727,N6728,
N6729,N6730,N6731,N6732,N6733,N6734,N6735,N6736,N6737,N6738,
N6739,N6740,N6741,N6742,N6743,N6744,N6745,N6746,N6747,N6748,
N6749,N6750,N6751,N6752,N6753,N6754,N6755,N6756,N6757,N6758,
N6759,N6760,N6761,N6762,N6763,N6764,N6765,N6766,N6767,N6768,
N6769,N6770,N6771,N6772,N6773,N6774,N6775,N6776,N6777,N6778,
N6779,N6780,N6781,N6782,N6783,N6784,N6785,N6786,N6787,N6788,
N6789,N6790,N6791,N6792,N6793,N6794,N6795,N6796,N6797,N6798,
N6799,N6800,N6801,N6802,N6803,N6804,N6805,N6806,N6807,N6808,
N6809,N6810,N6811,N6812,N6813,N6814,N6815,N6816,N6817,N6818,
N6819,N6820,N6821,N6822,N6823,N6824,N6825,N6826,N6827,N6828,
N6829,N6830,N6831,N6832,N6833,N6834,N6835,N6836,N6837,N6838,
N6839,N6840,N6841,N6842,N6843,N6844,N6845,N6846,N6847,N6848,
N6849,N6850,N6851,N6852,N6853,N6854,N6855,N6856,N6857,N6858,
N6859,N6860,N6861,N6862,N6863,N6864,N6865,N6866,N6867,N6868,
N6869,N6870,N6871,N6872,N6873,N6874,N6875,N6876,N6877,N6878,
N6879,N6880,N6881,N6882,N6883,N6884,N6885,N6886,N6887,N6888,
N6889,N6890,N6891,N6892,N6893,N6894,N6895,N6896,N6897,N6898,
N6899,N6900,N6901,N6902,N6903,N6904,N6905,N6906,N6907,N6908,
N6909,N6910,N6911,N6912,N6913,N6914,N6915,N6916,N6917,N6918,
N6919,N6920,N6921,N6922,N6923,N6924,N6925,N6926,N6927,N6928,
N6929,N6930,N6931,N6932,N6933,N6934,N6935,N6936,N6937,N6938,
N6939,N6940,N6941,N6942,N6943,N6944,N6945,N6946,N6947,N6948,
N6949,N6950,N6951,N6952,N6953,N6954,N6955,N6956,N6957,N6958,
N6959,N6960,N6961,N6962,N6963,N6964,N6965,N6966,N6967,N6968,
N6969,N6970,N6971,N6972,N6973,N6974,N6975,N6976,N6977,N6978,
N6979,N6980,N6981,N6982,N6983,N6984,N6985,N6986,N6987,N6988,
N6989,N6990,N6991,N6992,N6993,N6994,N6995,N6996,N6997,N6998,
N6999,N7000,N7001,N7002,N7003,N7004,N7005,N7006,N7007,N7008,
N7009,N7010,N7011,N7012,N7013,N7014,N7015,N7016,N7017,N7018,
N7019,N7020,N7021,N7022,N7023,N7024,N7025,N7026,N7027,N7028,
N7029,N7030,N7031,N7032,N7033,N7034,N7035,N7036,N7037,N7038,
N7039,N7040,N7041,N7042,N7043,N7044,N7045,N7046,N7047,N7048,
N7049,N7050,N7051,N7052,N7053,N7054,N7055,N7056,N7057,N7058,
N7059,N7060,N7061,N7062,N7063,N7064,N7065,N7066,N7067,N7068,
N7069,N7070,N7071,N7072,N7073,N7074,N7075,N7076,N7077,N7078,
N7079,N7080,N7081,N7082,N7083,N7084,N7085,N7086,N7087,N7088,
N7089,N7090,N7091,N7092,N7093,N7094,N7095,N7096,N7097,N7098,
N7099,N7100,N7101,N7102,N7103,N7104,N7105,N7106,N7107,N7108,
N7109,N7110,N7111,N7112,N7113,N7114,N7115,N7116,N7117,N7118,
N7119,N7120,N7121,N7122,N7123,N7124,N7125,N7126,N7127,N7128,
N7129,N7130,N7131,N7132,N7133,N7134,N7135,N7136,N7137,N7138,
N7139,N7140,N7141,N7142,N7143,N7144,N7145,N7146,N7147,N7148,
N7149,N7150,N7151,N7152,N7153,N7154,N7155,N7156,N7157,N7158,
N7159,N7160,N7161,N7162,N7163,N7164,N7165,N7166,N7167,N7168,
N7169,N7170,N7171,N7172,N7173,N7174,N7175,N7176,N7177,N7178,
N7179,N7180,N7181,N7182,N7183,N7184,N7185,N7186,N7187,N7188,
N7189,N7190,N7191,N7192,N7193,N7194,N7195,N7196,N7197,N7198,
N7199,N7200,N7201,N7202,N7203,N7204,N7205,N7206,N7207,N7208,
N7209,N7210,N7211,N7212,N7213,N7214,N7215,N7216,N7217,N7218,
N7219,N7220,N7221,N7222,N7223,N7224,N7225,N7226,N7227,N7228,
N7229,N7230,N7231,N7232,N7233,N7234,N7235,N7236,N7237,N7238,
N7239,N7240,N7241,N7242,N7243,N7244,N7245,N7246,N7247,N7248,
N7249,N7250,N7251,N7252,N7253,N7254,N7255,N7256,N7257,N7258,
N7259,N7260,N7261,N7262,N7263,N7264,N7265,N7266,N7267,N7268,
N7269,N7270,N7271,N7272,N7273,N7274,N7275,N7276,N7277,N7278,
N7279,N7280,N7281,N7282,N7283,N7284,N7285,N7286,N7287,N7288,
N7289,N7290,N7291,N7292,N7293,N7294,N7295,N7296,N7297,N7298,
N7299,N7300,N7301,N7302,N7303,N7304,N7305,N7306,N7307,N7308,
N7309,N7310,N7311,N7312,N7313,N7314,N7315,N7316,N7317,N7318,
N7319,N7320,N7321,N7322,N7323,N7324,N7325,N7326,N7327,N7328,
N7329,N7330,N7331,N7332,N7333,N7334,N7335,N7336,N7337,N7338,
N7339,N7340,N7341,N7342,N7343,N7344,N7345,N7346,N7347,N7348,
N7349,N7350,N7351,N7352,N7353,N7354,N7355,N7356,N7357,N7358,
N7359,N7360,N7361,N7362,N7363,N7364,N7365,N7366,N7367,N7368,
N7369,N7370,N7371,N7372,N7373,N7374,N7375,N7376,N7377,N7378,
N7379,N7380,N7381,N7382,N7383,N7384,N7385,N7386,N7387,N7388,
N7389,N7390,N7391,N7392,N7393,N7394,N7395,N7396,N7397,N7398,
N7399,N7400,N7401,N7402,N7403,N7404,N7405,N7406,N7407,N7408,
N7409,N7410,N7411,N7412,N7413,N7414,N7415,N7416,N7417,N7418,
N7419,N7420,N7421,N7422,N7423,N7424,N7425,N7426,N7427,N7428,
N7429,N7430,N7431,N7432,N7433,N7434,N7435,N7436,N7437,N7438,
N7439,N7440,N7441,N7442,N7443,N7444,N7445,N7446,N7447,N7448,
N7449,N7450,N7451,N7452,N7453,N7454,N7455,N7456,N7457,N7458,
N7459,N7460,N7461,N7462,N7463,N7464,N7465,N7466,N7467,N7468,
N7469,N7470,N7471,N7472,N7473,N7474,N7475,N7476,N7477,N7478,
N7479,N7480,N7481,N7482,N7483,N7484,N7485,N7486,N7487,N7488,
N7489,N7490,N7491,N7492,N7493,N7494,N7495,N7496,N7497,N7498,
N7499,N7500,N7501,N7502,N7503,N7504,N7505,N7506,N7507,N7508,
N7509,N7510,N7511,N7512,N7513,N7514,N7515,N7516,N7517,N7518,
N7519,N7520,N7521,N7522,N7523,N7524,N7525,N7526,N7527,N7528,
N7529,N7530,N7531,N7532,N7533,N7534,N7535,N7536,N7537,N7538,
N7539,N7540,N7541,N7542,N7543,N7544,N7545,N7546,N7547,N7548,
N7549,N7550,N7551,N7552,N7553,N7554,N7555,N7556,N7557,N7558,
N7559,N7560,N7561,N7562,N7563,N7564,N7565,N7566,N7567,N7568,
N7569,N7570,N7571,N7572,N7573,N7574,N7575,N7576,N7577,N7578,
N7579,N7580,N7581,N7582,N7583,N7584,N7585,N7586,N7587,N7588,
N7589,N7590,N7591,N7592,N7593,N7594,N7595,N7596,N7597,N7598,
N7599,N7600,N7601,N7602,N7603,N7604,N7605,N7606,N7607,N7608,
N7609,N7610,N7611,N7612,N7613,N7614,N7615,N7616,N7617,N7618,
N7619,N7620,N7621,N7622,N7623,N7624,N7625,N7626,N7627,N7628,
N7629,N7630,N7631,N7632,N7633,N7634,N7635,N7636,N7637,N7638,
N7639,N7640,N7641,N7642,N7643,N7644,N7645,N7646,N7647,N7648,
N7649,N7650,N7651,N7652,N7653,N7654,N7655,N7656,N7657,N7658,
N7659,N7660,N7661,N7662,N7663,N7664,N7665,N7666,N7667,N7668,
N7669,N7670,N7671,N7672,N7673,N7674,N7675,N7676,N7677,N7678,
N7679,N7680,N7681,N7682,N7683,N7684,N7685,N7686,N7687,N7688,
N7689,N7690,N7691,N7692,N7693,N7694,N7695,N7696,N7697,N7698,
N7699,N7700,N7701,N7702,N7703,N7704,N7705,N7706,N7707,N7708,
N7709,N7710,N7711,N7712,N7713,N7714,N7715,N7716,N7717,N7718,
N7719,N7720,N7721,N7722,N7723,N7724,N7725,N7726,N7727,N7728,
N7729,N7730,N7731,N7732,N7733,N7734,N7735,N7736,N7737,N7738,
N7739,N7740,N7741,N7742,N7743,N7744,N7745,N7746,N7747,N7748,
N7749,N7750,N7751,N7752,N7753,N7754,N7755,N7756,N7757,N7758,
N7759,N7760,N7761,N7762,N7763,N7764,N7765,N7766,N7767,N7768,
N7769,N7770,N7771,N7772,N7773,N7774,N7775,N7776,N7777,N7778,
N7779,N7780,N7781,N7782,N7783,N7784,N7785,N7786,N7787,N7788,
N7789,N7790,N7791,N7792,N7793,N7794,N7795,N7796,N7797,N7798,
N7799,N7800,N7801,N7802,N7803,N7804,N7805,N7806,N7807,N7808,
N7809,N7810,N7811,N7812,N7813,N7814,N7815,N7816,N7817,N7818,
N7819,N7820,N7821,N7822,N7823,N7824,N7825,N7826,N7827,N7828,
N7829,N7830,N7831,N7832,N7833,N7834,N7835,N7836,N7837,N7838,
N7839,N7840,N7841,N7842,N7843,N7844,N7845,N7846,N7847,N7848,
N7849,N7850,N7851,N7852,N7853,N7854,N7855,N7856,N7857,N7858,
N7859,N7860,N7861,N7862,N7863,N7864,N7865,N7866,N7867,N7868,
N7869,N7870,N7871,N7872,N7873,N7874,N7875,N7876,N7877,N7878,
N7879,N7880,N7881,N7882,N7883,N7884,N7885,N7886,N7887,N7888,
N7889,N7890,N7891,N7892,N7893,N7894,N7895,N7896,N7897,N7898,
N7899,N7900,N7901,N7902,N7903,N7904,N7905,N7906,N7907,N7908,
N7909,N7910,N7911,N7912,N7913,N7914,N7915,N7916,N7917,N7918,
N7919,N7920,N7921,N7922,N7923,N7924,N7925,N7926,N7927,N7928,
N7929,N7930,N7931,N7932,N7933,N7934,N7935,N7936,N7937,N7938,
N7939,N7940,N7941,N7942,N7943,N7944,N7945,N7946,N7947,N7948,
N7949,N7950,N7951,N7952,N7953,N7954,N7955,N7956,N7957,N7958,
N7959,N7960,N7961,N7962,N7963,N7964,N7965,N7966,N7967,N7968,
N7969,N7970,N7971,N7972,N7973,N7974,N7975,N7976,N7977,N7978,
N7979,N7980,N7981,N7982,N7983,N7984,N7985,N7986,N7987,N7988,
N7989,N7990,N7991,N7992,N7993,N7994,N7995,N7996,N7997,N7998,
N7999,N8000,N8001,N8002,N8003,N8004,N8005,N8006,N8007,N8008,
N8009,N8010,N8011,N8012,N8013,N8014,N8015,N8016,N8017,N8018,
N8019,N8020,N8021,N8022,N8023,N8024,N8025,N8026,N8027,N8028,
N8029,N8030,N8031,N8032,N8033,N8034,N8035,N8036,N8037,N8038,
N8039,N8040,N8041,N8042,N8043,N8044,N8045,N8046,N8047,N8048,
N8049,N8050,N8051,N8052,N8053,N8054,N8055,N8056,N8057,N8058,
N8059,N8060,N8061,N8062,N8063,N8064,N8065,N8066,N8067,N8068,
N8069,N8070,N8071,N8072,N8073,N8074,N8075,N8076,N8077,N8078,
N8079,N8080,N8081,N8082,N8083,N8084,N8085,N8086,N8087,N8088,
N8089,N8090,N8091,N8092,N8093,N8094,N8095,N8096,N8097,N8098,
N8099,N8100,N8101,N8102,N8103,N8104,N8105,N8106,N8107,N8108,
N8109,N8110,N8111,N8112,N8113,N8114,N8115,N8116,N8117,N8118,
N8119,N8120,N8121,N8122,N8123,N8124,N8125,N8126,N8127,N8128,
N8129,N8130,N8131,N8132,N8133,N8134,N8135,N8136,N8137,N8138,
N8139,N8140,N8141,N8142,N8143,N8144,N8145,N8146,N8147,N8148,
N8149,N8150,N8151,N8152,N8153,N8154,N8155,N8156,N8157,N8158,
N8159,N8160,N8161,N8162,N8163,N8164,N8165,N8166,N8167,N8168,
N8169,N8170,N8171,N8172,N8173,N8174,N8175,N8176,N8177,N8178,
N8179,N8180,N8181,N8182,N8183,N8184,N8185,N8186,N8187,N8188,
N8189,N8190,N8191,N8192,N8193,N8194,N8195,N8196,N8197,N8198,
N8199,N8200,N8201,N8202,N8203,N8204,N8205,N8206,N8207,N8208,
N8209,N8210,N8211,N8212,N8213,N8214,N8215,N8216,N8217,N8218,
N8219,N8220,N8221,N8222,N8223,N8224,N8225,N8226,N8227,N8228,
N8229,N8230,N8231,N8232,N8233,N8234,N8235,N8236,N8237,N8238,
N8239,N8240,N8241,N8242,N8243,N8244,N8245,N8246,N8247,N8248,
N8249,N8250,N8251,N8252,N8253,N8254,N8255,N8256,N8257,N8258,
N8259,N8260,N8261,N8262,N8263,N8264,N8265,N8266,N8267,N8268,
N8269,N8270,N8271,N8272,N8273,N8274,N8275,N8276,N8277,N8278,
N8279,N8280,N8281,N8282,N8283,N8284,N8285,N8286,N8287,N8288,
N8289,N8290,N8291,N8292,N8293,N8294,N8295,N8296,N8297,N8298,
N8299,N8300,N8301,N8302,N8303,N8304,N8305,N8306,N8307,N8308,
N8309,N8310,N8311,N8312,N8313,N8314,N8315,N8316,N8317,N8318,
N8319,N8320,N8321,N8322,N8323,N8324,N8325,N8326,N8327,N8328,
N8329,N8330,N8331,N8332,N8333,N8334,N8335,N8336,N8337,N8338,
N8339,N8340,N8341,N8342,N8343,N8344,N8345,N8346,N8347,N8348,
N8349,N8350,N8351,N8352,N8353,N8354,N8355,N8356,N8357,N8358,
N8359,N8360,N8361,N8362,N8363,N8364,N8365,N8366,N8367,N8368,
N8369,N8370,N8371,N8372,N8373,N8374,N8375,N8376,N8377,N8378,
N8379,N8380,N8381,N8382,N8383,N8384,N8385,N8386,N8387,N8388,
N8389,N8390,N8391,N8392,N8393,N8394,N8395,N8396,N8397,N8398,
N8399,N8400,N8401,N8402,N8403,N8404,N8405,N8406,N8407,N8408,
N8409,N8410,N8411,N8412,N8413,N8414,N8415,N8416,N8417,N8418,
N8419,N8420,N8421,N8422,N8423,N8424,N8425,N8426,N8427,N8428,
N8429,N8430,N8431,N8432,N8433,N8434,N8435,N8436,N8437,N8438,
N8439,N8440,N8441,N8442,N8443,N8444,N8445,N8446,N8447,N8448,
N8449,N8450,N8451,N8452,N8453,N8454,N8455,N8456,N8457,N8458,
N8459,N8460,N8461,N8462,N8463,N8464,N8465,N8466,N8467,N8468,
N8469,N8470,N8471,N8472,N8473,N8474,N8475,N8476,N8477,N8478,
N8479,N8480,N8481,N8482,N8483,N8484,N8485,N8486,N8487,N8488,
N8489,N8490,N8491,N8492,N8493,N8494,N8495,N8496,N8497,N8498,
N8499,N8500,N8501,N8502,N8503,N8504,N8505,N8506,N8507,N8508,
N8509,N8510,N8511,N8512,N8513,N8514,N8515,N8516,N8517,N8518,
N8519,N8520,N8521,N8522,N8523,N8524,N8525,N8526,N8527,N8528,
N8529,N8530,N8531,N8532,N8533,N8534,N8535,N8536,N8537,N8538,
N8539,N8540,N8541,N8542,N8543,N8544,N8545,N8546,N8547,N8548,
N8549,N8550,N8551,N8552,N8553,N8554,N8555,N8556,N8557,N8558,
N8559,N8560,N8561,N8562,N8563,N8564,N8565,N8566,N8567,N8568,
N8569,N8570,N8571,N8572,N8573,N8574,N8575,N8576,N8577,N8578,
N8579,N8580,N8581,N8582,N8583,N8584,N8585,N8586,N8587,N8588,
N8589,N8590,N8591,N8592,N8593,N8594,N8595,N8596,N8597,N8598,
N8599,N8600,N8601,N8602,N8603,N8604,N8605,N8606,N8607,N8608,
N8609,N8610,N8611,N8612,N8613,N8614,N8615,N8616,N8617,N8618,
N8619,N8620,N8621,N8622,N8623,N8624,N8625,N8626,N8627,N8628,
N8629,N8630,N8631,N8632,N8633,N8634,N8635,N8636,N8637,N8638,
N8639,N8640,N8641,N8642,N8643,N8644,N8645,N8646,N8647,N8648,
N8649,N8650,N8651,N8652,N8653,N8654,N8655,N8656,N8657,N8658,
N8659,N8660,N8661,N8662,N8663,N8664,N8665,N8666,N8667,N8668,
N8669,N8670,N8671,N8672,N8673,N8674,N8675,N8676,N8677,N8678,
N8679,N8680,N8681,N8682,N8683,N8684,N8685,N8686,N8687,N8688,
N8689,N8690,N8691,N8692,N8693,N8694,N8695,N8696,N8697,N8698,
N8699,N8700,N8701,N8702,N8703,N8704,N8705,N8706,N8707,N8708,
N8709,N8710,N8711,N8712,N8713,N8714,N8715,N8716,N8717,N8718,
N8719,N8720,N8721,N8722,N8723,N8724,N8725,N8726,N8727,N8728,
N8729,N8730,N8731,N8732,N8733,N8734,N8735,N8736,N8737,N8738,
N8739,N8740,N8741,N8742,N8743,N8744,N8745,N8746,N8747,N8748,
N8749,N8750,N8751,N8752,N8753,N8754,N8755,N8756,N8757,N8758,
N8759,N8760,N8761,N8762,N8763,N8764,N8765,N8766,N8767,N8768,
N8769,N8770,N8771,N8772,N8773,N8774,N8775,N8776,N8777,N8778,
N8779,N8780,N8781,N8782,N8783,N8784,N8785,N8786,N8787,N8788,
N8789,N8790,N8791,N8792,N8793,N8794,N8795,N8796,N8797,N8798,
N8799,N8800,N8801,N8802,N8803,N8804,N8805,N8806,N8807,N8808,
N8809,N8810,N8811,N8812,N8813,N8814,N8815,N8816,N8817,N8818,
N8819,N8820,N8821,N8822,N8823,N8824,N8825,N8826,N8827,N8828,
N8829,N8830,N8831,N8832,N8833,N8834,N8835,N8836,N8837,N8838,
N8839,N8840,N8841,N8842,N8843,N8844,N8845,N8846,N8847,N8848,
N8849,N8850,N8851,N8852,N8853,N8854,N8855,N8856,N8857,N8858,
N8859,N8860,N8861,N8862,N8863,N8864,N8865,N8866,N8867,N8868,
N8869,N8870,N8871,N8872,N8873,N8874,N8875,N8876,N8877,N8878,
N8879,N8880,N8881,N8882,N8883,N8884,N8885,N8886,N8887,N8888,
N8889,N8890,N8891,N8892,N8893,N8894,N8895,N8896,N8897,N8898,
N8899,N8900,N8901,N8902,N8903,N8904,N8905,N8906,N8907,N8908,
N8909,N8910,N8911,N8912,N8913,N8914,N8915,N8916,N8917,N8918,
N8919,N8920,N8921,N8922,N8923,N8924,N8925,N8926,N8927,N8928,
N8929,N8930,N8931,N8932,N8933,N8934,N8935,N8936,N8937,N8938,
N8939,N8940,N8941,N8942,N8943,N8944,N8945,N8946,N8947,N8948,
N8949,N8950,N8951,N8952,N8953,N8954,N8955,N8956,N8957,N8958,
N8959,N8960,N8961,N8962,N8963,N8964,N8965,N8966,N8967,N8968,
N8969,N8970,N8971,N8972,N8973,N8974,N8975,N8976,N8977,N8978,
N8979,N8980,N8981,N8982,N8983,N8984,N8985,N8986,N8987,N8988,
N8989,N8990,N8991,N8992,N8993,N8994,N8995,N8996,N8997,N8998,
N8999,N9000,N9001,N9002,N9003,N9004,N9005,N9006,N9007,N9008,
N9009,N9010,N9011,N9012,N9013,N9014,N9015,N9016,N9017,N9018,
N9019,N9020,N9021,N9022,N9023,N9024,N9025,N9026,N9027,N9028,
N9029,N9030,N9031,N9032,N9033,N9034,N9035,N9036,N9037,N9038,
N9039,N9040,N9041,N9042,N9043,N9044,N9045,N9046,N9047,N9048,
N9049,N9050,N9051,N9052,N9053,N9054,N9055,N9056,N9057,N9058,
N9059,N9060,N9061,N9062,N9063,N9064,N9065,N9066,N9067,N9068,
N9069,N9070,N9071,N9072,N9073,N9074,N9075,N9076,N9077,N9078,
N9079,N9080,N9081,N9082,N9083,N9084,N9085,N9086,N9087,N9088,
N9089,N9090,N9091,N9092,N9093,N9094,N9095,N9096,N9097,N9098,
N9099,N9100,N9101,N9102,N9103,N9104,N9105,N9106,N9107,N9108,
N9109,N9110,N9111,N9112,N9113,N9114,N9115,N9116,N9117,N9118,
N9119,N9120,N9121,N9122,N9123,N9124,N9125,N9126,N9127,N9128,
N9129,N9130,N9131,N9132,N9133,N9134,N9135,N9136,N9137,N9138,
N9139,N9140,N9141,N9142,N9143,N9144,N9145,N9146,N9147,N9148,
N9149,N9150,N9151,N9152,N9153,N9154,N9155,N9156,N9157,N9158,
N9159,N9160,N9161,N9162,N9163,N9164,N9165,N9166,N9167,N9168,
N9169,N9170,N9171,N9172,N9173,N9174,N9175,N9176,N9177,N9178,
N9179,N9180,N9181,N9182,N9183,N9184,N9185,N9186,N9187,N9188,
N9189,N9190,N9191,N9192,N9193,N9194,N9195,N9196,N9197,N9198,
N9199,N9200,N9201,N9202,N9203,N9204,N9205,N9206,N9207,N9208,
N9209,N9210,N9211,N9212,N9213,N9214,N9215,N9216,N9217,N9218,
N9219,N9220,N9221,N9222,N9223,N9224,N9225,N9226,N9227,N9228,
N9229,N9230,N9231,N9232,N9233,N9234,N9235,N9236,N9237,N9238,
N9239,N9240,N9241,N9242,N9243,N9244,N9245,N9246,N9247,N9248,
N9249,N9250,N9251,N9252,N9253,N9254,N9255,N9256,N9257,N9258,
N9259,N9260,N9261,N9262,N9263,N9264,N9265,N9266,N9267,N9268,
N9269,N9270,N9271,N9272,N9273,N9274,N9275,N9276,N9277,N9278,
N9279,N9280,N9281,N9282,N9283,N9284,N9285,N9286,N9287,N9288,
N9289,N9290,N9291,N9292,N9293,N9294,N9295,N9296,N9297,N9298,
N9299,N9300,N9301,N9302,N9303,N9304,N9305,N9306,N9307,N9308,
N9309,N9310,N9311,N9312,N9313,N9314,N9315,N9316,N9317,N9318,
N9319,N9320,N9321,N9322,N9323,N9324,N9325,N9326,N9327,N9328,
N9329,N9330,N9331,N9332,N9333,N9334,N9335,N9336,N9337,N9338,
N9339,N9340,N9341,N9342,N9343,N9344,N9345,N9346,N9347,N9348,
N9349,N9350,N9351,N9352,N9353,N9354,N9355,N9356,N9357,N9358,
N9359,N9360,N9361,N9362,N9363,N9364,N9365,N9366,N9367,N9368,
N9369,N9370,N9371,N9372,N9373,N9374,N9375,N9376,N9377,N9378,
N9379,N9380,N9381,N9382,N9383,N9384,N9385,N9386,N9387,N9388,
N9389,N9390,N9391,N9392,N9393,N9394,N9395,N9396,N9397,N9398,
N9399,N9400,N9401,N9402,N9403,N9404,N9405,N9406,N9407,N9408,
N9409,N9410,N9411,N9412,N9413,N9414,N9415,N9416,N9417,N9418,
N9419,N9420,N9421,N9422,N9423,N9424,N9425,N9426,N9427,N9428,
N9429,N9430,N9431,N9432,N9433,N9434,N9435,N9436,N9437,N9438,
N9439,N9440,N9441,N9442,N9443,N9444,N9445,N9446,N9447,N9448,
N9449,N9450,N9451,N9452,N9453,N9454,N9455,N9456,N9457,N9458,
N9459,N9460,N9461,N9462,N9463,N9464,N9465,N9466,N9467,N9468,
N9469,N9470,N9471,N9472,N9473,N9474,N9475,N9476,N9477,N9478,
N9479,N9480,N9481,N9482,N9483,N9484,N9485,N9486,N9487,N9488,
N9489,N9490,N9491,N9492,N9493,N9494,N9495,N9496,N9497,N9498,
N9499,N9500,N9501,N9502,N9503,N9504,N9505,N9506,N9507,N9508,
N9509,N9510,N9511,N9512,N9513,N9514,N9515,N9516,N9517,N9518,
N9519,N9520,N9521,N9522,N9523,N9524,N9525,N9526,N9527,N9528,
N9529,N9530,N9531,N9532,N9533,N9534,N9535,N9536,N9537,N9538,
N9539,N9540,N9541,N9542,N9543,N9544,N9545,N9546,N9547,N9548,
N9549,N9550,N9551,N9552,N9553,N9554,N9555,N9556,N9557,N9558,
N9559,N9560,N9561,N9562,N9563,N9564,N9565,N9566,N9567,N9568,
N9569,N9570,N9571,N9572,N9573,N9574,N9575,N9576,N9577,N9578,
N9579,N9580,N9581,N9582,N9583,N9584,N9585,N9586,N9587,N9588,
N9589,N9590,N9591,N9592,N9593,N9594,N9595,N9596,N9597,N9598,
N9599,N9600,N9601,N9602,N9603,N9604,N9605,N9606,N9607,N9608,
N9609,N9610,N9611,N9612,N9613,N9614,N9615,N9616,N9617,N9618,
N9619,N9620,N9621,N9622,N9623,N9624,N9625,N9626,N9627,N9628,
N9629,N9630,N9631,N9632,N9633,N9634,N9635,N9636,N9637,N9638,
N9639,N9640,N9641,N9642,N9643,N9644,N9645,N9646,N9647,N9648,
N9649,N9650,N9651,N9652,N9653,N9654,N9655,N9656,N9657,N9658,
N9659,N9660,N9661,N9662,N9663,N9664,N9665,N9666,N9667,N9668,
N9669,N9670,N9671,N9672,N9673,N9674,N9675,N9676,N9677,N9678,
N9679,N9680,N9681,N9682,N9683,N9684,N9685,N9686,N9687,N9688,
N9689,N9690,N9691,N9692,N9693,N9694,N9695,N9696,N9697,N9698,
N9699,N9700,N9701,N9702,N9703,N9704,N9705,N9706,N9707,N9708,
N9709,N9710,N9711,N9712,N9713,N9714,N9715,N9716,N9717,N9718,
N9719,N9720,N9721,N9722,N9723,N9724,N9725,N9726,N9727,N9728,
N9729,N9730,N9731,N9732,N9733,N9734,N9735,N9736,N9737,N9738,
N9739,N9740,N9741,N9742,N9743,N9744,N9745,N9746,N9747,N9748,
N9749,N9750,N9751,N9752,N9753,N9754,N9755,N9756,N9757,N9758,
N9759,N9760,N9761,N9762,N9763,N9764,N9765,N9766,N9767,N9768,
N9769,N9770,N9771,N9772,N9773,N9774,N9775,N9776,N9777,N9778,
N9779,N9780,N9781,N9782,N9783,N9784,N9785,N9786,N9787,N9788,
N9789,N9790,N9791,N9792,N9793,N9794,N9795,N9796,N9797,N9798,
N9799,N9800,N9801,N9802,N9803,N9804,N9805,N9806,N9807,N9808,
N9809,N9810,N9811,N9812,N9813,N9814,N9815,N9816,N9817,N9818,
N9819,N9820,N9821,N9822,N9823,N9824,N9825,N9826,N9827,N9828,
N9829,N9830,N9831,N9832,N9833,N9834,N9835,N9836,N9837,N9838,
N9839,N9840,N9841,N9842,N9843,N9844,N9845,N9846,N9847,N9848,
N9849,N9850,N9851,N9852,N9853,N9854,N9855,N9856,N9857,N9858,
N9859,N9860,N9861,N9862,N9863,N9864,N9865,N9866,N9867,N9868,
N9869,N9870,N9871,N9872,N9873,N9874,N9875,N9876,N9877,N9878,
N9879,N9880,N9881,N9882,N9883,N9884,N9885,N9886,N9887,N9888,
N9889,N9890,N9891,N9892,N9893,N9894,N9895,N9896,N9897,N9898,
N9899,N9900,N9901,N9902,N9903,N9904,N9905,N9906,N9907,N9908,
N9909,N9910,N9911,N9912,N9913,N9914,N9915,N9916,N9917,N9918,
N9919,N9920,N9921,N9922,N9923,N9924,N9925,N9926,N9927,N9928,
N9929,N9930,N9931,N9932,N9933,N9934,N9935,N9936,N9937,N9938,
N9939,N9940,N9941,N9942,N9943,N9944,N9945,N9946,N9947,N9948,
N9949,N9950,N9951,N9952,N9953,N9954,N9955,N9956,N9957,N9958,
N9959,N9960,N9961,N9962,N9963,N9964,N9965,N9966,N9967,N9968,
N9969,N9970,N9971,N9972,N9973,N9974,N9975,N9976,N9977,N9978,
N9979,N9980,N9981,N9982,N9983,N9984,N9985,N9986,N9987,N9988,
N9989,N9990,N9991,N9992,N9993,N9994,N9995,N9996,N9997,N9998,
N9999,N10000,N10001,N10002,N10003,N10004,N10005,N10006,N10007,N10008,
N10009,N10010,N10011,N10012,N10013,N10014,N10015,N10016,N10017,N10018,
N10019,N10020,N10021,N10022,N10023,N10024,N10025,N10026,N10027,N10028,
N10029,N10030,N10031,N10032,N10033,N10034,N10035,N10036,N10037,N10038,
N10039,N10040,N10041,N10042,N10043,N10044,N10045,N10046,N10047,N10048,
N10049,N10050,N10051,N10052,N10053,N10054,N10055,N10056,N10057,N10058,
N10059,N10060,N10061,N10062,N10063,N10064,N10065,N10066,N10067,N10068,
N10069,N10070,N10071,N10072,N10073,N10074,N10075,N10076,N10077,N10078,
N10079,N10080,N10081,N10082,N10083,N10084,N10085,N10086,N10087,N10088,
N10089,N10090,N10091,N10092,N10093,N10094,N10095,N10096,N10097,N10098,
N10099,N10100,N10101,N10102,N10103,N10104,N10105,N10106,N10107,N10108,
N10109,N10110,N10111,N10112,N10113,N10114,N10115,N10116,N10117,N10118,
N10119,N10120,N10121,N10122,N10123,N10124,N10125,N10126,N10127,N10128,
N10129,N10130,N10131,N10132,N10133,N10134,N10135,N10136,N10137,N10138,
N10139,N10140,N10141,N10142,N10143,N10144,N10145,N10146,N10147,N10148,
N10149,N10150,N10151,N10152,N10153,N10154,N10155,N10156,N10157,N10158,
N10159,N10160,N10161,N10162,N10163,N10164,N10165,N10166,N10167,N10168,
N10169,N10170,N10171,N10172,N10173,N10174,N10175,N10176,N10177,N10178,
N10179,N10180,N10181,N10182,N10183,N10184,N10185,N10186,N10187,N10188,
N10189,N10190,N10191,N10192,N10193,N10194,N10195,N10196,N10197,N10198,
N10199,N10200,N10201,N10202,N10203,N10204,N10205,N10206,N10207,N10208,
N10209,N10210,N10211,N10212,N10213,N10214,N10215,N10216,N10217,N10218,
N10219,N10220,N10221,N10222,N10223,N10224,N10225,N10226,N10227,N10228,
N10229,N10230,N10231,N10232,N10233,N10234,N10235,N10236,N10237,N10238,
N10239,N10240,N10241,N10242,N10243,N10244,N10245,N10246,N10247,N10248,
N10249,N10250,N10251,N10252,N10253,N10254,N10255,N10256,N10257,N10258,
N10259,N10260,N10261,N10262,N10263,N10264,N10265,N10266,N10267,N10268,
N10269,N10270,N10271,N10272,N10273,N10274,N10275,N10276,N10277,N10278,
N10279,N10280,N10281,N10282,N10283,N10284,N10285,N10286,N10287,N10288,
N10289,N10290,N10291,N10292,N10293,N10294,N10295,N10296,N10297,N10298,
N10299,N10300,N10301,N10302,N10303,N10304,N10305,N10306,N10307,N10308,
N10309,N10310,N10311,N10312,N10313,N10314,N10315,N10316,N10317,N10318,
N10319,N10320,N10321,N10322,N10323,N10324,N10325,N10326,N10327,N10328,
N10329,N10330,N10331,N10332,N10333,N10334,N10335,N10336,N10337,N10338,
N10339,N10340,N10341,N10342,N10343,N10344,N10345,N10346,N10347,N10348,
N10349,N10350,N10351,N10352,N10353,N10354,N10355,N10356,N10357,N10358,
N10359,N10360,N10361,N10362,N10363,N10364,N10365,N10366,N10367,N10368,
N10369,N10370,N10371,N10372,N10373,N10374,N10375,N10376,N10377,N10378,
N10379,N10380,N10381,N10382,N10383,N10384,N10385,N10386,N10387,N10388,
N10389,N10390,N10391,N10392,N10393,N10394,N10395,N10396,N10397,N10398,
N10399,N10400,N10401,N10402,N10403,N10404,N10405,N10406,N10407,N10408,
N10409,N10410,N10411,N10412,N10413,N10414,N10415,N10416,N10417,N10418,
N10419,N10420,N10421,N10422,N10423,N10424,N10425,N10426,N10427,N10428,
N10429,N10430,N10431,N10432,N10433,N10434,N10435,N10436,N10437,N10438,
N10439,N10440,N10441,N10442,N10443,N10444,N10445,N10446,N10447,N10448,
N10449,N10450,N10451,N10452,N10453,N10454,N10455,N10456,N10457,N10458,
N10459,N10460,N10461,N10462,N10463,N10464,N10465,N10466,N10467,N10468,
N10469,N10470,N10471,N10472,N10473,N10474,N10475,N10476,N10477,N10478,
N10479,N10480,N10481,N10482,N10483,N10484,N10485,N10486,N10487,N10488,
N10489,N10490,N10491,N10492,N10493,N10494,N10495,N10496,N10497,N10498,
N10499,N10500,N10501,N10502,N10503,N10504,N10505,N10506,N10507,N10508,
N10509,N10510,N10511,N10512,N10513,N10514,N10515,N10516,N10517,N10518,
N10519,N10520,N10521,N10522,N10523,N10524,N10525,N10526,N10527,N10528,
N10529,N10530,N10531,N10532,N10533,N10534,N10535,N10536,N10537,N10538,
N10539,N10540,N10541,N10542,N10543,N10544,N10545,N10546,N10547,N10548,
N10549,N10550,N10551,N10552,N10553,N10554,N10555,N10556,N10557,N10558,
N10559,N10560,N10561,N10562,N10563,N10564,N10565,N10566,N10567,N10568,
N10569,N10570,N10571,N10572,N10573,N10574,N10575,N10576,N10577,N10578,
N10579,N10580,N10581,N10582,N10583,N10584,N10585,N10586,N10587,N10588,
N10589,N10590,N10591,N10592,N10593,N10594,N10595,N10596,N10597,N10598,
N10599,N10600,N10601,N10602,N10603,N10604,N10605,N10606,N10607,N10608,
N10609,N10610,N10611,N10612,N10613,N10614,N10615,N10616,N10617,N10618,
N10619,N10620,N10621,N10622,N10623,N10624,N10625,N10626,N10627,N10628,
N10629,N10630,N10631,N10632,N10633,N10634,N10635,N10636,N10637,N10638,
N10639,N10640,N10641,N10642,N10643,N10644,N10645,N10646,N10647,N10648,
N10649,N10650,N10651,N10652,N10653,N10654,N10655,N10656,N10657,N10658,
N10659,N10660,N10661,N10662,N10663,N10664,N10665,N10666,N10667,N10668,
N10669,N10670,N10671,N10672,N10673,N10674,N10675,N10676,N10677,N10678,
N10679,N10680,N10681,N10682,N10683,N10684,N10685,N10686,N10687,N10688,
N10689,N10690,N10691,N10692,N10693,N10694,N10695,N10696,N10697,N10698,
N10699,N10700,N10701,N10702,N10703,N10704,N10705,N10706,N10707,N10708,
N10709,N10710,N10711,N10712,N10713,N10714,N10715,N10716,N10717,N10718,
N10719,N10720,N10721,N10722,N10723,N10724,N10725,N10726,N10727,N10728,
N10729,N10730,N10731,N10732,N10733,N10734,N10735,N10736,N10737,N10738,
N10739,N10740,N10741,N10742,N10743,N10744,N10745,N10746,N10747,N10748,
N10749,N10750,N10751,N10752,N10753,N10754,N10755,N10756,N10757,N10758,
N10759,N10760,N10761,N10762,N10763,N10764,N10765,N10766,N10767,N10768,
N10769,N10770,N10771,N10772,N10773,N10774,N10775,N10776,N10777,N10778,
N10779,N10780,N10781,N10782,N10783,N10784,N10785,N10786,N10787,N10788,
N10789,N10790,N10791,N10792,N10793,N10794,N10795,N10796,N10797,N10798,
N10799,N10800,N10801,N10802,N10803,N10804,N10805,N10806,N10807,N10808,
N10809,N10810,N10811,N10812,N10813,N10814,N10815,N10816,N10817,N10818,
N10819,N10820,N10821,N10822,N10823,N10824,N10825,N10826,N10827,N10828,
N10829,N10830,N10831,N10832,N10833,N10834,N10835,N10836,N10837,N10838,
N10839,N10840,N10841,N10842,N10843,N10844,N10845,N10846,N10847,N10848,
N10849,N10850,N10851,N10852,N10853,N10854,N10855,N10856,N10857,N10858,
N10859,N10860,N10861,N10862,N10863,N10864,N10865,N10866,N10867,N10868,
N10869,N10870,N10871,N10872,N10873,N10874,N10875,N10876,N10877,N10878,
N10879,N10880,N10881,N10882,N10883,N10884,N10885,N10886,N10887,N10888,
N10889,N10890,N10891,N10892,N10893,N10894,N10895,N10896,N10897,N10898,
N10899,N10900,N10901,N10902,N10903,N10904,N10905,N10906,N10907,N10908,
N10909,N10910,N10911,N10912,N10913,N10914,N10915,N10916,N10917,N10918,
N10919,N10920,N10921,N10922,N10923,N10924,N10925,N10926,N10927,N10928,
N10929,N10930,N10931,N10932,N10933,N10934,N10935,N10936,N10937,N10938,
N10939,N10940,N10941,N10942,N10943,N10944,N10945,N10946,N10947,N10948,
N10949,N10950,N10951,N10952,N10953,N10954,N10955,N10956,N10957,N10958,
N10959,N10960,N10961,N10962,N10963,N10964,N10965,N10966,N10967,N10968,
N10969,N10970,N10971,N10972,N10973,N10974,N10975,N10976,N10977,N10978,
N10979,N10980,N10981,N10982,N10983,N10984,N10985,N10986,N10987,N10988,
N10989,N10990,N10991,N10992,N10993,N10994,N10995,N10996,N10997,N10998,
N10999,N11000,N11001,N11002,N11003,N11004,N11005,N11006,N11007,N11008,
N11009,N11010,N11011,N11012,N11013,N11014,N11015,N11016,N11017,N11018,
N11019,N11020,N11021,N11022,N11023,N11024,N11025,N11026,N11027,N11028,
N11029,N11030,N11031,N11032,N11033,N11034,N11035,N11036,N11037,N11038,
N11039,N11040,N11041,N11042,N11043,N11044,N11045,N11046,N11047,N11048,
N11049,N11050,N11051,N11052,N11053,N11054,N11055,N11056,N11057,N11058,
N11059,N11060,N11061,N11062,N11063,N11064,N11065,N11066,N11067,N11068,
N11069,N11070,N11071,N11072,N11073,N11074,N11075,N11076,N11077,N11078,
N11079,N11080,N11081,N11082,N11083,N11084,N11085,N11086,N11087,N11088,
N11089,N11090,N11091,N11092,N11093,N11094,N11095,N11096,N11097,N11098,
N11099,N11100,N11101,N11102,N11103,N11104,N11105,N11106,N11107,N11108,
N11109,N11110,N11111,N11112,N11113,N11114,N11115,N11116,N11117,N11118,
N11119,N11120,N11121,N11122,N11123,N11124,N11125,N11126,N11127,N11128,
N11129,N11130,N11131,N11132,N11133,N11134,N11135,N11136,N11137,N11138,
N11139,N11140,N11141,N11142,N11143,N11144,N11145,N11146,N11147,N11148,
N11149,N11150,N11151,N11152,N11153,N11154,N11155,N11156,N11157,N11158,
N11159,N11160,N11161,N11162,N11163,N11164,N11165,N11166,N11167,N11168,
N11169,N11170,N11171,N11172,N11173,N11174,N11175,N11176,N11177,N11178,
N11179,N11180,N11181,N11182,N11183,N11184,N11185,N11186,N11187,N11188,
N11189,N11190,N11191,N11192,N11193,N11194,N11195,N11196,N11197,N11198,
N11199,N11200,N11201,N11202,N11203,N11204,N11205,N11206,N11207,N11208,
N11209,N11210,N11211,N11212,N11213,N11214,N11215,N11216,N11217,N11218,
N11219,N11220,N11221,N11222,N11223,N11224,N11225,N11226,N11227,N11228,
N11229,N11230,N11231,N11232,N11233,N11234,N11235,N11236,N11237,N11238,
N11239,N11240,N11241,N11242,N11243,N11244,N11245,N11246,N11247,N11248,
N11249,N11250,N11251,N11252,N11253,N11254,N11255,N11256,N11257,N11258,
N11259,N11260,N11261,N11262,N11263,N11264,N11265,N11266,N11267,N11268,
N11269,N11270,N11271,N11272,N11273,N11274,N11275,N11276,N11277,N11278,
N11279,N11280,N11281,N11282,N11283,N11284,N11285,N11286,N11287,N11288,
N11289,N11290,N11291,N11292,N11293,N11294,N11295,N11296,N11297,N11298,
N11299,N11300,N11301,N11302,N11303,N11304,N11305,N11306,N11307,N11308,
N11309,N11310,N11311,N11312,N11313,N11314,N11315,N11316,N11317,N11318,
N11319,N11320,N11321,N11322,N11323,N11324,N11325,N11326,N11327,N11328,
N11329,N11330,N11331,N11332,N11333,N11334,N11335,N11336,N11337,N11338,
N11339,N11340,N11341,N11342,N11343,N11344,N11345,N11346,N11347,N11348,
N11349,N11350,N11351,N11352,N11353,N11354,N11355,N11356,N11357,N11358,
N11359,N11360,N11361,N11362,N11363,N11364,N11365,N11366,N11367,N11368,
N11369,N11370,N11371,N11372,N11373,N11374,N11375,N11376,N11377,N11378,
N11379,N11380,N11381,N11382,N11383,N11384,N11385,N11386,N11387,N11388,
N11389,N11390,N11391,N11392,N11393,N11394,N11395,N11396,N11397,N11398,
N11399,N11400,N11401,N11402,N11403,N11404,N11405,N11406,N11407,N11408,
N11409,N11410,N11411,N11412,N11413,N11414,N11415,N11416,N11417,N11418,
N11419,N11420,N11421,N11422,N11423,N11424,N11425,N11426,N11427,N11428,
N11429,N11430,N11431,N11432,N11433,N11434,N11435,N11436,N11437,N11438,
N11439,N11440,N11441,N11442,N11443,N11444,N11445,N11446,N11447,N11448,
N11449,N11450,N11451,N11452,N11453,N11454,N11455,N11456,N11457,N11458,
N11459,N11460,N11461,N11462,N11463,N11464,N11465,N11466,N11467,N11468,
N11469,N11470,N11471,N11472,N11473,N11474,N11475,N11476,N11477,N11478,
N11479,N11480,N11481,N11482,N11483,N11484,N11485,N11486,N11487,N11488,
N11489,N11490,N11491,N11492,N11493,N11494,N11495,N11496,N11497,N11498,
N11499,N11500,N11501,N11502,N11503,N11504,N11505,N11506,N11507,N11508,
N11509,N11510,N11511,N11512,N11513,N11514,N11515,N11516,N11517,N11518,
N11519,N11520,N11521,N11522,N11523,N11524,N11525,N11526,N11527,N11528,
N11529,N11530,N11531,N11532,N11533,N11534,N11535,N11536,N11537,N11538,
N11539,N11540,N11541,N11542,N11543,N11544,N11545,N11546,N11547,N11548,
N11549,N11550,N11551,N11552,N11553,N11554,N11555,N11556,N11557,N11558,
N11559,N11560,N11561,N11562,N11563,N11564,N11565,N11566,N11567,N11568,
N11569,N11570,N11571,N11572,N11573,N11574,N11575,N11576,N11577,N11578,
N11579,N11580,N11581,N11582,N11583,N11584,N11585,N11586,N11587,N11588,
N11589,N11590,N11591,N11592,N11593,N11594,N11595,N11596,N11597,N11598,
N11599,N11600,N11601,N11602,N11603,N11604,N11605,N11606,N11607,N11608,
N11609,N11610,N11611,N11612,N11613,N11614,N11615,N11616,N11617,N11618,
N11619,N11620,N11621,N11622,N11623,N11624,N11625,N11626,N11627,N11628,
N11629,N11630,N11631,N11632,N11633,N11634,N11635,N11636,N11637,N11638,
N11639,N11640,N11641,N11642,N11643,N11644,N11645,N11646,N11647,N11648,
N11649,N11650,N11651,N11652,N11653,N11654,N11655,N11656,N11657,N11658,
N11659,N11660,N11661,N11662,N11663,N11664,N11665,N11666,N11667,N11668,
N11669,N11670,N11671,N11672,N11673,N11674,N11675,N11676,N11677,N11678,
N11679,N11680,N11681,N11682,N11683,N11684,N11685,N11686,N11687,N11688,
N11689,N11690,N11691,N11692,N11693,N11694,N11695,N11696,N11697,N11698,
N11699,N11700,N11701,N11702,N11703,N11704,N11705,N11706,N11707,N11708,
N11709,N11710,N11711,N11712,N11713,N11714,N11715,N11716,N11717,N11718,
N11719,N11720,N11721,N11722,N11723,N11724,N11725,N11726,N11727,N11728,
N11729,N11730,N11731,N11732,N11733,N11734,N11735,N11736,N11737,N11738,
N11739,N11740,N11741,N11742,N11743,N11744,N11745,N11746,N11747,N11748,
N11749,N11750,N11751,N11752,N11753,N11754,N11755,N11756,N11757,N11758,
N11759,N11760,N11761,N11762,N11763,N11764,N11765,N11766,N11767,N11768,
N11769,N11770,N11771,N11772,N11773,N11774,N11775,N11776,N11777,N11778,
N11779,N11780,N11781,N11782,N11783,N11784,N11785,N11786,N11787,N11788,
N11789,N11790,N11791,N11792,N11793,N11794,N11795,N11796,N11797,N11798,
N11799,N11800,N11801,N11802,N11803,N11804,N11805,N11806,N11807,N11808,
N11809,N11810,N11811,N11812,N11813,N11814,N11815,N11816,N11817,N11818,
N11819,N11820,N11821,N11822,N11823,N11824,N11825,N11826,N11827,N11828,
N11829,N11830,N11831,N11832,N11833,N11834,N11835,N11836,N11837,N11838,
N11839,N11840,N11841,N11842,N11843,N11844,N11845,N11846,N11847,N11848,
N11849,N11850,N11851,N11852,N11853,N11854,N11855,N11856,N11857,N11858,
N11859,N11860,N11861,N11862,N11863,N11864,N11865,N11866,N11867,N11868,
N11869,N11870,N11871,N11872,N11873,N11874,N11875,N11876,N11877,N11878,
N11879,N11880,N11881,N11882,N11883,N11884,N11885,N11886,N11887,N11888,
N11889,N11890,N11891,N11892,N11893,N11894,N11895,N11896,N11897,N11898,
N11899,N11900,N11901,N11902,N11903,N11904,N11905,N11906,N11907,N11908,
N11909,N11910,N11911,N11912,N11913,N11914,N11915,N11916,N11917,N11918,
N11919,N11920,N11921,N11922,N11923,N11924,N11925,N11926,N11927,N11928,
N11929,N11930,N11931,N11932,N11933,N11934,N11935,N11936,N11937,N11938,
N11939,N11940,N11941,N11942,N11943,N11944,N11945,N11946,N11947,N11948,
N11949,N11950,N11951,N11952,N11953,N11954,N11955,N11956,N11957,N11958,
N11959,N11960,N11961,N11962,N11963,N11964,N11965,N11966,N11967,N11968,
N11969,N11970,N11971,N11972,N11973,N11974,N11975,N11976,N11977,N11978,
N11979,N11980,N11981,N11982,N11983,N11984,N11985,N11986,N11987,N11988,
N11989,N11990,N11991,N11992,N11993,N11994,N11995,N11996,N11997,N11998,
N11999,N12000,N12001,N12002,N12003,N12004,N12005,N12006,N12007,N12008,
N12009,N12010,N12011,N12012,N12013,N12014,N12015,N12016,N12017,N12018,
N12019,N12020,N12021,N12022,N12023,N12024,N12025,N12026,N12027,N12028,
N12029,N12030,N12031,N12032,N12033,N12034,N12035,N12036,N12037,N12038,
N12039,N12040,N12041,N12042,N12043,N12044,N12045,N12046,N12047,N12048,
N12049,N12050,N12051,N12052,N12053,N12054,N12055,N12056,N12057,N12058,
N12059,N12060,N12061,N12062,N12063,N12064,N12065,N12066,N12067,N12068,
N12069,N12070,N12071,N12072,N12073,N12074,N12075,N12076,N12077,N12078,
N12079,N12080,N12081,N12082,N12083,N12084,N12085,N12086,N12087,N12088,
N12089,N12090,N12091,N12092,N12093,N12094,N12095,N12096,N12097,N12098,
N12099,N12100,N12101,N12102,N12103,N12104,N12105,N12106,N12107,N12108,
N12109,N12110,N12111,N12112,N12113,N12114,N12115,N12116,N12117,N12118,
N12119,N12120,N12121,N12122,N12123,N12124,N12125,N12126,N12127,N12128,
N12129,N12130,N12131,N12132,N12133,N12134,N12135,N12136,N12137,N12138,
N12139,N12140,N12141,N12142,N12143,N12144,N12145,N12146,N12147,N12148,
N12149,N12150,N12151,N12152,N12153,N12154,N12155,N12156,N12157,N12158,
N12159,N12160,N12161,N12162,N12163,N12164,N12165,N12166,N12167,N12168,
N12169,N12170,N12171,N12172,N12173,N12174,N12175,N12176,N12177,N12178,
N12179,N12180,N12181,N12182,N12183,N12184,N12185,N12186,N12187,N12188,
N12189,N12190,N12191,N12192,N12193,N12194,N12195,N12196,N12197,N12198,
N12199,N12200,N12201,N12202,N12203,N12204,N12205,N12206,N12207,N12208,
N12209,N12210,N12211,N12212,N12213,N12214,N12215,N12216,N12217,N12218,
N12219,N12220,N12221,N12222,N12223,N12224,N12225,N12226,N12227,N12228,
N12229,N12230,N12231,N12232,N12233,N12234,N12235,N12236,N12237,N12238,
N12239,N12240,N12241,N12242,N12243,N12244,N12245,N12246,N12247,N12248,
N12249,N12250,N12251,N12252,N12253,N12254,N12255,N12256,N12257,N12258,
N12259,N12260,N12261,N12262,N12263,N12264,N12265,N12266,N12267,N12268,
N12269,N12270,N12271,N12272,N12273,N12274,N12275,N12276,N12277,N12278,
N12279,N12280,N12281,N12282,N12283,N12284,N12285,N12286,N12287,N12288,
N12289,N12290,N12291,N12292,N12293,N12294,N12295,N12296,N12297,N12298,
N12299,N12300,N12301,N12302,N12303,N12304,N12305,N12306,N12307,N12308,
N12309,N12310,N12311,N12312,N12313,N12314,N12315,N12316,N12317,N12318,
N12319,N12320,N12321,N12322,N12323,N12324,N12325,N12326,N12327,N12328,
N12329,N12330,N12331,N12332,N12333,N12334,N12335,N12336,N12337,N12338,
N12339,N12340,N12341,N12342,N12343,N12344,N12345,N12346,N12347,N12348,
N12349,N12350,N12351,N12352,N12353,N12354,N12355,N12356,N12357,N12358,
N12359,N12360,N12361,N12362,N12363,N12364,N12365,N12366,N12367,N12368,
N12369,N12370,N12371,N12372,N12373,N12374,N12375,N12376,N12377,N12378,
N12379,N12380,N12381,N12382,N12383,N12384,N12385,N12386,N12387,N12388,
N12389,N12390,N12391,N12392,N12393,N12394,N12395,N12396,N12397,N12398,
N12399,N12400,N12401,N12402,N12403,N12404,N12405,N12406,N12407,N12408,
N12409,N12410,N12411,N12412,N12413,N12414,N12415,N12416,N12417,N12418,
N12419,N12420,N12421,N12422,N12423,N12424,N12425,N12426,N12427,N12428,
N12429,N12430,N12431,N12432,N12433,N12434,N12435,N12436,N12437,N12438,
N12439,N12440,N12441,N12442,N12443,N12444,N12445,N12446,N12447,N12448,
N12449,N12450,N12451,N12452,N12453,N12454,N12455,N12456,N12457,N12458,
N12459,N12460,N12461,N12462,N12463,N12464,N12465,N12466,N12467,N12468,
N12469,N12470,N12471,N12472,N12473,N12474,N12475,N12476,N12477,N12478,
N12479,N12480,N12481,N12482,N12483,N12484,N12485,N12486,N12487,N12488,
N12489,N12490,N12491,N12492,N12493,N12494,N12495,N12496,N12497,N12498,
N12499,N12500,N12501,N12502,N12503,N12504,N12505,N12506,N12507,N12508,
N12509,N12510,N12511,N12512,N12513,N12514,N12515,N12516,N12517,N12518,
N12519,N12520,N12521,N12522,N12523,N12524,N12525,N12526,N12527,N12528,
N12529,N12530,N12531,N12532,N12533,N12534,N12535,N12536,N12537,N12538,
N12539,N12540,N12541,N12542,N12543,N12544,N12545,N12546,N12547,N12548,
N12549,N12550,N12551,N12552,N12553,N12554,N12555,N12556,N12557,N12558,
N12559,N12560,N12561,N12562,N12563,N12564,N12565,N12566,N12567,N12568,
N12569,N12570,N12571,N12572,N12573,N12574,N12575,N12576,N12577,N12578,
N12579,N12580,N12581,N12582,N12583,N12584,N12585,N12586,N12587,N12588,
N12589,N12590,N12591,N12592,N12593,N12594,N12595,N12596,N12597,N12598,
N12599,N12600,N12601,N12602,N12603,N12604,N12605,N12606,N12607,N12608,
N12609,N12610,N12611,N12612,N12613,N12614,N12615,N12616,N12617,N12618,
N12619,N12620,N12621,N12622,N12623,N12624,N12625,N12626,N12627,N12628,
N12629,N12630,N12631,N12632,N12633,N12634,N12635,N12636,N12637,N12638,
N12639,N12640,N12641,N12642,N12643,N12644,N12645,N12646,N12647,N12648,
N12649,N12650,N12651,N12652,N12653,N12654,N12655,N12656,N12657,N12658,
N12659,N12660,N12661,N12662,N12663,N12664,N12665,N12666,N12667,N12668,
N12669,N12670,N12671,N12672,N12673,N12674,N12675,N12676,N12677,N12678,
N12679,N12680,N12681,N12682,N12683,N12684,N12685,N12686,N12687,N12688,
N12689,N12690,N12691,N12692,N12693,N12694,N12695,N12696,N12697,N12698,
N12699,N12700,N12701,N12702,N12703,N12704,N12705,N12706,N12707,N12708,
N12709,N12710,N12711,N12712,N12713,N12714,N12715,N12716,N12717,N12718,
N12719,N12720,N12721,N12722,N12723,N12724,N12725,N12726,N12727,N12728,
N12729,N12730,N12731,N12732,N12733,N12734,N12735,N12736,N12737,N12738,
N12739,N12740,N12741,N12742,N12743,N12744,N12745,N12746,N12747,N12748,
N12749,N12750,N12751,N12752,N12753,N12754,N12755,N12756,N12757,N12758,
N12759,N12760,N12761,N12762,N12763,N12764,N12765,N12766,N12767,N12768,
N12769,N12770,N12771,N12772,N12773,N12774,N12775,N12776,N12777,N12778,
N12779,N12780,N12781,N12782,N12783,N12784,N12785,N12786,N12787,N12788,
N12789,N12790,N12791,N12792,N12793,N12794,N12795,N12796,N12797,N12798,
N12799,N12800,N12801,N12802,N12803,N12804,N12805,N12806,N12807,N12808,
N12809,N12810,N12811,N12812,N12813,N12814,N12815,N12816,N12817,N12818,
N12819,N12820,N12821,N12822,N12823,N12824,N12825,N12826,N12827,N12828,
N12829,N12830,N12831,N12832,N12833,N12834,N12835,N12836,N12837,N12838,
N12839,N12840,N12841,N12842,N12843,N12844,N12845,N12846,N12847,N12848,
N12849,N12850,N12851,N12852,N12853,N12854,N12855,N12856,N12857,N12858,
N12859,N12860,N12861,N12862,N12863,N12864,N12865,N12866,N12867,N12868,
N12869,N12870,N12871,N12872,N12873,N12874,N12875,N12876,N12877,N12878,
N12879,N12880,N12881,N12882,N12883,N12884,N12885,N12886,N12887,N12888,
N12889,N12890,N12891,N12892,N12893,N12894,N12895,N12896,N12897,N12898,
N12899,N12900,N12901,N12902,N12903,N12904,N12905,N12906,N12907,N12908,
N12909,N12910,N12911,N12912,N12913,N12914,N12915,N12916,N12917,N12918,
N12919,N12920,N12921,N12922,N12923,N12924,N12925,N12926,N12927,N12928,
N12929,N12930,N12931,N12932,N12933,N12934,N12935,N12936,N12937,N12938,
N12939,N12940,N12941,N12942,N12943,N12944,N12945,N12946,N12947,N12948,
N12949,N12950,N12951,N12952,N12953,N12954,N12955,N12956,N12957,N12958,
N12959,N12960,N12961,N12962,N12963,N12964,N12965,N12966,N12967,N12968,
N12969,N12970,N12971,N12972,N12973,N12974,N12975,N12976,N12977,N12978,
N12979,N12980,N12981,N12982,N12983,N12984,N12985,N12986,N12987,N12988,
N12989,N12990,N12991,N12992,N12993,N12994,N12995,N12996,N12997,N12998,
N12999,N13000,N13001,N13002,N13003,N13004,N13005,N13006,N13007,N13008,
N13009,N13010,N13011,N13012,N13013,N13014,N13015,N13016,N13017,N13018,
N13019,N13020,N13021,N13022,N13023,N13024,N13025,N13026,N13027,N13028,
N13029,N13030,N13031,N13032,N13033,N13034,N13035,N13036,N13037,N13038,
N13039,N13040,N13041,N13042,N13043,N13044,N13045,N13046,N13047,N13048,
N13049,N13050,N13051,N13052,N13053,N13054,N13055,N13056,N13057,N13058,
N13059,N13060,N13061,N13062,N13063,N13064,N13065,N13066,N13067,N13068,
N13069,N13070,N13071,N13072,N13073,N13074,N13075,N13076,N13077,N13078,
N13079,N13080,N13081,N13082,N13083,N13084,N13085,N13086,N13087,N13088,
N13089,N13090,N13091,N13092,N13093,N13094,N13095,N13096,N13097,N13098,
N13099,N13100,N13101,N13102,N13103,N13104,N13105,N13106,N13107,N13108,
N13109,N13110,N13111,N13112,N13113,N13114,N13115,N13116,N13117,N13118,
N13119,N13120,N13121,N13122,N13123,N13124,N13125,N13126,N13127,N13128,
N13129,N13130,N13131,N13132,N13133,N13134,N13135,N13136,N13137,N13138,
N13139,N13140,N13141,N13142,N13143,N13144,N13145,N13146,N13147,N13148,
N13149,N13150,N13151,N13152,N13153,N13154,N13155,N13156,N13157,N13158,
N13159,N13160,N13161,N13162,N13163,N13164,N13165,N13166,N13167,N13168,
N13169,N13170,N13171,N13172,N13173,N13174,N13175,N13176,N13177,N13178,
N13179,N13180,N13181,N13182,N13183,N13184,N13185,N13186,N13187,N13188,
N13189,N13190,N13191,N13192,N13193,N13194,N13195,N13196,N13197,N13198,
N13199,N13200,N13201,N13202,N13203,N13204,N13205,N13206,N13207,N13208,
N13209,N13210,N13211,N13212,N13213,N13214,N13215,N13216,N13217,N13218,
N13219,N13220,N13221,N13222,N13223,N13224,N13225,N13226,N13227,N13228,
N13229,N13230,N13231,N13232,N13233,N13234,N13235,N13236,N13237,N13238,
N13239,N13240,N13241,N13242,N13243,N13244,N13245,N13246,N13247,N13248,
N13249,N13250,N13251,N13252,N13253,N13254,N13255,N13256,N13257,N13258,
N13259,N13260,N13261,N13262,N13263,N13264,N13265,N13266,N13267,N13268,
N13269,N13270,N13271,N13272,N13273,N13274,N13275,N13276,N13277,N13278,
N13279,N13280,N13281,N13282,N13283,N13284,N13285,N13286,N13287,N13288,
N13289,N13290,N13291,N13292,N13293,N13294,N13295,N13296,N13297,N13298,
N13299,N13300,N13301,N13302,N13303,N13304,N13305,N13306,N13307,N13308,
N13309,N13310,N13311,N13312,N13313,N13314,N13315,N13316,N13317,N13318,
N13319,N13320,N13321,N13322,N13323,N13324,N13325,N13326,N13327,N13328,
N13329,N13330,N13331,N13332,N13333,N13334,N13335,N13336,N13337,N13338,
N13339,N13340,N13341,N13342,N13343,N13344,N13345,N13346,N13347,N13348,
N13349,N13350,N13351,N13352,N13353,N13354,N13355,N13356,N13357,N13358,
N13359,N13360,N13361,N13362,N13363,N13364,N13365,N13366,N13367,N13368,
N13369,N13370,N13371,N13372,N13373,N13374,N13375,N13376,N13377,N13378,
N13379,N13380,N13381,N13382,N13383,N13384,N13385,N13386,N13387,N13388,
N13389,N13390,N13391,N13392,N13393,N13394,N13395,N13396,N13397,N13398,
N13399,N13400,N13401,N13402,N13403,N13404,N13405,N13406,N13407,N13408,
N13409,N13410,N13411,N13412,N13413,N13414,N13415,N13416,N13417,N13418,
N13419,N13420,N13421,N13422,N13423,N13424,N13425,N13426,N13427,N13428,
N13429,N13430,N13431,N13432,N13433,N13434,N13435,N13436,N13437,N13438,
N13439,N13440,N13441,N13442,N13443,N13444,N13445,N13446,N13447,N13448,
N13449,N13450,N13451,N13452,N13453,N13454,N13455,N13456,N13457,N13458,
N13459,N13460,N13461,N13462,N13463,N13464,N13465,N13466,N13467,N13468,
N13469,N13470,N13471,N13472,N13473,N13474,N13475,N13476,N13477,N13478,
N13479,N13480,N13481,N13482,N13483,N13484,N13485,N13486,N13487,N13488,
N13489,N13490,N13491,N13492,N13493,N13494,N13495,N13496,N13497,N13498,
N13499,N13500,N13501,N13502,N13503,N13504,N13505,N13506,N13507,N13508,
N13509,N13510,N13511,N13512,N13513,N13514,N13515,N13516,N13517,N13518,
N13519,N13520,N13521,N13522,N13523,N13524,N13525,N13526,N13527,N13528,
N13529,N13530,N13531,N13532,N13533,N13534,N13535,N13536,N13537,N13538,
N13539,N13540,N13541,N13542,N13543,N13544,N13545,N13546,N13547,N13548,
N13549,N13550,N13551,N13552,N13553,N13554,N13555,N13556,N13557,N13558,
N13559,N13560,N13561,N13562,N13563,N13564,N13565,N13566,N13567,N13568,
N13569,N13570,N13571,N13572,N13573,N13574,N13575,N13576,N13577,N13578,
N13579,N13580,N13581,N13582,N13583,N13584,N13585,N13586,N13587,N13588,
N13589,N13590,N13591,N13592,N13593,N13594,N13595,N13596,N13597,N13598,
N13599,N13600,N13601,N13602,N13603,N13604,N13605,N13606,N13607,N13608,
N13609,N13610,N13611,N13612,N13613,N13614,N13615,N13616,N13617,N13618,
N13619,N13620,N13621,N13622,N13623,N13624,N13625,N13626,N13627,N13628,
N13629,N13630,N13631,N13632,N13633,N13634,N13635,N13636,N13637,N13638,
N13639,N13640,N13641,N13642,N13643,N13644,N13645,N13646,N13647,N13648,
N13649,N13650,N13651,N13652,N13653,N13654,N13655,N13656,N13657,N13658,
N13659,N13660,N13661,N13662,N13663,N13664,N13665,N13666,N13667,N13668,
N13669,N13670,N13671,N13672,N13673,N13674,N13675,N13676,N13677,N13678,
N13679,N13680,N13681,N13682,N13683,N13684,N13685,N13686,N13687,N13688,
N13689,N13690,N13691,N13692,N13693,N13694,N13695,N13696,N13697,N13698,
N13699,N13700,N13701,N13702,N13703,N13704,N13705,N13706,N13707,N13708,
N13709,N13710,N13711,N13712,N13713,N13714,N13715,N13716,N13717,N13718,
N13719,N13720,N13721,N13722,N13723,N13724,N13725,N13726,N13727,N13728,
N13729,N13730,N13731,N13732,N13733,N13734,N13735,N13736,N13737,N13738,
N13739,N13740,N13741,N13742,N13743,N13744,N13745,N13746,N13747,N13748,
N13749,N13750,N13751,N13752,N13753,N13754,N13755,N13756,N13757,N13758,
N13759,N13760,N13761,N13762,N13763,N13764,N13765,N13766,N13767,N13768,
N13769,N13770,N13771,N13772,N13773,N13774,N13775,N13776,N13777,N13778,
N13779,N13780,N13781,N13782,N13783,N13784,N13785,N13786,N13787,N13788,
N13789,N13790,N13791,N13792,N13793,N13794,N13795,N13796,N13797,N13798,
N13799,N13800,N13801,N13802,N13803,N13804,N13805,N13806,N13807,N13808,
N13809,N13810,N13811,N13812,N13813,N13814,N13815,N13816,N13817,N13818,
N13819,N13820,N13821,N13822,N13823,N13824,N13825,N13826,N13827,N13828,
N13829,N13830,N13831,N13832,N13833,N13834,N13835,N13836,N13837,N13838,
N13839,N13840,N13841,N13842,N13843,N13844,N13845,N13846,N13847,N13848,
N13849,N13850,N13851,N13852,N13853,N13854,N13855,N13856,N13857,N13858,
N13859,N13860,N13861,N13862,N13863,N13864,N13865,N13866,N13867,N13868,
N13869,N13870,N13871,N13872,N13873,N13874,N13875,N13876,N13877,N13878,
N13879,N13880,N13881,N13882,N13883,N13884,N13885,N13886,N13887,N13888,
N13889,N13890,N13891,N13892,N13893,N13894,N13895,N13896,N13897,N13898,
N13899,N13900,N13901,N13902,N13903,N13904,N13905,N13906,N13907,N13908,
N13909,N13910,N13911,N13912,N13913,N13914,N13915,N13916,N13917,N13918,
N13919,N13920,N13921,N13922,N13923,N13924,N13925,N13926,N13927,N13928,
N13929,N13930,N13931,N13932,N13933,N13934,N13935,N13936,N13937,N13938,
N13939,N13940,N13941,N13942,N13943,N13944,N13945,N13946,N13947,N13948,
N13949,N13950,N13951,N13952,N13953,N13954,N13955,N13956,N13957,N13958,
N13959,N13960,N13961,N13962,N13963,N13964,N13965,N13966,N13967,N13968,
N13969,N13970,N13971,N13972,N13973,N13974,N13975,N13976,N13977,N13978,
N13979,N13980,N13981,N13982,N13983,N13984,N13985,N13986,N13987,N13988,
N13989,N13990,N13991,N13992,N13993,N13994,N13995,N13996,N13997,N13998,
N13999,N14000,N14001,N14002,N14003,N14004,N14005,N14006,N14007,N14008,
N14009,N14010,N14011,N14012,N14013,N14014,N14015,N14016,N14017,N14018,
N14019,N14020,N14021,N14022,N14023,N14024,N14025,N14026,N14027,N14028,
N14029,N14030,N14031,N14032,N14033,N14034,N14035,N14036,N14037,N14038,
N14039,N14040,N14041,N14042,N14043,N14044,N14045,N14046,N14047,N14048,
N14049,N14050,N14051,N14052,N14053,N14054,N14055,N14056,N14057,N14058,
N14059,N14060,N14061,N14062,N14063,N14064,N14065,N14066,N14067,N14068,
N14069,N14070,N14071,N14072,N14073,N14074,N14075,N14076,N14077,N14078,
N14079,N14080,N14081,N14082,N14083,N14084,N14085,N14086,N14087,N14088,
N14089,N14090,N14091,N14092,N14093,N14094,N14095,N14096,N14097,N14098,
N14099,N14100,N14101,N14102,N14103,N14104,N14105,N14106,N14107,N14108,
N14109,N14110,N14111,N14112,N14113,N14114,N14115,N14116,N14117,N14118,
N14119,N14120,N14121,N14122,N14123,N14124,N14125,N14126,N14127,N14128,
N14129,N14130,N14131,N14132,N14133,N14134,N14135,N14136,N14137,N14138,
N14139,N14140,N14141,N14142,N14143,N14144,N14145,N14146,N14147,N14148,
N14149,N14150,N14151,N14152,N14153,N14154,N14155,N14156,N14157,N14158,
N14159,N14160,N14161,N14162,N14163,N14164,N14165,N14166,N14167,N14168,
N14169,N14170,N14171,N14172,N14173,N14174,N14175,N14176,N14177,N14178,
N14179,N14180,N14181,N14182,N14183,N14184,N14185,N14186,N14187,N14188,
N14189,N14190,N14191,N14192,N14193,N14194,N14195,N14196,N14197,N14198,
N14199,N14200,N14201,N14202,N14203,N14204,N14205,N14206,N14207,N14208,
N14209,N14210,N14211,N14212,N14213,N14214,N14215,N14216,N14217,N14218,
N14219,N14220,N14221,N14222,N14223,N14224,N14225,N14226,N14227,N14228,
N14229,N14230,N14231,N14232,N14233,N14234,N14235,N14236,N14237,N14238,
N14239,N14240,N14241,N14242,N14243,N14244,N14245,N14246,N14247,N14248,
N14249,N14250,N14251,N14252,N14253,N14254,N14255,N14256,N14257,N14258,
N14259,N14260,N14261,N14262,N14263,N14264,N14265,N14266,N14267,N14268,
N14269,N14270,N14271,N14272,N14273,N14274,N14275,N14276,N14277,N14278,
N14279,N14280,N14281,N14282,N14283,N14284,N14285,N14286,N14287,N14288,
N14289,N14290,N14291,N14292,N14293,N14294,N14295,N14296,N14297,N14298,
N14299,N14300,N14301,N14302,N14303,N14304,N14305,N14306,N14307,N14308,
N14309,N14310,N14311,N14312,N14313,N14314,N14315,N14316,N14317,N14318,
N14319,N14320,N14321,N14322,N14323,N14324,N14325,N14326,N14327,N14328,
N14329,N14330,N14331,N14332,N14333,N14334,N14335,N14336,N14337,N14338,
N14339,N14340,N14341,N14342,N14343,N14344,N14345,N14346,N14347,N14348,
N14349,N14350,N14351,N14352,N14353,N14354,N14355,N14356,N14357,N14358,
N14359,N14360,N14361,N14362,N14363,N14364,N14365,N14366,N14367,N14368,
N14369,N14370,N14371,N14372,N14373,N14374,N14375,N14376,N14377,N14378,
N14379,N14380,N14381,N14382,N14383,N14384,N14385,N14386,N14387,N14388,
N14389,N14390,N14391,N14392,N14393,N14394,N14395,N14396,N14397,N14398,
N14399,N14400,N14401,N14402,N14403,N14404,N14405,N14406,N14407,N14408,
N14409,N14410,N14411,N14412,N14413,N14414,N14415,N14416,N14417,N14418,
N14419,N14420,N14421,N14422,N14423,N14424,N14425,N14426,N14427,N14428,
N14429,N14430,N14431,N14432,N14433,N14434,N14435,N14436,N14437,N14438,
N14439,N14440,N14441,N14442,N14443,N14444,N14445,N14446,N14447,N14448,
N14449,N14450,N14451,N14452,N14453,N14454,N14455,N14456,N14457,N14458,
N14459,N14460,N14461,N14462,N14463,N14464,N14465,N14466,N14467,N14468,
N14469,N14470,N14471,N14472,N14473,N14474,N14475,N14476,N14477,N14478,
N14479,N14480,N14481,N14482,N14483,N14484,N14485,N14486,N14487,N14488,
N14489,N14490,N14491,N14492,N14493,N14494,N14495,N14496,N14497,N14498,
N14499,N14500,N14501,N14502,N14503,N14504,N14505,N14506,N14507,N14508,
N14509,N14510,N14511,N14512,N14513,N14514,N14515,N14516,N14517,N14518,
N14519,N14520,N14521,N14522,N14523,N14524,N14525,N14526,N14527,N14528,
N14529,N14530,N14531,N14532,N14533,N14534,N14535,N14536,N14537,N14538,
N14539,N14540,N14541,N14542,N14543,N14544,N14545,N14546,N14547,N14548,
N14549,N14550,N14551,N14552,N14553,N14554,N14555,N14556,N14557,N14558,
N14559,N14560,N14561,N14562,N14563,N14564,N14565,N14566,N14567,N14568,
N14569,N14570,N14571,N14572,N14573,N14574,N14575,N14576,N14577,N14578,
N14579,N14580,N14581,N14582,N14583,N14584,N14585,N14586,N14587,N14588,
N14589,N14590,N14591,N14592,N14593,N14594,N14595,N14596,N14597,N14598,
N14599,N14600,N14601,N14602,N14603,N14604,N14605,N14606,N14607,N14608,
N14609,N14610,N14611,N14612,N14613,N14614,N14615,N14616,N14617,N14618,
N14619,N14620,N14621,N14622,N14623,N14624,N14625,N14626,N14627,N14628,
N14629,N14630,N14631,N14632,N14633,N14634,N14635,N14636,N14637,N14638,
N14639,N14640,N14641,N14642,N14643,N14644,N14645,N14646,N14647,N14648,
N14649,N14650,N14651,N14652,N14653,N14654,N14655,N14656,N14657,N14658,
N14659,N14660,N14661,N14662,N14663,N14664,N14665,N14666,N14667,N14668,
N14669,N14670,N14671,N14672,N14673,N14674,N14675,N14676,N14677,N14678,
N14679,N14680,N14681,N14682,N14683,N14684,N14685,N14686,N14687,N14688,
N14689,N14690,N14691,N14692,N14693,N14694,N14695,N14696,N14697,N14698,
N14699,N14700,N14701,N14702,N14703,N14704,N14705,N14706,N14707,N14708,
N14709,N14710,N14711,N14712,N14713,N14714,N14715,N14716,N14717,N14718,
N14719,N14720,N14721,N14722,N14723,N14724,N14725,N14726,N14727,N14728,
N14729,N14730,N14731,N14732,N14733,N14734,N14735,N14736,N14737,N14738,
N14739,N14740,N14741,N14742,N14743,N14744,N14745,N14746,N14747,N14748,
N14749,N14750,N14751,N14752,N14753,N14754,N14755,N14756,N14757,N14758,
N14759,N14760,N14761,N14762,N14763,N14764,N14765,N14766,N14767,N14768,
N14769,N14770,N14771,N14772,N14773,N14774,N14775,N14776,N14777,N14778,
N14779,N14780,N14781,N14782,N14783,N14784,N14785,N14786,N14787,N14788,
N14789,N14790,N14791,N14792,N14793,N14794,N14795,N14796,N14797,N14798,
N14799,N14800,N14801,N14802,N14803,N14804,N14805,N14806,N14807,N14808,
N14809,N14810,N14811,N14812,N14813,N14814,N14815,N14816,N14817,N14818,
N14819,N14820,N14821,N14822,N14823,N14824,N14825,N14826,N14827,N14828,
N14829,N14830,N14831,N14832,N14833,N14834,N14835,N14836,N14837,N14838,
N14839,N14840,N14841,N14842,N14843,N14844,N14845,N14846,N14847,N14848,
N14849,N14850,N14851,N14852,N14853,N14854,N14855,N14856,N14857,N14858,
N14859,N14860,N14861,N14862,N14863,N14864,N14865,N14866,N14867,N14868,
N14869,N14870,N14871,N14872,N14873,N14874,N14875,N14876,N14877,N14878,
N14879,N14880,N14881,N14882,N14883,N14884,N14885,N14886,N14887,N14888,
N14889,N14890,N14891,N14892,N14893,N14894,N14895,N14896,N14897,N14898,
N14899,N14900,N14901,N14902,N14903,N14904,N14905,N14906,N14907,N14908,
N14909,N14910,N14911,N14912,N14913,N14914,N14915,N14916,N14917,N14918,
N14919,N14920,N14921,N14922,N14923,N14924,N14925,N14926,N14927,N14928,
N14929,N14930,N14931,N14932,N14933,N14934,N14935,N14936,N14937,N14938,
N14939,N14940,N14941,N14942,N14943,N14944,N14945,N14946,N14947,N14948,
N14949,N14950,N14951,N14952,N14953,N14954,N14955,N14956,N14957,N14958,
N14959,N14960,N14961,N14962,N14963,N14964,N14965,N14966,N14967,N14968,
N14969,N14970,N14971,N14972,N14973,N14974,N14975,N14976,N14977,N14978,
N14979,N14980,N14981,N14982,N14983,N14984,N14985,N14986,N14987,N14988,
N14989,N14990,N14991,N14992,N14993,N14994,N14995,N14996,N14997,N14998,
N14999,N15000,N15001,N15002,N15003,N15004,N15005,N15006,N15007,N15008,
N15009,N15010,N15011,N15012,N15013,N15014,N15015,N15016,N15017,N15018,
N15019,N15020,N15021,N15022,N15023,N15024,N15025,N15026,N15027,N15028,
N15029,N15030,N15031,N15032,N15033,N15034,N15035,N15036,N15037,N15038,
N15039,N15040,N15041,N15042,N15043,N15044,N15045,N15046,N15047,N15048,
N15049,N15050,N15051,N15052,N15053,N15054,N15055,N15056,N15057,N15058,
N15059,N15060,N15061,N15062,N15063,N15064,N15065,N15066,N15067,N15068,
N15069,N15070,N15071,N15072,N15073,N15074,N15075,N15076,N15077,N15078,
N15079,N15080,N15081,N15082,N15083,N15084,N15085,N15086,N15087,N15088,
N15089,N15090,N15091,N15092,N15093,N15094,N15095,N15096,N15097,N15098,
N15099,N15100,N15101,N15102,N15103,N15104,N15105,N15106,N15107,N15108,
N15109,N15110,N15111,N15112,N15113,N15114,N15115,N15116,N15117,N15118,
N15119,N15120,N15121,N15122,N15123,N15124,N15125,N15126,N15127,N15128,
N15129,N15130,N15131,N15132,N15133,N15134,N15135,N15136,N15137,N15138,
N15139,N15140,N15141,N15142,N15143,N15144,N15145,N15146,N15147,N15148,
N15149,N15150,N15151,N15152,N15153,N15154,N15155,N15156,N15157,N15158,
N15159,N15160,N15161,N15162,N15163,N15164,N15165,N15166,N15167,N15168,
N15169,N15170,N15171,N15172,N15173,N15174,N15175,N15176,N15177,N15178,
N15179,N15180,N15181,N15182,N15183,N15184,N15185,N15186,N15187,N15188,
N15189,N15190,N15191,N15192,N15193,N15194,N15195,N15196,N15197,N15198,
N15199,N15200,N15201,N15202,N15203,N15204,N15205,N15206,N15207,N15208,
N15209,N15210,N15211,N15212,N15213,N15214,N15215,N15216,N15217,N15218,
N15219,N15220,N15221,N15222,N15223,N15224,N15225,N15226,N15227,N15228,
N15229,N15230,N15231,N15232,N15233,N15234,N15235,N15236,N15237,N15238,
N15239,N15240,N15241,N15242,N15243,N15244,N15245,N15246,N15247,N15248,
N15249,N15250,N15251,N15252,N15253,N15254,N15255,N15256,N15257,N15258,
N15259,N15260,N15261,N15262,N15263,N15264,N15265,N15266,N15267,N15268,
N15269,N15270,N15271,N15272,N15273,N15274,N15275,N15276,N15277,N15278,
N15279,N15280,N15281,N15282,N15283,N15284,N15285,N15286,N15287,N15288,
N15289,N15290,N15291,N15292,N15293,N15294,N15295,N15296,N15297,N15298,
N15299,N15300,N15301,N15302,N15303,N15304,N15305,N15306,N15307,N15308,
N15309,N15310,N15311,N15312,N15313,N15314,N15315,N15316,N15317,N15318,
N15319,N15320,N15321,N15322,N15323,N15324,N15325,N15326,N15327,N15328,
N15329,N15330,N15331,N15332,N15333,N15334,N15335,N15336,N15337,N15338,
N15339,N15340,N15341,N15342,N15343,N15344,N15345,N15346,N15347,N15348,
N15349,N15350,N15351,N15352,N15353,N15354,N15355,N15356,N15357,N15358,
N15359,N15360,N15361,N15362,N15363,N15364,N15365,N15366,N15367,N15368,
N15369,N15370,N15371,N15372,N15373,N15374,N15375,N15376,N15377,N15378,
N15379,N15380,N15381,N15382,N15383,N15384,N15385,N15386,N15387,N15388,
N15389,N15390,N15391,N15392,N15393,N15394,N15395,N15396,N15397,N15398,
N15399,N15400,N15401,N15402,N15403,N15404,N15405,N15406,N15407,N15408,
N15409,N15410,N15411,N15412,N15413,N15414,N15415,N15416,N15417,N15418,
N15419,N15420,N15421,N15422,N15423,N15424,N15425,N15426,N15427,N15428,
N15429,N15430,N15431,N15432,N15433,N15434,N15435,N15436,N15437,N15438,
N15439,N15440,N15441,N15442,N15443,N15444,N15445,N15446,N15447,N15448,
N15449,N15450,N15451,N15452,N15453,N15454,N15455,N15456,N15457,N15458,
N15459,N15460,N15461,N15462,N15463,N15464,N15465,N15466,N15467,N15468,
N15469,N15470,N15471,N15472,N15473,N15474,N15475,N15476,N15477,N15478,
N15479,N15480,N15481,N15482,N15483,N15484,N15485,N15486,N15487,N15488,
N15489,N15490,N15491,N15492,N15493,N15494,N15495,N15496,N15497,N15498,
N15499,N15500,N15501,N15502,N15503,N15504,N15505,N15506,N15507,N15508,
N15509,N15510,N15511,N15512,N15513,N15514,N15515,N15516,N15517,N15518,
N15519,N15520,N15521,N15522,N15523,N15524,N15525,N15526,N15527,N15528,
N15529,N15530,N15531,N15532,N15533,N15534,N15535,N15536,N15537,N15538,
N15539,N15540,N15541,N15542,N15543,N15544,N15545,N15546,N15547,N15548,
N15549,N15550,N15551,N15552,N15553,N15554,N15555,N15556,N15557,N15558,
N15559,N15560,N15561,N15562,N15563,N15564,N15565,N15566,N15567,N15568,
N15569,N15570,N15571,N15572,N15573,N15574,N15575,N15576,N15577,N15578,
N15579,N15580,N15581,N15582,N15583,N15584,N15585,N15586,N15587,N15588,
N15589,N15590,N15591,N15592,N15593,N15594,N15595,N15596,N15597,N15598,
N15599,N15600,N15601,N15602,N15603,N15604,N15605,N15606,N15607,N15608,
N15609,N15610,N15611,N15612,N15613,N15614,N15615,N15616,N15617,N15618,
N15619,N15620,N15621,N15622,N15623,N15624,N15625,N15626,N15627,N15628,
N15629,N15630,N15631,N15632,N15633,N15634,N15635,N15636,N15637,N15638,
N15639,N15640,N15641,N15642,N15643,N15644,N15645,N15646,N15647,N15648,
N15649,N15650,N15651,N15652,N15653,N15654,N15655,N15656,N15657,N15658,
N15659,N15660,N15661,N15662,N15663,N15664,N15665,N15666,N15667,N15668,
N15669,N15670,N15671,N15672,N15673,N15674,N15675,N15676,N15677,N15678,
N15679,N15680,N15681,N15682,N15683,N15684,N15685,N15686,N15687,N15688,
N15689,N15690,N15691,N15692,N15693,N15694,N15695,N15696,N15697,N15698,
N15699,N15700,N15701,N15702,N15703,N15704,N15705,N15706,N15707,N15708,
N15709,N15710,N15711,N15712,N15713,N15714,N15715,N15716,N15717,N15718,
N15719,N15720,N15721,N15722,N15723,N15724,N15725,N15726,N15727,N15728,
N15729,N15730,N15731,N15732,N15733,N15734,N15735,N15736,N15737,N15738,
N15739,N15740,N15741,N15742,N15743,N15744,N15745,N15746,N15747,N15748,
N15749,N15750,N15751,N15752,N15753,N15754,N15755,N15756,N15757,N15758,
N15759,N15760,N15761,N15762,N15763,N15764,N15765,N15766,N15767,N15768,
N15769,N15770,N15771,N15772,N15773,N15774,N15775,N15776,N15777,N15778,
N15779,N15780,N15781,N15782,N15783,N15784,N15785,N15786,N15787,N15788,
N15789,N15790,N15791,N15792,N15793,N15794,N15795,N15796,N15797,N15798,
N15799,N15800,N15801,N15802,N15803,N15804,N15805,N15806,N15807,N15808,
N15809,N15810,N15811,N15812,N15813,N15814,N15815,N15816,N15817,N15818,
N15819,N15820,N15821,N15822,N15823,N15824,N15825,N15826,N15827,N15828,
N15829,N15830,N15831,N15832,N15833,N15834,N15835,N15836,N15837,N15838,
N15839,N15840,N15841,N15842,N15843,N15844,N15845,N15846,N15847,N15848,
N15849,N15850,N15851,N15852,N15853,N15854,N15855,N15856,N15857,N15858,
N15859,N15860,N15861,N15862,N15863,N15864,N15865,N15866,N15867,N15868,
N15869,N15870,N15871,N15872,N15873,N15874,N15875,N15876,N15877,N15878,
N15879,N15880,N15881,N15882,N15883,N15884,N15885,N15886,N15887,N15888,
N15889,N15890,N15891,N15892,N15893,N15894,N15895,N15896,N15897,N15898,
N15899,N15900,N15901,N15902,N15903,N15904,N15905,N15906,N15907,N15908,
N15909,N15910,N15911,N15912,N15913,N15914,N15915,N15916,N15917,N15918,
N15919,N15920,N15921,N15922,N15923,N15924,N15925,N15926,N15927,N15928,
N15929,N15930,N15931,N15932,N15933,N15934,N15935,N15936,N15937,N15938,
N15939,N15940,N15941,N15942,N15943,N15944,N15945,N15946,N15947,N15948,
N15949,N15950,N15951,N15952,N15953,N15954,N15955,N15956,N15957,N15958,
N15959,N15960,N15961,N15962,N15963,N15964,N15965,N15966,N15967,N15968,
N15969,N15970,N15971,N15972,N15973,N15974,N15975,N15976,N15977,N15978,
N15979,N15980,N15981,N15982,N15983,N15984,N15985,N15986,N15987,N15988,
N15989,N15990,N15991,N15992,N15993,N15994,N15995,N15996,N15997,N15998,
N15999,N16000,N16001,N16002,N16003,N16004,N16005,N16006,N16007,N16008,
N16009,N16010,N16011,N16012,N16013,N16014,N16015,N16016,N16017,N16018,
N16019,N16020,N16021,N16022,N16023,N16024,N16025,N16026,N16027,N16028,
N16029,N16030,N16031,N16032,N16033,N16034,N16035,N16036,N16037,N16038,
N16039,N16040,N16041,N16042,N16043,N16044,N16045,N16046,N16047,N16048,
N16049,N16050,N16051,N16052,N16053,N16054,N16055,N16056,N16057,N16058,
N16059,N16060,N16061,N16062,N16063,N16064,N16065,N16066,N16067,N16068,
N16069,N16070,N16071,N16072,N16073,N16074,N16075,N16076,N16077,N16078,
N16079,N16080,N16081,N16082,N16083,N16084,N16085,N16086,N16087,N16088,
N16089,N16090,N16091,N16092,N16093,N16094,N16095,N16096,N16097,N16098,
N16099,N16100,N16101,N16102,N16103,N16104,N16105,N16106,N16107,N16108,
N16109,N16110,N16111,N16112,N16113,N16114,N16115,N16116,N16117,N16118,
N16119,N16120,N16121,N16122,N16123,N16124,N16125,N16126,N16127,N16128,
N16129,N16130,N16131,N16132,N16133,N16134,N16135,N16136,N16137,N16138,
N16139,N16140,N16141,N16142,N16143,N16144,N16145,N16146,N16147,N16148,
N16149,N16150,N16151,N16152,N16153,N16154,N16155,N16156,N16157,N16158,
N16159,N16160,N16161,N16162,N16163,N16164,N16165,N16166,N16167,N16168,
N16169,N16170,N16171,N16172,N16173,N16174,N16175,N16176,N16177,N16178,
N16179,N16180,N16181,N16182,N16183,N16184,N16185,N16186,N16187,N16188,
N16189,N16190,N16191,N16192,N16193,N16194,N16195,N16196,N16197,N16198,
N16199,N16200,N16201,N16202,N16203,N16204,N16205,N16206,N16207,N16208,
N16209,N16210,N16211,N16212,N16213,N16214,N16215,N16216,N16217,N16218,
N16219,N16220,N16221,N16222,N16223,N16224,N16225,N16226,N16227,N16228,
N16229,N16230,N16231,N16232,N16233,N16234,N16235,N16236,N16237,N16238,
N16239,N16240,N16241,N16242,N16243,N16244,N16245,N16246,N16247,N16248,
N16249,N16250,N16251,N16252,N16253,N16254,N16255,N16256,N16257,N16258,
N16259,N16260,N16261,N16262,N16263,N16264,N16265,N16266,N16267,N16268,
N16269,N16270,N16271,N16272,N16273,N16274,N16275,N16276,N16277,N16278,
N16279,N16280,N16281,N16282,N16283,N16284,N16285,N16286,N16287,N16288,
N16289,N16290,N16291,N16292,N16293,N16294,N16295,N16296,N16297,N16298,
N16299,N16300,N16301,N16302,N16303,N16304,N16305,N16306,N16307,N16308,
N16309,N16310,N16311,N16312,N16313,N16314,N16315,N16316,N16317,N16318,
N16319,N16320,N16321,N16322,N16323,N16324,N16325,N16326,N16327,N16328,
N16329,N16330,N16331,N16332,N16333,N16334,N16335,N16336,N16337,N16338,
N16339,N16340,N16341,N16342,N16343,N16344,N16345,N16346,N16347,N16348,
N16349,N16350,N16351,N16352,N16353,N16354,N16355,N16356,N16357,N16358,
N16359,N16360,N16361,N16362,N16363,N16364,N16365,N16366,N16367,N16368,
N16369,N16370,N16371,N16372,N16373,N16374,N16375,N16376,N16377,N16378,
N16379,N16380,N16381,N16382,N16383,N16384,N16385,N16386,N16387,N16388,
N16389,N16390,N16391,N16392,N16393,N16394,N16395,N16396,N16397,N16398,
N16399,N16400,N16401,N16402,N16403,N16404,N16405,N16406,N16407,N16408,
N16409,N16410,N16411,N16412,N16413,N16414,N16415,N16416,N16417,N16418,
N16419,N16420,N16421,N16422,N16423,N16424,N16425,N16426,N16427,N16428,
N16429,N16430,N16431,N16432,N16433,N16434,N16435,N16436,N16437,N16438,
N16439,N16440,N16441,N16442,N16443,N16444,N16445,N16446,N16447,N16448,
N16449,N16450,N16451,N16452,N16453,N16454,N16455,N16456,N16457,N16458,
N16459,N16460,N16461,N16462,N16463,N16464,N16465,N16466,N16467,N16468,
N16469,N16470,N16471,N16472,N16473,N16474,N16475,N16476,N16477,N16478,
N16479,N16480,N16481,N16482,N16483,N16484,N16485,N16486,N16487,N16488,
N16489,N16490,N16491,N16492,N16493,N16494,N16495,N16496,N16497,N16498,
N16499,N16500,N16501,N16502,N16503,N16504,N16505,N16506,N16507,N16508,
N16509,N16510,N16511,N16512,N16513,N16514,N16515,N16516,N16517,N16518,
N16519,N16520,N16521,N16522,N16523,N16524,N16525,N16526,N16527,N16528,
N16529,N16530,N16531,N16532,N16533,N16534,N16535,N16536,N16537,N16538,
N16539,N16540,N16541,N16542,N16543,N16544,N16545,N16546,N16547,N16548,
N16549,N16550,N16551,N16552,N16553,N16554,N16555,N16556,N16557,N16558,
N16559,N16560,N16561,N16562,N16563,N16564,N16565,N16566,N16567,N16568,
N16569,N16570,N16571,N16572,N16573,N16574,N16575,N16576,N16577,N16578,
N16579,N16580,N16581,N16582,N16583,N16584,N16585,N16586,N16587,N16588,
N16589,N16590,N16591,N16592,N16593,N16594,N16595,N16596,N16597,N16598,
N16599,N16600,N16601,N16602,N16603,N16604,N16605,N16606,N16607,N16608,
N16609,N16610,N16611,N16612,N16613,N16614,N16615,N16616,N16617,N16618,
N16619,N16620,N16621,N16622,N16623,N16624,N16625,N16626,N16627,N16628,
N16629,N16630,N16631,N16632,N16633,N16634,N16635,N16636,N16637,N16638,
N16639,N16640,N16641,N16642,N16643,N16644,N16645,N16646,N16647,N16648,
N16649,N16650,N16651,N16652,N16653,N16654,N16655,N16656,N16657,N16658,
N16659,N16660,N16661,N16662,N16663,N16664,N16665,N16666,N16667,N16668,
N16669,N16670,N16671,N16672,N16673,N16674,N16675,N16676,N16677,N16678,
N16679,N16680,N16681,N16682,N16683,N16684,N16685,N16686,N16687,N16688,
N16689,N16690,N16691,N16692,N16693,N16694,N16695,N16696,N16697,N16698,
N16699,N16700,N16701,N16702,N16703,N16704,N16705,N16706,N16707,N16708,
N16709,N16710,N16711,N16712,N16713,N16714,N16715,N16716,N16717,N16718,
N16719,N16720,N16721,N16722,N16723,N16724,N16725,N16726,N16727,N16728,
N16729,N16730,N16731,N16732,N16733,N16734,N16735,N16736,N16737,N16738,
N16739,N16740,N16741,N16742,N16743,N16744,N16745,N16746,N16747,N16748,
N16749,N16750,N16751,N16752,N16753,N16754,N16755,N16756,N16757,N16758,
N16759,N16760,N16761,N16762,N16763,N16764,N16765,N16766,N16767,N16768,
N16769,N16770,N16771,N16772,N16773,N16774,N16775,N16776,N16777,N16778,
N16779,N16780,N16781,N16782,N16783,N16784,N16785,N16786,N16787,N16788,
N16789,N16790,N16791,N16792,N16793,N16794,N16795,N16796,N16797,N16798,
N16799,N16800,N16801,N16802,N16803,N16804,N16805,N16806,N16807,N16808,
N16809,N16810,N16811,N16812,N16813,N16814,N16815,N16816,N16817,N16818,
N16819,N16820,N16821,N16822,N16823,N16824,N16825,N16826,N16827,N16828,
N16829,N16830,N16831,N16832,N16833,N16834,N16835,N16836,N16837,N16838,
N16839,N16840,N16841,N16842,N16843,N16844,N16845,N16846,N16847,N16848,
N16849,N16850,N16851,N16852,N16853,N16854,N16855,N16856,N16857,N16858,
N16859,N16860,N16861,N16862,N16863,N16864,N16865,N16866,N16867,N16868,
N16869,N16870,N16871,N16872,N16873,N16874,N16875,N16876,N16877,N16878,
N16879,N16880,N16881,N16882,N16883,N16884,N16885,N16886,N16887,N16888,
N16889,N16890,N16891,N16892,N16893,N16894,N16895,N16896,N16897,N16898,
N16899,N16900,N16901,N16902,N16903,N16904,N16905,N16906,N16907,N16908,
N16909,N16910,N16911,N16912,N16913,N16914,N16915,N16916,N16917,N16918,
N16919,N16920,N16921,N16922,N16923,N16924,N16925,N16926,N16927,N16928,
N16929,N16930,N16931,N16932,N16933,N16934,N16935,N16936,N16937,N16938,
N16939,N16940,N16941,N16942,N16943,N16944,N16945,N16946,N16947,N16948,
N16949,N16950,N16951,N16952,N16953,N16954,N16955,N16956,N16957,N16958,
N16959,N16960,N16961,N16962,N16963,N16964,N16965,N16966,N16967,N16968,
N16969,N16970,N16971,N16972,N16973,N16974,N16975,N16976,N16977,N16978,
N16979,N16980,N16981,N16982,N16983,N16984,N16985,N16986,N16987,N16988,
N16989,N16990,N16991,N16992,N16993,N16994,N16995,N16996,N16997,N16998,
N16999,N17000,N17001,N17002,N17003,N17004,N17005,N17006,N17007,N17008,
N17009,N17010,N17011,N17012,N17013,N17014,N17015,N17016,N17017,N17018,
N17019,N17020,N17021,N17022,N17023,N17024,N17025,N17026,N17027,N17028,
N17029,N17030,N17031,N17032,N17033,N17034,N17035,N17036,N17037,N17038,
N17039,N17040,N17041,N17042,N17043,N17044,N17045,N17046,N17047,N17048,
N17049,N17050,N17051,N17052,N17053,N17054,N17055,N17056,N17057,N17058,
N17059,N17060,N17061,N17062,N17063,N17064,N17065,N17066,N17067,N17068,
N17069,N17070,N17071,N17072,N17073,N17074,N17075,N17076,N17077,N17078,
N17079,N17080,N17081,N17082,N17083,N17084,N17085,N17086,N17087,N17088,
N17089,N17090,N17091,N17092,N17093,N17094,N17095,N17096,N17097,N17098,
N17099,N17100,N17101,N17102,N17103,N17104,N17105,N17106,N17107,N17108,
N17109,N17110,N17111,N17112,N17113,N17114,N17115,N17116,N17117,N17118,
N17119,N17120,N17121,N17122,N17123,N17124,N17125,N17126,N17127,N17128,
N17129,N17130,N17131,N17132,N17133,N17134,N17135,N17136,N17137,N17138,
N17139,N17140,N17141,N17142,N17143,N17144,N17145,N17146,N17147,N17148,
N17149,N17150,N17151,N17152,N17153,N17154,N17155,N17156,N17157,N17158,
N17159,N17160,N17161,N17162,N17163,N17164,N17165,N17166,N17167,N17168,
N17169,N17170,N17171,N17172,N17173,N17174,N17175,N17176,N17177,N17178,
N17179,N17180,N17181,N17182,N17183,N17184,N17185,N17186,N17187,N17188,
N17189,N17190,N17191,N17192,N17193,N17194,N17195,N17196,N17197,N17198,
N17199,N17200,N17201,N17202,N17203,N17204,N17205,N17206,N17207,N17208,
N17209,N17210,N17211,N17212,N17213,N17214,N17215,N17216,N17217,N17218,
N17219,N17220,N17221,N17222,N17223,N17224,N17225,N17226,N17227,N17228,
N17229,N17230,N17231,N17232,N17233,N17234,N17235,N17236,N17237,N17238,
N17239,N17240,N17241,N17242,N17243,N17244,N17245,N17246,N17247,N17248,
N17249,N17250,N17251,N17252,N17253,N17254,N17255,N17256,N17257,N17258,
N17259,N17260,N17261,N17262,N17263,N17264,N17265,N17266,N17267,N17268,
N17269,N17270,N17271,N17272,N17273,N17274,N17275,N17276,N17277,N17278,
N17279,N17280,N17281,N17282,N17283,N17284,N17285,N17286,N17287,N17288,
N17289,N17290,N17291,N17292,N17293,N17294,N17295,N17296,N17297,N17298,
N17299,N17300,N17301,N17302,N17303,N17304,N17305,N17306,N17307,N17308,
N17309,N17310,N17311,N17312,N17313,N17314,N17315,N17316,N17317,N17318,
N17319,N17320,N17321,N17322,N17323,N17324,N17325,N17326,N17327,N17328,
N17329,N17330,N17331,N17332,N17333,N17334,N17335,N17336,N17337,N17338,
N17339,N17340,N17341,N17342,N17343,N17344,N17345,N17346,N17347,N17348,
N17349,N17350,N17351,N17352,N17353,N17354,N17355,N17356,N17357,N17358,
N17359,N17360,N17361,N17362,N17363,N17364,N17365,N17366,N17367,N17368,
N17369,N17370,N17371,N17372,N17373,N17374,N17375,N17376,N17377,N17378,
N17379,N17380,N17381,N17382,N17383,N17384,N17385,N17386,N17387,N17388,
N17389,N17390,N17391,N17392,N17393,N17394,N17395,N17396,N17397,N17398,
N17399,N17400,N17401,N17402,N17403,N17404,N17405,N17406,N17407,N17408,
N17409,N17410,N17411,N17412,N17413,N17414,N17415,N17416,N17417,N17418,
N17419,N17420,N17421,N17422,N17423,N17424,N17425,N17426,N17427,N17428,
N17429,N17430,N17431,N17432,N17433,N17434,N17435,N17436,N17437,N17438,
N17439,N17440,N17441,N17442,N17443,N17444,N17445,N17446,N17447,N17448,
N17449,N17450,N17451,N17452,N17453,N17454,N17455,N17456,N17457,N17458,
N17459,N17460,N17461,N17462,N17463,N17464,N17465,N17466,N17467,N17468,
N17469,N17470,N17471,N17472,N17473,N17474,N17475,N17476,N17477,N17478,
N17479,N17480,N17481,N17482,N17483,N17484,N17485,N17486,N17487,N17488,
N17489,N17490,N17491,N17492,N17493,N17494,N17495,N17496,N17497,N17498,
N17499,N17500,N17501,N17502,N17503,N17504,N17505,N17506,N17507,N17508,
N17509,N17510,N17511,N17512,N17513,N17514,N17515,N17516,N17517,N17518,
N17519,N17520,N17521,N17522,N17523,N17524,N17525,N17526,N17527,N17528,
N17529,N17530,N17531,N17532,N17533,N17534,N17535,N17536,N17537,N17538,
N17539,N17540,N17541,N17542,N17543,N17544,N17545,N17546,N17547,N17548,
N17549,N17550,N17551,N17552,N17553,N17554,N17555,N17556,N17557,N17558,
N17559,N17560,N17561,N17562,N17563,N17564,N17565,N17566,N17567,N17568,
N17569,N17570,N17571,N17572,N17573,N17574,N17575,N17576,N17577,N17578,
N17579,N17580,N17581,N17582,N17583,N17584,N17585,N17586,N17587,N17588,
N17589,N17590,N17591,N17592,N17593,N17594,N17595,N17596,N17597,N17598,
N17599,N17600,N17601,N17602,N17603,N17604,N17605,N17606,N17607,N17608,
N17609,N17610,N17611,N17612,N17613,N17614,N17615,N17616,N17617,N17618,
N17619,N17620,N17621,N17622,N17623,N17624,N17625,N17626,N17627,N17628,
N17629,N17630,N17631,N17632,N17633,N17634,N17635,N17636,N17637,N17638,
N17639,N17640,N17641,N17642,N17643,N17644,N17645,N17646,N17647,N17648,
N17649,N17650,N17651,N17652,N17653,N17654,N17655,N17656,N17657,N17658,
N17659,N17660,N17661,N17662,N17663,N17664,N17665,N17666,N17667,N17668,
N17669,N17670,N17671,N17672,N17673,N17674,N17675,N17676,N17677,N17678,
N17679,N17680,N17681,N17682,N17683,N17684,N17685,N17686,N17687,N17688,
N17689,N17690,N17691,N17692,N17693,N17694,N17695,N17696,N17697,N17698,
N17699,N17700,N17701,N17702,N17703,N17704,N17705,N17706,N17707,N17708,
N17709,N17710,N17711,N17712,N17713,N17714,N17715,N17716,N17717,N17718,
N17719,N17720,N17721,N17722,N17723,N17724,N17725,N17726,N17727,N17728,
N17729,N17730,N17731,N17732,N17733,N17734,N17735,N17736,N17737,N17738,
N17739,N17740,N17741,N17742,N17743,N17744,N17745,N17746,N17747,N17748,
N17749,N17750,N17751,N17752,N17753,N17754,N17755,N17756,N17757,N17758,
N17759,N17760,N17761,N17762,N17763,N17764,N17765,N17766,N17767,N17768,
N17769,N17770,N17771,N17772,N17773,N17774,N17775,N17776,N17777,N17778,
N17779,N17780,N17781,N17782,N17783,N17784,N17785,N17786,N17787,N17788,
N17789,N17790,N17791,N17792,N17793,N17794,N17795,N17796,N17797,N17798,
N17799,N17800,N17801,N17802,N17803,N17804,N17805,N17806,N17807,N17808,
N17809,N17810,N17811,N17812,N17813,N17814,N17815,N17816,N17817,N17818,
N17819,N17820,N17821,N17822,N17823,N17824,N17825,N17826,N17827,N17828,
N17829,N17830,N17831,N17832,N17833,N17834,N17835,N17836,N17837,N17838,
N17839,N17840,N17841,N17842,N17843,N17844,N17845,N17846,N17847,N17848,
N17849,N17850,N17851,N17852,N17853,N17854,N17855,N17856,N17857,N17858,
N17859,N17860,N17861,N17862,N17863,N17864,N17865,N17866,N17867,N17868,
N17869,N17870,N17871,N17872,N17873,N17874,N17875,N17876,N17877,N17878,
N17879,N17880,N17881,N17882,N17883,N17884,N17885,N17886,N17887,N17888,
N17889,N17890,N17891,N17892,N17893,N17894,N17895,N17896,N17897,N17898,
N17899,N17900,N17901,N17902,N17903,N17904,N17905,N17906,N17907,N17908,
N17909,N17910,N17911,N17912,N17913,N17914,N17915,N17916,N17917,N17918,
N17919,N17920,N17921,N17922,N17923,N17924,N17925,N17926,N17927,N17928,
N17929,N17930,N17931,N17932,N17933,N17934,N17935,N17936,N17937,N17938,
N17939,N17940,N17941,N17942,N17943,N17944,N17945,N17946,N17947,N17948,
N17949,N17950,N17951,N17952,N17953,N17954,N17955,N17956,N17957,N17958,
N17959,N17960,N17961,N17962,N17963,N17964,N17965,N17966,N17967,N17968,
N17969,N17970,N17971,N17972,N17973,N17974,N17975,N17976,N17977,N17978,
N17979,N17980,N17981,N17982,N17983,N17984,N17985,N17986,N17987,N17988,
N17989,N17990,N17991,N17992,N17993,N17994,N17995,N17996,N17997,N17998,
N17999,N18000,N18001,N18002,N18003,N18004,N18005,N18006,N18007,N18008,
N18009,N18010,N18011,N18012,N18013,N18014,N18015,N18016,N18017,N18018,
N18019,N18020,N18021,N18022,N18023,N18024,N18025,N18026,N18027,N18028,
N18029,N18030,N18031,N18032,N18033,N18034,N18035,N18036,N18037,N18038,
N18039,N18040,N18041,N18042,N18043,N18044,N18045,N18046,N18047,N18048,
N18049,N18050,N18051,N18052,N18053,N18054,N18055,N18056,N18057,N18058,
N18059,N18060,N18061,N18062,N18063,N18064,N18065,N18066,N18067,N18068,
N18069,N18070,N18071,N18072,N18073,N18074,N18075,N18076,N18077,N18078,
N18079,N18080,N18081,N18082,N18083,N18084,N18085,N18086,N18087,N18088,
N18089,N18090,N18091,N18092,N18093,N18094,N18095,N18096,N18097,N18098,
N18099,N18100,N18101,N18102,N18103,N18104,N18105,N18106,N18107,N18108,
N18109,N18110,N18111,N18112,N18113,N18114,N18115,N18116,N18117,N18118,
N18119,N18120,N18121,N18122,N18123,N18124,N18125,N18126,N18127,N18128,
N18129,N18130,N18131,N18132,N18133,N18134,N18135,N18136,N18137,N18138,
N18139,N18140,N18141,N18142,N18143,N18144,N18145,N18146,N18147,N18148,
N18149,N18150,N18151,N18152,N18153,N18154,N18155,N18156,N18157,N18158,
N18159,N18160,N18161,N18162,N18163,N18164,N18165,N18166,N18167,N18168,
N18169,N18170,N18171,N18172,N18173,N18174,N18175,N18176,N18177,N18178,
N18179,N18180,N18181,N18182,N18183,N18184,N18185,N18186,N18187,N18188,
N18189,N18190,N18191,N18192,N18193,N18194,N18195,N18196,N18197,N18198,
N18199,N18200,N18201,N18202,N18203,N18204,N18205,N18206,N18207,N18208,
N18209,N18210,N18211,N18212,N18213,N18214,N18215,N18216,N18217,N18218,
N18219,N18220,N18221,N18222,N18223,N18224,N18225,N18226,N18227,N18228,
N18229,N18230,N18231,N18232,N18233,N18234,N18235,N18236,N18237,N18238,
N18239,N18240,N18241,N18242,N18243,N18244,N18245,N18246,N18247,N18248,
N18249,N18250,N18251,N18252,N18253,N18254,N18255,N18256,N18257,N18258,
N18259,N18260,N18261,N18262,N18263,N18264,N18265,N18266,N18267,N18268,
N18269,N18270,N18271,N18272,N18273,N18274,N18275,N18276,N18277,N18278,
N18279,N18280,N18281,N18282,N18283,N18284,N18285,N18286,N18287,N18288,
N18289,N18290,N18291,N18292,N18293,N18294,N18295,N18296,N18297,N18298,
N18299,N18300,N18301,N18302,N18303,N18304,N18305,N18306,N18307,N18308,
N18309,N18310,N18311,N18312,N18313,N18314,N18315,N18316,N18317,N18318,
N18319,N18320,N18321,N18322,N18323,N18324,N18325,N18326,N18327,N18328,
N18329,N18330,N18331,N18332,N18333,N18334,N18335,N18336,N18337,N18338,
N18339,N18340,N18341,N18342,N18343,N18344,N18345,N18346,N18347,N18348,
N18349,N18350,N18351,N18352,N18353,N18354,N18355,N18356,N18357,N18358,
N18359,N18360,N18361,N18362,N18363,N18364,N18365,N18366,N18367,N18368,
N18369,N18370,N18371,N18372,N18373,N18374,N18375,N18376,N18377,N18378,
N18379,N18380,N18381,N18382,N18383,N18384,N18385,N18386,N18387,N18388,
N18389,N18390,N18391,N18392,N18393,N18394,N18395,N18396,N18397,N18398,
N18399,N18400,N18401,N18402,N18403,N18404,N18405,N18406,N18407,N18408,
N18409,N18410,N18411,N18412,N18413,N18414,N18415,N18416,N18417,N18418,
N18419,N18420,N18421,N18422,N18423,N18424,N18425,N18426,N18427,N18428,
N18429,N18430,N18431,N18432,N18433,N18434,N18435,N18436,N18437,N18438,
N18439,N18440,N18441,N18442,N18443,N18444,N18445,N18446,N18447,N18448,
N18449,N18450,N18451,N18452,N18453,N18454,N18455,N18456,N18457,N18458,
N18459,N18460,N18461,N18462,N18463,N18464,N18465,N18466,N18467,N18468,
N18469,N18470,N18471,N18472,N18473,N18474,N18475,N18476,N18477,N18478,
N18479,N18480,N18481,N18482,N18483,N18484,N18485,N18486,N18487,N18488,
N18489,N18490,N18491,N18492,N18493,N18494,N18495,N18496,N18497,N18498,
N18499,N18500,N18501,N18502,N18503,N18504,N18505,N18506,N18507,N18508,
N18509,N18510,N18511,N18512,N18513,N18514,N18515,N18516,N18517,N18518,
N18519,N18520,N18521,N18522,N18523,N18524,N18525,N18526,N18527,N18528,
N18529,N18530,N18531,N18532,N18533,N18534,N18535,N18536,N18537,N18538,
N18539,N18540,N18541,N18542,N18543,N18544,N18545,N18546,N18547,N18548,
N18549,N18550,N18551,N18552,N18553,N18554,N18555,N18556,N18557,N18558,
N18559,N18560,N18561,N18562,N18563,N18564,N18565,N18566,N18567,N18568,
N18569,N18570,N18571,N18572,N18573,N18574,N18575,N18576,N18577,N18578,
N18579,N18580,N18581,N18582,N18583,N18584,N18585,N18586,N18587,N18588,
N18589,N18590,N18591,N18592,N18593,N18594,N18595,N18596,N18597,N18598,
N18599,N18600,N18601,N18602,N18603,N18604,N18605,N18606,N18607,N18608,
N18609,N18610,N18611,N18612,N18613,N18614,N18615,N18616,N18617,N18618,
N18619,N18620,N18621,N18622,N18623,N18624,N18625,N18626,N18627,N18628,
N18629,N18630,N18631,N18632,N18633,N18634,N18635,N18636,N18637,N18638,
N18639,N18640,N18641,N18642,N18643,N18644,N18645,N18646,N18647,N18648,
N18649,N18650,N18651,N18652,N18653,N18654,N18655,N18656,N18657,N18658,
N18659,N18660,N18661,N18662,N18663,N18664,N18665,N18666,N18667,N18668,
N18669,N18670,N18671,N18672,N18673,N18674,N18675,N18676,N18677,N18678,
N18679,N18680,N18681,N18682,N18683,N18684,N18685,N18686,N18687,N18688,
N18689,N18690,N18691,N18692,N18693,N18694,N18695,N18696,N18697,N18698,
N18699,N18700,N18701,N18702,N18703,N18704,N18705,N18706,N18707,N18708,
N18709,N18710,N18711,N18712,N18713,N18714,N18715,N18716,N18717,N18718,
N18719,N18720,N18721,N18722,N18723,N18724,N18725,N18726,N18727,N18728,
N18729,N18730,N18731,N18732,N18733,N18734,N18735,N18736,N18737,N18738,
N18739,N18740,N18741,N18742,N18743,N18744,N18745,N18746,N18747,N18748,
N18749,N18750,N18751,N18752,N18753,N18754,N18755,N18756,N18757,N18758,
N18759,N18760,N18761,N18762,N18763,N18764,N18765,N18766,N18767,N18768,
N18769,N18770,N18771,N18772,N18773,N18774,N18775,N18776,N18777,N18778,
N18779,N18780,N18781,N18782,N18783,N18784,N18785,N18786,N18787,N18788,
N18789,N18790,N18791,N18792,N18793,N18794,N18795,N18796,N18797,N18798,
N18799,N18800,N18801,N18802,N18803,N18804,N18805,N18806,N18807,N18808,
N18809,N18810,N18811,N18812,N18813,N18814,N18815,N18816,N18817,N18818,
N18819,N18820,N18821,N18822,N18823,N18824,N18825,N18826,N18827,N18828,
N18829,N18830,N18831,N18832,N18833,N18834,N18835,N18836,N18837,N18838,
N18839,N18840,N18841,N18842,N18843,N18844,N18845,N18846,N18847,N18848,
N18849,N18850,N18851,N18852,N18853,N18854,N18855,N18856,N18857,N18858,
N18859,N18860,N18861,N18862,N18863,N18864,N18865,N18866,N18867,N18868,
N18869,N18870,N18871,N18872,N18873,N18874,N18875,N18876,N18877,N18878,
N18879,N18880,N18881,N18882,N18883,N18884,N18885,N18886,N18887,N18888,
N18889,N18890,N18891,N18892,N18893,N18894,N18895,N18896,N18897,N18898,
N18899,N18900,N18901,N18902,N18903,N18904,N18905,N18906,N18907,N18908,
N18909,N18910,N18911,N18912,N18913,N18914,N18915,N18916,N18917,N18918,
N18919,N18920,N18921,N18922,N18923,N18924,N18925,N18926,N18927,N18928,
N18929,N18930,N18931,N18932,N18933,N18934,N18935,N18936,N18937,N18938,
N18939,N18940,N18941,N18942,N18943,N18944,N18945,N18946,N18947,N18948,
N18949,N18950,N18951,N18952,N18953,N18954,N18955,N18956,N18957,N18958,
N18959,N18960,N18961,N18962,N18963,N18964,N18965,N18966,N18967,N18968,
N18969,N18970,N18971,N18972,N18973,N18974,N18975,N18976,N18977,N18978,
N18979,N18980,N18981,N18982,N18983,N18984,N18985,N18986,N18987,N18988,
N18989,N18990,N18991,N18992,N18993,N18994,N18995,N18996,N18997,N18998,
N18999,N19000,N19001,N19002,N19003,N19004,N19005,N19006,N19007,N19008,
N19009,N19010,N19011,N19012,N19013,N19014,N19015,N19016,N19017,N19018,
N19019,N19020,N19021,N19022,N19023,N19024,N19025,N19026,N19027,N19028,
N19029,N19030,N19031,N19032,N19033,N19034,N19035,N19036,N19037,N19038,
N19039,N19040,N19041,N19042,N19043,N19044,N19045,N19046,N19047,N19048,
N19049,N19050,N19051,N19052,N19053,N19054,N19055,N19056,N19057,N19058,
N19059,N19060,N19061,N19062,N19063,N19064,N19065,N19066,N19067,N19068,
N19069,N19070,N19071,N19072,N19073,N19074,N19075,N19076,N19077,N19078,
N19079,N19080,N19081,N19082,N19083,N19084,N19085,N19086,N19087,N19088,
N19089,N19090,N19091,N19092,N19093,N19094,N19095,N19096,N19097,N19098,
N19099,N19100,N19101,N19102,N19103,N19104,N19105,N19106,N19107,N19108,
N19109,N19110,N19111,N19112,N19113,N19114,N19115,N19116,N19117,N19118,
N19119,N19120,N19121,N19122,N19123,N19124,N19125,N19126,N19127,N19128,
N19129,N19130,N19131,N19132,N19133,N19134,N19135,N19136,N19137,N19138,
N19139,N19140,N19141,N19142,N19143,N19144,N19145,N19146,N19147,N19148,
N19149,N19150,N19151,N19152,N19153,N19154,N19155,N19156,N19157,N19158,
N19159,N19160,N19161,N19162,N19163,N19164,N19165,N19166,N19167,N19168,
N19169,N19170,N19171,N19172,N19173,N19174,N19175,N19176,N19177,N19178,
N19179,N19180,N19181,N19182,N19183,N19184,N19185,N19186,N19187,N19188,
N19189,N19190,N19191,N19192,N19193,N19194,N19195,N19196,N19197,N19198,
N19199,N19200,N19201,N19202,N19203,N19204,N19205,N19206,N19207,N19208,
N19209,N19210,N19211,N19212,N19213,N19214,N19215,N19216,N19217,N19218,
N19219,N19220,N19221,N19222,N19223,N19224,N19225,N19226,N19227,N19228,
N19229,N19230,N19231,N19232,N19233,N19234,N19235,N19236,N19237,N19238,
N19239,N19240,N19241,N19242,N19243,N19244,N19245,N19246,N19247,N19248,
N19249,N19250,N19251,N19252,N19253,N19254,N19255,N19256,N19257,N19258,
N19259,N19260,N19261,N19262,N19263,N19264,N19265,N19266,N19267,N19268,
N19269,N19270,N19271,N19272,N19273,N19274,N19275,N19276,N19277,N19278,
N19279,N19280,N19281,N19282,N19283,N19284,N19285,N19286,N19287,N19288,
N19289,N19290,N19291,N19292,N19293,N19294,N19295,N19296,N19297,N19298,
N19299,N19300,N19301,N19302,N19303,N19304,N19305,N19306,N19307,N19308,
N19309,N19310,N19311,N19312,N19313,N19314,N19315,N19316,N19317,N19318,
N19319,N19320,N19321,N19322,N19323,N19324,N19325,N19326,N19327,N19328,
N19329,N19330,N19331,N19332,N19333,N19334,N19335,N19336,N19337,N19338,
N19339,N19340,N19341,N19342,N19343,N19344,N19345,N19346,N19347,N19348,
N19349,N19350,N19351,N19352,N19353,N19354,N19355,N19356,N19357,N19358,
N19359,N19360,N19361,N19362,N19363,N19364,N19365,N19366,N19367,N19368,
N19369,N19370,N19371,N19372,N19373,N19374,N19375,N19376,N19377,N19378,
N19379,N19380,N19381,N19382,N19383,N19384,N19385,N19386,N19387,N19388,
N19389,N19390,N19391,N19392,N19393,N19394,N19395,N19396,N19397,N19398,
N19399,N19400,N19401,N19402,N19403,N19404,N19405,N19406,N19407,N19408,
N19409,N19410,N19411,N19412,N19413,N19414,N19415,N19416,N19417,N19418,
N19419,N19420,N19421,N19422,N19423,N19424,N19425,N19426,N19427,N19428,
N19429,N19430,N19431,N19432,N19433,N19434,N19435,N19436,N19437,N19438,
N19439,N19440,N19441,N19442,N19443,N19444,N19445,N19446,N19447,N19448,
N19449,N19450,N19451,N19452,N19453,N19454,N19455,N19456,N19457,N19458,
N19459,N19460,N19461,N19462,N19463,N19464,N19465,N19466,N19467,N19468,
N19469,N19470,N19471,N19472,N19473,N19474,N19475,N19476,N19477,N19478,
N19479,N19480,N19481,N19482,N19483,N19484,N19485,N19486,N19487,N19488,
N19489,N19490,N19491,N19492,N19493,N19494,N19495,N19496,N19497,N19498,
N19499,N19500,N19501,N19502,N19503,N19504,N19505,N19506,N19507,N19508,
N19509,N19510,N19511,N19512,N19513,N19514,N19515,N19516,N19517,N19518,
N19519,N19520,N19521,N19522,N19523,N19524,N19525,N19526,N19527,N19528,
N19529,N19530,N19531,N19532,N19533,N19534,N19535,N19536,N19537,N19538,
N19539,N19540,N19541,N19542,N19543,N19544,N19545,N19546,N19547,N19548,
N19549,N19550,N19551,N19552,N19553,N19554,N19555,N19556,N19557,N19558,
N19559,N19560,N19561,N19562,N19563,N19564,N19565,N19566,N19567,N19568,
N19569,N19570,N19571,N19572,N19573,N19574,N19575,N19576,N19577,N19578,
N19579,N19580,N19581,N19582,N19583,N19584,N19585,N19586,N19587,N19588,
N19589,N19590,N19591,N19592,N19593,N19594,N19595,N19596,N19597,N19598,
N19599,N19600,N19601,N19602,N19603,N19604,N19605,N19606,N19607,N19608,
N19609,N19610,N19611,N19612,N19613,N19614,N19615,N19616,N19617,N19618,
N19619,N19620,N19621,N19622,N19623,N19624,N19625,N19626,N19627,N19628,
N19629,N19630,N19631,N19632,N19633,N19634,N19635,N19636,N19637,N19638,
N19639,N19640,N19641,N19642,N19643,N19644,N19645,N19646,N19647,N19648,
N19649,N19650,N19651,N19652,N19653,N19654,N19655,N19656,N19657,N19658,
N19659,N19660,N19661,N19662,N19663,N19664,N19665,N19666,N19667,N19668,
N19669,N19670,N19671,N19672,N19673,N19674,N19675,N19676,N19677,N19678,
N19679,N19680,N19681,N19682,N19683,N19684,N19685,N19686,N19687,N19688,
N19689,N19690,N19691,N19692,N19693,N19694,N19695,N19696,N19697,N19698,
N19699,N19700,N19701,N19702,N19703,N19704,N19705,N19706,N19707,N19708,
N19709,N19710,N19711,N19712,N19713,N19714,N19715,N19716,N19717,N19718,
N19719,N19720,N19721,N19722,N19723,N19724,N19725,N19726,N19727,N19728,
N19729,N19730,N19731,N19732,N19733,N19734,N19735,N19736,N19737,N19738,
N19739,N19740,N19741,N19742,N19743,N19744,N19745,N19746,N19747,N19748,
N19749,N19750,N19751,N19752,N19753,N19754,N19755,N19756,N19757,N19758,
N19759,N19760,N19761,N19762,N19763,N19764,N19765,N19766,N19767,N19768,
N19769,N19770,N19771,N19772,N19773,N19774,N19775,N19776,N19777,N19778,
N19779,N19780,N19781,N19782,N19783,N19784,N19785,N19786,N19787,N19788,
N19789,N19790,N19791,N19792,N19793,N19794,N19795,N19796,N19797,N19798,
N19799,N19800,N19801,N19802,N19803,N19804,N19805,N19806,N19807,N19808,
N19809,N19810,N19811,N19812,N19813,N19814,N19815,N19816,N19817,N19818,
N19819,N19820,N19821,N19822,N19823,N19824,N19825,N19826,N19827,N19828,
N19829,N19830,N19831,N19832,N19833,N19834,N19835,N19836,N19837,N19838,
N19839,N19840,N19841,N19842,N19843,N19844,N19845,N19846,N19847,N19848,
N19849,N19850,N19851,N19852,N19853,N19854,N19855,N19856,N19857,N19858,
N19859,N19860,N19861,N19862,N19863,N19864,N19865,N19866,N19867,N19868,
N19869,N19870,N19871,N19872,N19873,N19874,N19875,N19876,N19877,N19878,
N19879,N19880,N19881,N19882,N19883,N19884,N19885,N19886,N19887,N19888,
N19889,N19890,N19891,N19892,N19893,N19894,N19895,N19896,N19897,N19898,
N19899,N19900,N19901,N19902,N19903,N19904,N19905,N19906,N19907,N19908,
N19909,N19910,N19911,N19912,N19913,N19914,N19915,N19916,N19917,N19918,
N19919,N19920,N19921,N19922,N19923,N19924,N19925,N19926,N19927,N19928,
N19929,N19930,N19931,N19932,N19933,N19934,N19935,N19936,N19937,N19938,
N19939,N19940,N19941,N19942,N19943,N19944,N19945,N19946,N19947,N19948,
N19949,N19950,N19951,N19952,N19953,N19954,N19955,N19956,N19957,N19958,
N19959,N19960,N19961,N19962,N19963,N19964,N19965,N19966,N19967,N19968,
N19969,N19970,N19971,N19972,N19973,N19974,N19975,N19976,N19977,N19978,
N19979,N19980,N19981,N19982,N19983,N19984,N19985,N19986,N19987,N19988,
N19989,N19990,N19991,N19992,N19993,N19994,N19995,N19996,N19997,N19998,
N19999,N20000,N20001,N20002,N20003,N20004,N20005,N20006,N20007,N20008,
N20009,N20010,N20011,N20012,N20013,N20014,N20015,N20016,N20017,N20018,
N20019,N20020,N20021,N20022,N20023,N20024,N20025,N20026,N20027,N20028,
N20029,N20030,N20031,N20032,N20033,N20034,N20035,N20036,N20037,N20038,
N20039,N20040,N20041,N20042,N20043,N20044,N20045,N20046,N20047,N20048,
N20049,N20050,N20051,N20052,N20053,N20054,N20055,N20056,N20057,N20058,
N20059,N20060,N20061,N20062,N20063,N20064,N20065,N20066,N20067,N20068,
N20069,N20070,N20071,N20072,N20073,N20074,N20075,N20076,N20077,N20078,
N20079,N20080,N20081,N20082,N20083,N20084,N20085,N20086,N20087,N20088,
N20089,N20090,N20091,N20092,N20093,N20094,N20095,N20096,N20097,N20098,
N20099,N20100,N20101,N20102,N20103,N20104,N20105,N20106,N20107,N20108,
N20109,N20110,N20111,N20112,N20113,N20114,N20115,N20116,N20117,N20118,
N20119,N20120,N20121,N20122,N20123,N20124,N20125,N20126,N20127,N20128,
N20129,N20130,N20131,N20132,N20133,N20134,N20135,N20136,N20137,N20138,
N20139,N20140,N20141,N20142,N20143,N20144,N20145,N20146,N20147,N20148,
N20149,N20150,N20151,N20152,N20153,N20154,N20155,N20156,N20157,N20158,
N20159,N20160,N20161,N20162,N20163,N20164,N20165,N20166,N20167,N20168,
N20169,N20170,N20171,N20172,N20173,N20174,N20175,N20176,N20177,N20178,
N20179,N20180,N20181,N20182,N20183,N20184,N20185,N20186,N20187,N20188,
N20189,N20190,N20191,N20192,N20193,N20194,N20195,N20196,N20197,N20198,
N20199,N20200,N20201,N20202,N20203,N20204,N20205,N20206,N20207,N20208,
N20209,N20210,N20211,N20212,N20213,N20214,N20215,N20216,N20217,N20218,
N20219,N20220,N20221,N20222,N20223,N20224,N20225,N20226,N20227,N20228,
N20229,N20230,N20231,N20232,N20233,N20234,N20235,N20236,N20237,N20238,
N20239,N20240,N20241,N20242,N20243,N20244,N20245,N20246,N20247,N20248,
N20249,N20250,N20251,N20252,N20253,N20254,N20255,N20256,N20257,N20258,
N20259,N20260,N20261,N20262,N20263,N20264,N20265,N20266,N20267,N20268,
N20269,N20270,N20271,N20272,N20273,N20274,N20275,N20276,N20277,N20278,
N20279,N20280,N20281,N20282,N20283,N20284,N20285,N20286,N20287,N20288,
N20289,N20290,N20291,N20292,N20293,N20294,N20295,N20296,N20297,N20298,
N20299,N20300,N20301,N20302,N20303,N20304,N20305,N20306,N20307,N20308,
N20309,N20310,N20311,N20312,N20313,N20314,N20315,N20316,N20317,N20318,
N20319,N20320,N20321,N20322,N20323,N20324,N20325,N20326,N20327,N20328,
N20329,N20330,N20331,N20332,N20333,N20334,N20335,N20336,N20337,N20338,
N20339,N20340,N20341,N20342,N20343,N20344,N20345,N20346,N20347,N20348,
N20349,N20350,N20351,N20352,N20353,N20354,N20355,N20356,N20357,N20358,
N20359,N20360,N20361,N20362,N20363,N20364,N20365,N20366,N20367,N20368,
N20369,N20370,N20371,N20372,N20373,N20374,N20375,N20376,N20377,N20378,
N20379,N20380,N20381,N20382,N20383,N20384,N20385,N20386,N20387,N20388,
N20389,N20390,N20391,N20392,N20393,N20394,N20395,N20396,N20397,N20398,
N20399,N20400,N20401,N20402,N20403,N20404,N20405,N20406,N20407,N20408,
N20409,N20410,N20411,N20412,N20413,N20414,N20415,N20416,N20417,N20418,
N20419,N20420,N20421,N20422,N20423,N20424,N20425,N20426,N20427,N20428,
N20429,N20430,N20431,N20432,N20433,N20434,N20435,N20436,N20437,N20438,
N20439,N20440,N20441,N20442,N20443,N20444,N20445,N20446,N20447,N20448,
N20449,N20450,N20451,N20452,N20453,N20454,N20455,N20456,N20457,N20458,
N20459,N20460,N20461,N20462,N20463,N20464,N20465,N20466,N20467,N20468,
N20469,N20470,N20471,N20472,N20473,N20474,N20475,N20476,N20477,N20478,
N20479,N20480,N20481,N20482,N20483,N20484,N20485,N20486,N20487,N20488,
N20489,N20490,N20491,N20492,N20493,N20494,N20495,N20496,N20497,N20498,
N20499,N20500,N20501,N20502,N20503,N20504,N20505,N20506,N20507,N20508,
N20509,N20510,N20511,N20512,N20513,N20514,N20515,N20516,N20517,N20518,
N20519,N20520,N20521,N20522,N20523,N20524,N20525,N20526,N20527,N20528,
N20529,N20530,N20531,N20532,N20533,N20534,N20535,N20536,N20537,N20538,
N20539,N20540,N20541,N20542,N20543,N20544,N20545,N20546,N20547,N20548,
N20549,N20550,N20551,N20552,N20553,N20554,N20555,N20556,N20557,N20558,
N20559,N20560,N20561,N20562,N20563,N20564,N20565,N20566,N20567,N20568,
N20569,N20570,N20571,N20572,N20573,N20574,N20575,N20576,N20577,N20578,
N20579,N20580,N20581,N20582,N20583,N20584,N20585,N20586,N20587,N20588,
N20589,N20590,N20591,N20592,N20593,N20594,N20595,N20596,N20597,N20598,
N20599,N20600,N20601,N20602,N20603,N20604,N20605,N20606,N20607,N20608,
N20609,N20610,N20611,N20612,N20613,N20614,N20615,N20616,N20617,N20618,
N20619,N20620,N20621,N20622,N20623,N20624,N20625,N20626,N20627,N20628,
N20629,N20630,N20631,N20632,N20633,N20634,N20635,N20636,N20637,N20638,
N20639,N20640,N20641,N20642,N20643,N20644,N20645,N20646,N20647,N20648,
N20649,N20650,N20651,N20652,N20653,N20654,N20655,N20656,N20657,N20658,
N20659,N20660,N20661,N20662,N20663,N20664,N20665,N20666,N20667,N20668,
N20669,N20670,N20671,N20672,N20673,N20674,N20675,N20676,N20677,N20678,
N20679,N20680,N20681,N20682,N20683,N20684,N20685,N20686,N20687,N20688,
N20689,N20690,N20691,N20692,N20693,N20694,N20695,N20696,N20697,N20698,
N20699,N20700,N20701,N20702,N20703,N20704,N20705,N20706,N20707,N20708,
N20709,N20710,N20711,N20712,N20713,N20714,N20715,N20716,N20717,N20718,
N20719,N20720,N20721,N20722,N20723,N20724,N20725,N20726,N20727,N20728,
N20729,N20730,N20731,N20732,N20733,N20734,N20735,N20736,N20737,N20738,
N20739,N20740,N20741,N20742,N20743,N20744,N20745,N20746,N20747,N20748,
N20749,N20750,N20751,N20752,N20753,N20754,N20755,N20756,N20757,N20758,
N20759,N20760,N20761,N20762,N20763,N20764,N20765,N20766,N20767,N20768,
N20769,N20770,N20771,N20772,N20773,N20774,N20775,N20776,N20777,N20778,
N20779,N20780,N20781,N20782,N20783,N20784,N20785,N20786,N20787,N20788,
N20789,N20790,N20791,N20792,N20793,N20794,N20795,N20796,N20797,N20798,
N20799,N20800,N20801,N20802,N20803,N20804,N20805,N20806,N20807,N20808,
N20809,N20810,N20811,N20812,N20813,N20814,N20815,N20816,N20817,N20818,
N20819,N20820,N20821,N20822,N20823,N20824,N20825,N20826,N20827,N20828,
N20829,N20830,N20831,N20832,N20833,N20834,N20835,N20836,N20837,N20838,
N20839,N20840,N20841,N20842,N20843,N20844,N20845,N20846,N20847,N20848,
N20849,N20850,N20851,N20852,N20853,N20854,N20855,N20856,N20857,N20858,
N20859,N20860,N20861,N20862,N20863,N20864,N20865,N20866,N20867,N20868,
N20869,N20870,N20871,N20872,N20873,N20874,N20875,N20876,N20877,N20878,
N20879,N20880,N20881,N20882,N20883,N20884,N20885,N20886,N20887,N20888,
N20889,N20890,N20891,N20892,N20893,N20894,N20895,N20896,N20897,N20898,
N20899,N20900,N20901,N20902,N20903,N20904,N20905,N20906,N20907,N20908,
N20909,N20910,N20911,N20912,N20913,N20914,N20915,N20916,N20917,N20918,
N20919,N20920,N20921,N20922,N20923,N20924,N20925,N20926,N20927,N20928,
N20929,N20930,N20931,N20932,N20933,N20934,N20935,N20936,N20937,N20938,
N20939,N20940,N20941,N20942,N20943,N20944,N20945,N20946,N20947,N20948,
N20949,N20950,N20951,N20952,N20953,N20954,N20955,N20956,N20957,N20958,
N20959,N20960,N20961,N20962,N20963,N20964,N20965,N20966,N20967,N20968,
N20969,N20970,N20971,N20972,N20973,N20974,N20975,N20976,N20977,N20978,
N20979,N20980,N20981,N20982,N20983,N20984,N20985,N20986,N20987,N20988,
N20989,N20990,N20991,N20992,N20993,N20994,N20995,N20996,N20997,N20998,
N20999,N21000,N21001,N21002,N21003,N21004,N21005,N21006,N21007,N21008,
N21009,N21010,N21011,N21012,N21013,N21014,N21015,N21016,N21017,N21018,
N21019,N21020,N21021,N21022,N21023,N21024,N21025,N21026,N21027,N21028,
N21029,N21030,N21031,N21032,N21033,N21034,N21035,N21036,N21037,N21038,
N21039,N21040,N21041,N21042,N21043,N21044,N21045,N21046,N21047,N21048,
N21049,N21050,N21051,N21052,N21053,N21054,N21055,N21056,N21057,N21058,
N21059,N21060,N21061,N21062,N21063,N21064,N21065,N21066,N21067,N21068,
N21069,N21070,N21071,N21072,N21073,N21074,N21075,N21076,N21077,N21078,
N21079,N21080,N21081,N21082,N21083,N21084,N21085,N21086,N21087,N21088,
N21089,N21090,N21091,N21092,N21093,N21094,N21095,N21096,N21097,N21098,
N21099,N21100,N21101,N21102,N21103,N21104,N21105,N21106,N21107,N21108,
N21109,N21110,N21111,N21112,N21113,N21114,N21115,N21116,N21117,N21118,
N21119,N21120,N21121,N21122,N21123,N21124,N21125,N21126,N21127,N21128,
N21129,N21130,N21131,N21132,N21133,N21134,N21135,N21136,N21137,N21138,
N21139,N21140,N21141,N21142,N21143,N21144,N21145,N21146,N21147,N21148,
N21149,N21150,N21151,N21152,N21153,N21154,N21155,N21156,N21157,N21158,
N21159,N21160,N21161,N21162,N21163,N21164,N21165,N21166,N21167,N21168,
N21169,N21170,N21171,N21172,N21173,N21174,N21175,N21176,N21177,N21178,
N21179,N21180,N21181,N21182,N21183,N21184,N21185,N21186,N21187,N21188,
N21189,N21190,N21191,N21192,N21193,N21194,N21195,N21196,N21197,N21198,
N21199,N21200,N21201,N21202,N21203,N21204,N21205,N21206,N21207,N21208,
N21209,N21210,N21211,N21212,N21213,N21214,N21215,N21216,N21217,N21218,
N21219,N21220,N21221,N21222,N21223,N21224,N21225,N21226,N21227,N21228,
N21229,N21230,N21231,N21232,N21233,N21234,N21235,N21236,N21237,N21238,
N21239,N21240,N21241,N21242,N21243,N21244,N21245,N21246,N21247,N21248,
N21249,N21250,N21251,N21252,N21253,N21254,N21255,N21256,N21257,N21258,
N21259,N21260,N21261,N21262,N21263,N21264,N21265,N21266,N21267,N21268,
N21269,N21270,N21271,N21272,N21273,N21274,N21275,N21276,N21277,N21278,
N21279,N21280,N21281,N21282,N21283,N21284,N21285,N21286,N21287,N21288,
N21289,N21290,N21291,N21292,N21293,N21294,N21295,N21296,N21297,N21298,
N21299,N21300,N21301,N21302,N21303,N21304,N21305,N21306,N21307,N21308,
N21309,N21310,N21311,N21312,N21313,N21314,N21315,N21316,N21317,N21318,
N21319,N21320,N21321,N21322,N21323,N21324,N21325,N21326,N21327,N21328,
N21329,N21330,N21331,N21332,N21333,N21334,N21335,N21336,N21337,N21338,
N21339,N21340,N21341,N21342,N21343,N21344,N21345,N21346,N21347,N21348,
N21349,N21350,N21351,N21352,N21353,N21354,N21355,N21356,N21357,N21358,
N21359,N21360,N21361,N21362,N21363,N21364,N21365,N21366,N21367,N21368,
N21369,N21370,N21371,N21372,N21373,N21374,N21375,N21376,N21377,N21378,
N21379,N21380,N21381,N21382,N21383,N21384,N21385,N21386,N21387,N21388,
N21389,N21390,N21391,N21392,N21393,N21394,N21395,N21396,N21397,N21398,
N21399,N21400,N21401,N21402,N21403,N21404,N21405,N21406,N21407,N21408,
N21409,N21410,N21411,N21412,N21413,N21414,N21415,N21416,N21417,N21418,
N21419,N21420,N21421,N21422,N21423,N21424,N21425,N21426,N21427,N21428,
N21429,N21430,N21431,N21432,N21433,N21434,N21435,N21436,N21437,N21438,
N21439,N21440,N21441,N21442,N21443,N21444,N21445,N21446,N21447,N21448,
N21449,N21450,N21451,N21452,N21453,N21454,N21455,N21456,N21457,N21458,
N21459,N21460,N21461,N21462,N21463,N21464,N21465,N21466,N21467,N21468,
N21469,N21470,N21471,N21472,N21473,N21474,N21475,N21476,N21477,N21478,
N21479,N21480,N21481,N21482,N21483,N21484,N21485,N21486,N21487,N21488,
N21489,N21490,N21491,N21492,N21493,N21494,N21495,N21496,N21497,N21498,
N21499,N21500,N21501,N21502,N21503,N21504,N21505,N21506,N21507,N21508,
N21509,N21510,N21511,N21512,N21513,N21514,N21515,N21516,N21517,N21518,
N21519,N21520,N21521,N21522,N21523,N21524,N21525,N21526,N21527,N21528,
N21529,N21530,N21531,N21532,N21533,N21534,N21535,N21536,N21537,N21538,
N21539,N21540,N21541,N21542,N21543,N21544,N21545,N21546,N21547,N21548,
N21549,N21550,N21551,N21552,N21553,N21554,N21555,N21556,N21557,N21558,
N21559,N21560,N21561,N21562,N21563,N21564,N21565,N21566,N21567,N21568,
N21569,N21570,N21571,N21572,N21573,N21574,N21575,N21576,N21577,N21578,
N21579,N21580,N21581,N21582,N21583,N21584,N21585,N21586,N21587,N21588,
N21589,N21590,N21591,N21592,N21593,N21594,N21595,N21596,N21597,N21598,
N21599,N21600,N21601,N21602,N21603,N21604,N21605,N21606,N21607,N21608,
N21609,N21610,N21611,N21612,N21613,N21614,N21615,N21616,N21617,N21618,
N21619,N21620,N21621,N21622,N21623,N21624,N21625,N21626,N21627,N21628,
N21629,N21630,N21631,N21632,N21633,N21634,N21635,N21636,N21637,N21638,
N21639,N21640,N21641,N21642,N21643,N21644,N21645,N21646,N21647,N21648,
N21649,N21650,N21651,N21652,N21653,N21654,N21655,N21656,N21657,N21658,
N21659,N21660,N21661,N21662,N21663,N21664,N21665,N21666,N21667,N21668,
N21669,N21670,N21671,N21672,N21673,N21674,N21675,N21676,N21677,N21678,
N21679,N21680,N21681,N21682,N21683,N21684,N21685,N21686,N21687,N21688,
N21689,N21690,N21691,N21692,N21693,N21694,N21695,N21696,N21697,N21698,
N21699,N21700,N21701,N21702,N21703,N21704,N21705,N21706,N21707,N21708,
N21709,N21710,N21711,N21712,N21713,N21714,N21715,N21716,N21717,N21718,
N21719,N21720,N21721,N21722,N21723,N21724,N21725,N21726,N21727,N21728,
N21729,N21730,N21731,N21732,N21733,N21734,N21735,N21736,N21737,N21738,
N21739,N21740,N21741,N21742,N21743,N21744,N21745,N21746,N21747,N21748,
N21749,N21750,N21751,N21752,N21753,N21754,N21755,N21756,N21757,N21758,
N21759,N21760,N21761,N21762,N21763,N21764,N21765,N21766,N21767,N21768,
N21769,N21770,N21771,N21772,N21773,N21774,N21775,N21776,N21777,N21778,
N21779,N21780,N21781,N21782,N21783,N21784,N21785,N21786,N21787,N21788,
N21789,N21790,N21791,N21792,N21793,N21794,N21795,N21796,N21797,N21798,
N21799,N21800,N21801,N21802,N21803,N21804,N21805,N21806,N21807,N21808,
N21809,N21810,N21811,N21812,N21813,N21814,N21815,N21816,N21817,N21818,
N21819,N21820,N21821,N21822,N21823,N21824,N21825,N21826,N21827,N21828,
N21829,N21830,N21831,N21832,N21833,N21834,N21835,N21836,N21837,N21838,
N21839,N21840,N21841,N21842,N21843,N21844,N21845,N21846,N21847,N21848,
N21849,N21850,N21851,N21852,N21853,N21854,N21855,N21856,N21857,N21858,
N21859,N21860,N21861,N21862,N21863,N21864,N21865,N21866,N21867,N21868,
N21869,N21870,N21871,N21872,N21873,N21874,N21875,N21876,N21877,N21878,
N21879,N21880,N21881,N21882,N21883,N21884,N21885,N21886,N21887,N21888,
N21889,N21890,N21891,N21892,N21893,N21894,N21895,N21896,N21897,N21898,
N21899,N21900,N21901,N21902,N21903,N21904,N21905,N21906,N21907,N21908,
N21909,N21910,N21911,N21912,N21913,N21914,N21915,N21916,N21917,N21918,
N21919,N21920,N21921,N21922,N21923,N21924,N21925,N21926,N21927,N21928,
N21929,N21930,N21931,N21932,N21933,N21934,N21935,N21936,N21937,N21938,
N21939,N21940,N21941,N21942,N21943,N21944,N21945,N21946,N21947,N21948,
N21949,N21950,N21951,N21952,N21953,N21954,N21955,N21956,N21957,N21958,
N21959,N21960,N21961,N21962,N21963,N21964,N21965,N21966,N21967,N21968,
N21969,N21970,N21971,N21972,N21973,N21974,N21975,N21976,N21977,N21978,
N21979,N21980,N21981,N21982,N21983,N21984,N21985,N21986,N21987,N21988,
N21989,N21990,N21991,N21992,N21993,N21994,N21995,N21996,N21997,N21998,
N21999,N22000,N22001,N22002,N22003,N22004,N22005,N22006,N22007,N22008,
N22009,N22010,N22011,N22012,N22013,N22014,N22015,N22016,N22017,N22018,
N22019,N22020,N22021,N22022,N22023,N22024,N22025,N22026,N22027,N22028,
N22029,N22030,N22031,N22032,N22033,N22034,N22035,N22036,N22037,N22038,
N22039,N22040,N22041,N22042,N22043,N22044,N22045,N22046,N22047,N22048,
N22049,N22050,N22051,N22052,N22053,N22054,N22055,N22056,N22057,N22058,
N22059,N22060,N22061,N22062,N22063,N22064,N22065,N22066,N22067,N22068,
N22069,N22070,N22071,N22072,N22073,N22074,N22075,N22076,N22077,N22078,
N22079,N22080,N22081,N22082,N22083,N22084,N22085,N22086,N22087,N22088,
N22089,N22090,N22091,N22092,N22093,N22094,N22095,N22096,N22097,N22098,
N22099,N22100,N22101,N22102,N22103,N22104,N22105,N22106,N22107,N22108,
N22109,N22110,N22111,N22112,N22113,N22114,N22115,N22116,N22117,N22118,
N22119,N22120,N22121,N22122,N22123,N22124,N22125,N22126,N22127,N22128,
N22129,N22130,N22131,N22132,N22133,N22134,N22135,N22136,N22137,N22138,
N22139,N22140,N22141,N22142,N22143,N22144,N22145,N22146,N22147,N22148,
N22149,N22150,N22151,N22152,N22153,N22154,N22155,N22156,N22157,N22158,
N22159,N22160,N22161,N22162,N22163,N22164,N22165,N22166,N22167,N22168,
N22169,N22170,N22171,N22172,N22173,N22174,N22175,N22176,N22177,N22178,
N22179,N22180,N22181,N22182,N22183,N22184,N22185,N22186,N22187,N22188,
N22189,N22190,N22191,N22192,N22193,N22194,N22195,N22196,N22197,N22198,
N22199,N22200,N22201,N22202,N22203,N22204,N22205,N22206,N22207,N22208,
N22209,N22210,N22211,N22212,N22213,N22214,N22215,N22216,N22217,N22218,
N22219,N22220,N22221,N22222,N22223,N22224,N22225,N22226,N22227,N22228,
N22229,N22230,N22231,N22232,N22233,N22234,N22235,N22236,N22237,N22238,
N22239,N22240,N22241,N22242,N22243,N22244,N22245,N22246,N22247,N22248,
N22249,N22250,N22251,N22252,N22253,N22254,N22255,N22256,N22257,N22258,
N22259,N22260,N22261,N22262,N22263,N22264,N22265,N22266,N22267,N22268,
N22269,N22270,N22271,N22272,N22273,N22274,N22275,N22276,N22277,N22278,
N22279,N22280,N22281,N22282,N22283,N22284,N22285,N22286,N22287,N22288,
N22289,N22290,N22291,N22292,N22293,N22294,N22295,N22296,N22297,N22298,
N22299,N22300,N22301,N22302,N22303,N22304,N22305,N22306,N22307,N22308,
N22309,N22310,N22311,N22312,N22313,N22314,N22315,N22316,N22317,N22318,
N22319,N22320,N22321,N22322,N22323,N22324,N22325,N22326,N22327,N22328,
N22329,N22330,N22331,N22332,N22333,N22334,N22335,N22336,N22337,N22338,
N22339,N22340,N22341,N22342,N22343,N22344,N22345,N22346,N22347,N22348,
N22349,N22350,N22351,N22352,N22353,N22354,N22355,N22356,N22357,N22358,
N22359,N22360,N22361,N22362,N22363,N22364,N22365,N22366,N22367,N22368,
N22369,N22370,N22371,N22372,N22373,N22374,N22375,N22376,N22377,N22378,
N22379,N22380,N22381,N22382,N22383,N22384,N22385,N22386,N22387,N22388,
N22389,N22390,N22391,N22392,N22393,N22394,N22395,N22396,N22397,N22398,
N22399,N22400,N22401,N22402,N22403,N22404,N22405,N22406,N22407,N22408,
N22409,N22410,N22411,N22412,N22413,N22414,N22415,N22416,N22417,N22418,
N22419,N22420,N22421,N22422,N22423,N22424,N22425,N22426,N22427,N22428,
N22429,N22430,N22431,N22432,N22433,N22434,N22435,N22436,N22437,N22438,
N22439,N22440,N22441,N22442,N22443,N22444,N22445,N22446,N22447,N22448,
N22449,N22450,N22451,N22452,N22453,N22454,N22455,N22456,N22457,N22458,
N22459,N22460,N22461,N22462,N22463,N22464,N22465,N22466,N22467,N22468,
N22469,N22470,N22471,N22472,N22473,N22474,N22475,N22476,N22477,N22478,
N22479,N22480,N22481,N22482,N22483,N22484,N22485,N22486,N22487,N22488,
N22489,N22490,N22491,N22492,N22493,N22494,N22495,N22496,N22497,N22498,
N22499,N22500,N22501,N22502,N22503,N22504,N22505,N22506,N22507,N22508,
N22509,N22510,N22511,N22512,N22513,N22514,N22515,N22516,N22517,N22518,
N22519,N22520,N22521,N22522,N22523,N22524,N22525,N22526,N22527,N22528,
N22529,N22530,N22531,N22532,N22533,N22534,N22535,N22536,N22537,N22538,
N22539,N22540,N22541,N22542,N22543,N22544,N22545,N22546,N22547,N22548,
N22549,N22550,N22551,N22552,N22553,N22554,N22555,N22556,N22557,N22558,
N22559,N22560,N22561,N22562,N22563,N22564,N22565,N22566,N22567,N22568,
N22569,N22570,N22571,N22572,N22573,N22574,N22575,N22576,N22577,N22578,
N22579,N22580,N22581,N22582,N22583,N22584,N22585,N22586,N22587,N22588,
N22589,N22590,N22591,N22592,N22593,N22594,N22595,N22596,N22597,N22598,
N22599,N22600,N22601,N22602,N22603,N22604,N22605,N22606,N22607,N22608,
N22609,N22610,N22611,N22612,N22613,N22614,N22615,N22616,N22617,N22618,
N22619,N22620,N22621,N22622,N22623,N22624,N22625,N22626,N22627,N22628,
N22629,N22630,N22631,N22632,N22633,N22634,N22635,N22636,N22637,N22638,
N22639,N22640,N22641,N22642,N22643,N22644,N22645,N22646,N22647,N22648,
N22649,N22650,N22651,N22652,N22653,N22654,N22655,N22656,N22657,N22658,
N22659,N22660,N22661,N22662,N22663,N22664,N22665,N22666,N22667,N22668,
N22669,N22670,N22671,N22672,N22673,N22674,N22675,N22676,N22677,N22678,
N22679,N22680,N22681,N22682,N22683,N22684,N22685,N22686,N22687,N22688,
N22689,N22690,N22691,N22692,N22693,N22694,N22695,N22696,N22697,N22698,
N22699,N22700,N22701,N22702,N22703,N22704,N22705,N22706,N22707,N22708,
N22709,N22710,N22711,N22712,N22713,N22714,N22715,N22716,N22717,N22718,
N22719,N22720,N22721,N22722,N22723,N22724,N22725,N22726,N22727,N22728,
N22729,N22730,N22731,N22732,N22733,N22734,N22735,N22736,N22737,N22738,
N22739,N22740,N22741,N22742,N22743,N22744,N22745,N22746,N22747,N22748,
N22749,N22750,N22751,N22752,N22753,N22754,N22755,N22756,N22757,N22758,
N22759,N22760,N22761,N22762,N22763,N22764,N22765,N22766,N22767,N22768,
N22769,N22770,N22771,N22772,N22773,N22774,N22775,N22776,N22777,N22778,
N22779,N22780,N22781,N22782,N22783,N22784,N22785,N22786,N22787,N22788,
N22789,N22790,N22791,N22792,N22793,N22794,N22795,N22796,N22797,N22798,
N22799,N22800,N22801,N22802,N22803,N22804,N22805,N22806,N22807,N22808,
N22809,N22810,N22811,N22812,N22813,N22814,N22815,N22816,N22817,N22818,
N22819,N22820,N22821,N22822,N22823,N22824,N22825,N22826,N22827,N22828,
N22829,N22830,N22831,N22832,N22833,N22834,N22835,N22836,N22837,N22838,
N22839,N22840,N22841,N22842,N22843,N22844,N22845,N22846,N22847,N22848,
N22849,N22850,N22851,N22852,N22853,N22854,N22855,N22856,N22857,N22858,
N22859,N22860,N22861,N22862,N22863,N22864,N22865,N22866,N22867,N22868,
N22869,N22870,N22871,N22872,N22873,N22874,N22875,N22876,N22877,N22878,
N22879,N22880,N22881,N22882,N22883,N22884,N22885,N22886,N22887,N22888,
N22889,N22890,N22891,N22892,N22893,N22894,N22895,N22896,N22897,N22898,
N22899,N22900,N22901,N22902,N22903,N22904,N22905,N22906,N22907,N22908,
N22909,N22910,N22911,N22912,N22913,N22914,N22915,N22916,N22917,N22918,
N22919,N22920,N22921,N22922,N22923,N22924,N22925,N22926,N22927,N22928,
N22929,N22930,N22931,N22932,N22933,N22934,N22935,N22936,N22937,N22938,
N22939,N22940,N22941,N22942,N22943,N22944,N22945,N22946,N22947,N22948,
N22949,N22950,N22951,N22952,N22953,N22954,N22955,N22956,N22957,N22958,
N22959,N22960,N22961,N22962,N22963,N22964,N22965,N22966,N22967,N22968,
N22969,N22970,N22971,N22972,N22973,N22974,N22975,N22976,N22977,N22978,
N22979,N22980,N22981,N22982,N22983,N22984,N22985,N22986,N22987,N22988,
N22989,N22990,N22991,N22992,N22993,N22994,N22995,N22996,N22997,N22998,
N22999,N23000,N23001,N23002,N23003,N23004,N23005,N23006,N23007,N23008,
N23009,N23010,N23011,N23012,N23013,N23014,N23015,N23016,N23017,N23018,
N23019,N23020,N23021,N23022,N23023,N23024,N23025,N23026,N23027,N23028,
N23029,N23030,N23031,N23032,N23033,N23034,N23035,N23036,N23037,N23038,
N23039,N23040,N23041,N23042,N23043,N23044,N23045,N23046,N23047,N23048,
N23049,N23050,N23051,N23052,N23053,N23054,N23055,N23056,N23057,N23058,
N23059,N23060,N23061,N23062,N23063,N23064,N23065,N23066,N23067,N23068,
N23069,N23070,N23071,N23072,N23073,N23074,N23075,N23076,N23077,N23078,
N23079,N23080,N23081,N23082,N23083,N23084,N23085,N23086,N23087,N23088,
N23089,N23090,N23091,N23092,N23093,N23094,N23095,N23096,N23097,N23098,
N23099,N23100,N23101,N23102,N23103,N23104,N23105,N23106,N23107,N23108,
N23109,N23110,N23111,N23112,N23113,N23114,N23115,N23116,N23117,N23118,
N23119,N23120,N23121,N23122,N23123,N23124,N23125,N23126,N23127,N23128,
N23129,N23130,N23131,N23132,N23133,N23134,N23135,N23136,N23137,N23138,
N23139,N23140,N23141,N23142,N23143,N23144,N23145,N23146,N23147,N23148,
N23149,N23150,N23151,N23152,N23153,N23154,N23155,N23156,N23157,N23158,
N23159,N23160,N23161,N23162,N23163,N23164,N23165,N23166,N23167,N23168,
N23169,N23170,N23171,N23172,N23173,N23174,N23175,N23176,N23177,N23178,
N23179,N23180,N23181,N23182,N23183,N23184,N23185,N23186,N23187,N23188,
N23189,N23190,N23191,N23192,N23193,N23194,N23195,N23196,N23197,N23198,
N23199,N23200,N23201,N23202,N23203,N23204,N23205,N23206,N23207,N23208,
N23209,N23210,N23211,N23212,N23213,N23214,N23215,N23216,N23217,N23218,
N23219,N23220,N23221,N23222,N23223,N23224,N23225,N23226,N23227,N23228,
N23229,N23230,N23231,N23232,N23233,N23234,N23235,N23236,N23237,N23238,
N23239,N23240,N23241,N23242,N23243,N23244,N23245,N23246,N23247,N23248,
N23249,N23250,N23251,N23252,N23253,N23254,N23255,N23256,N23257,N23258,
N23259,N23260,N23261,N23262,N23263,N23264,N23265,N23266,N23267,N23268,
N23269,N23270,N23271,N23272,N23273,N23274,N23275,N23276,N23277,N23278,
N23279,N23280,N23281,N23282,N23283,N23284,N23285,N23286,N23287,N23288,
N23289,N23290,N23291,N23292,N23293,N23294,N23295,N23296,N23297,N23298,
N23299,N23300,N23301,N23302,N23303,N23304,N23305,N23306,N23307,N23308,
N23309,N23310,N23311,N23312,N23313,N23314,N23315,N23316,N23317,N23318,
N23319,N23320,N23321,N23322,N23323,N23324,N23325,N23326,N23327,N23328,
N23329,N23330,N23331,N23332,N23333,N23334,N23335,N23336,N23337,N23338,
N23339,N23340,N23341,N23342,N23343,N23344,N23345,N23346,N23347,N23348,
N23349,N23350,N23351,N23352,N23353,N23354,N23355,N23356,N23357,N23358,
N23359,N23360,N23361,N23362,N23363,N23364,N23365,N23366,N23367,N23368,
N23369,N23370,N23371,N23372,N23373,N23374,N23375,N23376,N23377,N23378,
N23379,N23380,N23381,N23382,N23383,N23384,N23385,N23386,N23387,N23388,
N23389,N23390,N23391,N23392,N23393,N23394,N23395,N23396,N23397,N23398,
N23399,N23400,N23401,N23402,N23403,N23404,N23405,N23406,N23407,N23408,
N23409,N23410,N23411,N23412,N23413,N23414,N23415,N23416,N23417,N23418,
N23419,N23420,N23421,N23422,N23423,N23424,N23425,N23426,N23427,N23428,
N23429,N23430,N23431,N23432,N23433,N23434,N23435,N23436,N23437,N23438,
N23439,N23440,N23441,N23442,N23443,N23444,N23445,N23446,N23447,N23448,
N23449,N23450,N23451,N23452,N23453,N23454,N23455,N23456,N23457,N23458,
N23459,N23460,N23461,N23462,N23463,N23464,N23465,N23466,N23467,N23468,
N23469,N23470,N23471,N23472,N23473,N23474,N23475,N23476,N23477,N23478,
N23479,N23480,N23481,N23482,N23483,N23484,N23485,N23486,N23487,N23488,
N23489,N23490,N23491,N23492,N23493,N23494,N23495,N23496,N23497,N23498,
N23499,N23500,N23501,N23502,N23503,N23504,N23505,N23506,N23507,N23508,
N23509,N23510,N23511,N23512,N23513,N23514,N23515,N23516,N23517,N23518,
N23519,N23520,N23521,N23522,N23523,N23524,N23525,N23526,N23527,N23528,
N23529,N23530,N23531,N23532,N23533,N23534,N23535,N23536,N23537,N23538,
N23539,N23540,N23541,N23542,N23543,N23544,N23545,N23546,N23547,N23548,
N23549,N23550,N23551,N23552,N23553,N23554,N23555,N23556,N23557,N23558,
N23559,N23560,N23561,N23562,N23563,N23564,N23565,N23566,N23567,N23568,
N23569,N23570,N23571,N23572,N23573,N23574,N23575,N23576,N23577,N23578,
N23579,N23580,N23581,N23582,N23583,N23584,N23585,N23586,N23587,N23588,
N23589,N23590,N23591,N23592,N23593,N23594,N23595,N23596,N23597,N23598,
N23599,N23600,N23601,N23602,N23603,N23604,N23605,N23606,N23607,N23608,
N23609,N23610,N23611,N23612,N23613,N23614,N23615,N23616,N23617,N23618,
N23619,N23620,N23621,N23622,N23623,N23624,N23625,N23626,N23627,N23628,
N23629,N23630,N23631,N23632,N23633,N23634,N23635,N23636,N23637,N23638,
N23639,N23640,N23641,N23642,N23643,N23644,N23645,N23646,N23647,N23648,
N23649,N23650,N23651,N23652,N23653,N23654,N23655,N23656,N23657,N23658,
N23659,N23660,N23661,N23662,N23663,N23664,N23665,N23666,N23667,N23668,
N23669,N23670,N23671,N23672,N23673,N23674,N23675,N23676,N23677,N23678,
N23679,N23680,N23681,N23682,N23683,N23684,N23685,N23686,N23687,N23688,
N23689,N23690,N23691,N23692,N23693,N23694,N23695,N23696,N23697,N23698,
N23699,N23700,N23701,N23702,N23703,N23704,N23705,N23706,N23707,N23708,
N23709,N23710,N23711,N23712,N23713,N23714,N23715,N23716,N23717,N23718,
N23719,N23720,N23721,N23722,N23723,N23724,N23725,N23726,N23727,N23728,
N23729,N23730,N23731,N23732,N23733,N23734,N23735,N23736,N23737,N23738,
N23739,N23740,N23741,N23742,N23743,N23744,N23745,N23746,N23747,N23748,
N23749,N23750,N23751,N23752,N23753,N23754,N23755,N23756,N23757,N23758,
N23759,N23760,N23761,N23762,N23763,N23764,N23765,N23766,N23767,N23768,
N23769,N23770,N23771,N23772,N23773,N23774,N23775,N23776,N23777,N23778,
N23779,N23780,N23781,N23782,N23783,N23784,N23785,N23786,N23787,N23788,
N23789,N23790,N23791,N23792,N23793,N23794,N23795,N23796,N23797,N23798,
N23799,N23800,N23801,N23802,N23803,N23804,N23805,N23806,N23807,N23808,
N23809,N23810,N23811,N23812,N23813,N23814,N23815,N23816,N23817,N23818,
N23819,N23820,N23821,N23822,N23823,N23824,N23825,N23826,N23827,N23828,
N23829,N23830,N23831,N23832,N23833,N23834,N23835,N23836,N23837,N23838,
N23839,N23840,N23841,N23842,N23843,N23844,N23845,N23846,N23847,N23848,
N23849,N23850,N23851,N23852,N23853,N23854,N23855,N23856,N23857,N23858,
N23859,N23860,N23861,N23862,N23863,N23864,N23865,N23866,N23867,N23868,
N23869,N23870,N23871,N23872,N23873,N23874,N23875,N23876,N23877,N23878,
N23879,N23880,N23881,N23882,N23883,N23884,N23885,N23886,N23887,N23888,
N23889,N23890,N23891,N23892,N23893,N23894,N23895,N23896,N23897,N23898,
N23899,N23900,N23901,N23902,N23903,N23904,N23905,N23906,N23907,N23908,
N23909,N23910,N23911,N23912,N23913,N23914,N23915,N23916,N23917,N23918,
N23919,N23920,N23921,N23922,N23923,N23924,N23925,N23926,N23927,N23928,
N23929,N23930,N23931,N23932,N23933,N23934,N23935,N23936,N23937,N23938,
N23939,N23940,N23941,N23942,N23943,N23944,N23945,N23946,N23947,N23948,
N23949,N23950,N23951,N23952,N23953,N23954,N23955,N23956,N23957,N23958,
N23959,N23960,N23961,N23962,N23963,N23964,N23965,N23966,N23967,N23968,
N23969,N23970,N23971,N23972,N23973,N23974,N23975,N23976,N23977,N23978,
N23979,N23980,N23981,N23982,N23983,N23984,N23985,N23986,N23987,N23988,
N23989,N23990,N23991,N23992,N23993,N23994,N23995,N23996,N23997,N23998,
N23999,N24000,N24001,N24002,N24003,N24004,N24005,N24006,N24007,N24008,
N24009,N24010,N24011,N24012,N24013,N24014,N24015,N24016,N24017,N24018,
N24019,N24020,N24021,N24022,N24023,N24024,N24025,N24026,N24027,N24028,
N24029,N24030,N24031,N24032,N24033,N24034,N24035,N24036,N24037,N24038,
N24039,N24040,N24041,N24042,N24043,N24044,N24045,N24046,N24047,N24048,
N24049,N24050,N24051,N24052,N24053,N24054,N24055,N24056,N24057,N24058,
N24059,N24060,N24061,N24062,N24063,N24064,N24065,N24066,N24067,N24068,
N24069,N24070,N24071,N24072,N24073,N24074,N24075,N24076,N24077,N24078,
N24079,N24080,N24081,N24082,N24083,N24084,N24085,N24086,N24087,N24088,
N24089,N24090,N24091,N24092,N24093,N24094,N24095,N24096,N24097,N24098,
N24099,N24100,N24101,N24102,N24103,N24104,N24105,N24106,N24107,N24108,
N24109,N24110,N24111,N24112,N24113,N24114,N24115,N24116,N24117,N24118,
N24119,N24120,N24121,N24122,N24123,N24124,N24125,N24126,N24127,N24128,
N24129,N24130,N24131,N24132,N24133,N24134,N24135,N24136,N24137,N24138,
N24139,N24140,N24141,N24142,N24143,N24144,N24145,N24146,N24147,N24148,
N24149,N24150,N24151,N24152,N24153,N24154,N24155,N24156,N24157,N24158,
N24159,N24160,N24161,N24162,N24163,N24164,N24165,N24166,N24167,N24168,
N24169,N24170,N24171,N24172,N24173,N24174,N24175,N24176,N24177,N24178,
N24179,N24180,N24181,N24182,N24183,N24184,N24185,N24186,N24187,N24188,
N24189,N24190,N24191,N24192,N24193,N24194,N24195,N24196,N24197,N24198,
N24199,N24200,N24201,N24202,N24203,N24204,N24205,N24206,N24207,N24208,
N24209,N24210,N24211,N24212,N24213,N24214,N24215,N24216,N24217,N24218,
N24219,N24220,N24221,N24222,N24223,N24224,N24225,N24226,N24227,N24228,
N24229,N24230,N24231,N24232,N24233,N24234,N24235,N24236,N24237,N24238,
N24239,N24240,N24241,N24242,N24243,N24244,N24245,N24246,N24247,N24248,
N24249,N24250,N24251,N24252,N24253,N24254,N24255,N24256,N24257,N24258,
N24259,N24260,N24261,N24262,N24263,N24264,N24265,N24266,N24267,N24268,
N24269,N24270,N24271,N24272,N24273,N24274,N24275,N24276,N24277,N24278,
N24279,N24280,N24281,N24282,N24283,N24284,N24285,N24286,N24287,N24288,
N24289,N24290,N24291,N24292,N24293,N24294,N24295,N24296,N24297,N24298,
N24299,N24300,N24301,N24302,N24303,N24304,N24305,N24306,N24307,N24308,
N24309,N24310,N24311,N24312,N24313,N24314,N24315,N24316,N24317,N24318,
N24319,N24320,N24321,N24322,N24323,N24324,N24325,N24326,N24327,N24328,
N24329,N24330,N24331,N24332,N24333,N24334,N24335,N24336,N24337,N24338,
N24339,N24340,N24341,N24342,N24343,N24344,N24345,N24346,N24347,N24348,
N24349,N24350,N24351,N24352,N24353,N24354,N24355,N24356,N24357,N24358,
N24359,N24360,N24361,N24362,N24363,N24364,N24365,N24366,N24367,N24368,
N24369,N24370,N24371,N24372,N24373,N24374,N24375,N24376,N24377,N24378,
N24379,N24380,N24381,N24382,N24383,N24384,N24385,N24386,N24387,N24388,
N24389,N24390,N24391,N24392,N24393,N24394,N24395,N24396,N24397,N24398,
N24399,N24400,N24401,N24402,N24403,N24404,N24405,N24406,N24407,N24408,
N24409,N24410,N24411,N24412,N24413,N24414,N24415,N24416,N24417,N24418,
N24419,N24420,N24421,N24422,N24423,N24424,N24425,N24426,N24427,N24428,
N24429,N24430,N24431,N24432,N24433,N24434,N24435,N24436,N24437,N24438,
N24439,N24440,N24441,N24442,N24443,N24444,N24445,N24446,N24447,N24448,
N24449,N24450,N24451,N24452,N24453,N24454,N24455,N24456,N24457,N24458,
N24459,N24460,N24461,N24462,N24463,N24464,N24465,N24466,N24467,N24468,
N24469,N24470,N24471,N24472,N24473,N24474,N24475,N24476,N24477,N24478,
N24479,N24480,N24481,N24482,N24483,N24484,N24485,N24486,N24487,N24488,
N24489,N24490,N24491,N24492,N24493,N24494,N24495,N24496,N24497,N24498,
N24499,N24500,N24501,N24502,N24503,N24504,N24505,N24506,N24507,N24508,
N24509,N24510,N24511,N24512,N24513,N24514,N24515,N24516,N24517,N24518,
N24519,N24520,N24521,N24522,N24523,N24524,N24525,N24526,N24527,N24528,
N24529,N24530,N24531,N24532,N24533,N24534,N24535,N24536,N24537,N24538,
N24539,N24540,N24541,N24542,N24543,N24544,N24545,N24546,N24547,N24548,
N24549,N24550,N24551,N24552,N24553,N24554,N24555,N24556,N24557,N24558,
N24559,N24560,N24561,N24562,N24563,N24564,N24565,N24566,N24567,N24568,
N24569,N24570,N24571,N24572,N24573,N24574,N24575,N24576,N24577,N24578,
N24579,N24580,N24581,N24582,N24583,N24584,N24585,N24586,N24587,N24588,
N24589,N24590,N24591,N24592,N24593,N24594,N24595,N24596,N24597,N24598,
N24599,N24600,N24601,N24602,N24603,N24604,N24605,N24606,N24607,N24608,
N24609,N24610,N24611,N24612,N24613,N24614,N24615,N24616,N24617,N24618,
N24619,N24620,N24621,N24622,N24623,N24624,N24625,N24626,N24627,N24628,
N24629,N24630,N24631,N24632,N24633,N24634,N24635,N24636,N24637,N24638,
N24639,N24640,N24641,N24642,N24643,N24644,N24645,N24646,N24647,N24648,
N24649,N24650,N24651,N24652,N24653,N24654,N24655,N24656,N24657,N24658,
N24659,N24660,N24661,N24662,N24663,N24664,N24665,N24666,N24667,N24668,
N24669,N24670,N24671,N24672,N24673,N24674,N24675,N24676,N24677,N24678,
N24679,N24680,N24681,N24682,N24683,N24684,N24685,N24686,N24687,N24688,
N24689,N24690,N24691,N24692,N24693,N24694,N24695,N24696,N24697,N24698,
N24699,N24700,N24701,N24702,N24703,N24704,N24705,N24706,N24707,N24708,
N24709,N24710,N24711,N24712,N24713,N24714,N24715,N24716,N24717,N24718,
N24719,N24720,N24721,N24722,N24723,N24724,N24725,N24726,N24727,N24728,
N24729,N24730,N24731,N24732,N24733,N24734,N24735,N24736,N24737,N24738,
N24739,N24740,N24741,N24742,N24743,N24744,N24745,N24746,N24747,N24748,
N24749,N24750,N24751,N24752,N24753,N24754,N24755,N24756,N24757,N24758,
N24759,N24760,N24761,N24762,N24763,N24764,N24765,N24766,N24767,N24768,
N24769,N24770,N24771,N24772,N24773,N24774,N24775,N24776,N24777,N24778,
N24779,N24780,N24781,N24782,N24783,N24784,N24785,N24786,N24787,N24788,
N24789,N24790,N24791,N24792,N24793,N24794,N24795,N24796,N24797,N24798,
N24799,N24800,N24801,N24802,N24803,N24804,N24805,N24806,N24807,N24808,
N24809,N24810,N24811,N24812,N24813,N24814,N24815,N24816,N24817,N24818,
N24819,N24820,N24821,N24822,N24823,N24824,N24825,N24826,N24827,N24828,
N24829,N24830,N24831,N24832,N24833,N24834,N24835,N24836,N24837,N24838,
N24839,N24840,N24841,N24842,N24843,N24844,N24845,N24846,N24847,N24848,
N24849,N24850,N24851,N24852,N24853,N24854,N24855,N24856,N24857,N24858,
N24859,N24860,N24861,N24862,N24863,N24864,N24865,N24866,N24867,N24868,
N24869,N24870,N24871,N24872,N24873,N24874,N24875,N24876,N24877,N24878,
N24879,N24880,N24881,N24882,N24883,N24884,N24885,N24886,N24887,N24888,
N24889,N24890,N24891,N24892,N24893,N24894,N24895,N24896,N24897,N24898,
N24899,N24900,N24901,N24902,N24903,N24904,N24905,N24906,N24907,N24908,
N24909,N24910,N24911,N24912,N24913,N24914,N24915,N24916,N24917,N24918,
N24919,N24920,N24921,N24922,N24923,N24924,N24925,N24926,N24927,N24928,
N24929,N24930,N24931,N24932,N24933,N24934,N24935,N24936,N24937,N24938,
N24939,N24940,N24941,N24942,N24943,N24944,N24945,N24946,N24947,N24948,
N24949,N24950,N24951,N24952,N24953,N24954,N24955,N24956,N24957,N24958,
N24959,N24960,N24961,N24962,N24963,N24964,N24965,N24966,N24967,N24968,
N24969,N24970,N24971,N24972,N24973,N24974,N24975,N24976,N24977,N24978,
N24979,N24980,N24981,N24982,N24983,N24984,N24985,N24986,N24987,N24988,
N24989,N24990,N24991,N24992,N24993,N24994,N24995,N24996,N24997,N24998,
N24999,N25000,N25001,N25002,N25003,N25004,N25005,N25006,N25007,N25008,
N25009,N25010,N25011,N25012,N25013,N25014,N25015,N25016,N25017,N25018,
N25019,N25020,N25021,N25022,N25023,N25024,N25025,N25026,N25027,N25028,
N25029,N25030,N25031,N25032,N25033,N25034,N25035,N25036,N25037,N25038,
N25039,N25040,N25041,N25042,N25043,N25044,N25045,N25046,N25047,N25048,
N25049,N25050,N25051,N25052,N25053,N25054,N25055,N25056,N25057,N25058,
N25059,N25060,N25061,N25062,N25063,N25064,N25065,N25066,N25067,N25068,
N25069,N25070,N25071,N25072,N25073,N25074,N25075,N25076,N25077,N25078,
N25079,N25080,N25081,N25082,N25083,N25084,N25085,N25086,N25087,N25088,
N25089,N25090,N25091,N25092,N25093,N25094,N25095,N25096,N25097,N25098,
N25099,N25100,N25101,N25102,N25103,N25104,N25105,N25106,N25107,N25108,
N25109,N25110,N25111,N25112,N25113,N25114,N25115,N25116,N25117,N25118,
N25119,N25120,N25121,N25122,N25123,N25124,N25125,N25126,N25127,N25128,
N25129,N25130,N25131,N25132,N25133,N25134,N25135,N25136,N25137,N25138,
N25139,N25140,N25141,N25142,N25143,N25144,N25145,N25146,N25147,N25148,
N25149,N25150,N25151,N25152,N25153,N25154,N25155,N25156,N25157,N25158,
N25159,N25160,N25161,N25162,N25163,N25164,N25165,N25166,N25167,N25168,
N25169,N25170,N25171,N25172,N25173,N25174,N25175,N25176,N25177,N25178,
N25179,N25180,N25181,N25182,N25183,N25184,N25185,N25186,N25187,N25188,
N25189,N25190,N25191,N25192,N25193,N25194,N25195,N25196,N25197,N25198,
N25199,N25200,N25201,N25202,N25203,N25204,N25205,N25206,N25207,N25208,
N25209,N25210,N25211,N25212,N25213,N25214,N25215,N25216,N25217,N25218,
N25219,N25220,N25221,N25222,N25223,N25224,N25225,N25226,N25227,N25228,
N25229,N25230,N25231,N25232,N25233,N25234,N25235,N25236,N25237,N25238,
N25239,N25240,N25241,N25242,N25243,N25244,N25245,N25246,N25247,N25248,
N25249,N25250,N25251,N25252,N25253,N25254,N25255,N25256,N25257,N25258,
N25259,N25260,N25261,N25262,N25263,N25264,N25265,N25266,N25267,N25268,
N25269,N25270,N25271,N25272,N25273,N25274,N25275,N25276,N25277,N25278,
N25279,N25280,N25281,N25282,N25283,N25284,N25285,N25286,N25287,N25288,
N25289,N25290,N25291,N25292,N25293,N25294,N25295,N25296,N25297,N25298,
N25299,N25300,N25301,N25302,N25303,N25304,N25305,N25306,N25307,N25308,
N25309,N25310,N25311,N25312,N25313,N25314,N25315,N25316,N25317,N25318,
N25319,N25320,N25321,N25322,N25323,N25324,N25325,N25326,N25327,N25328,
N25329,N25330,N25331,N25332,N25333,N25334,N25335,N25336,N25337,N25338,
N25339,N25340,N25341,N25342,N25343,N25344,N25345,N25346,N25347,N25348,
N25349,N25350,N25351,N25352,N25353,N25354,N25355,N25356,N25357,N25358,
N25359,N25360,N25361,N25362,N25363,N25364,N25365,N25366,N25367,N25368,
N25369,N25370,N25371,N25372,N25373,N25374,N25375,N25376,N25377,N25378,
N25379,N25380,N25381,N25382,N25383,N25384,N25385,N25386,N25387,N25388,
N25389,N25390,N25391,N25392,N25393,N25394,N25395,N25396,N25397,N25398,
N25399,N25400,N25401,N25402,N25403,N25404,N25405,N25406,N25407,N25408,
N25409,N25410,N25411,N25412,N25413,N25414,N25415,N25416,N25417,N25418,
N25419,N25420,N25421,N25422,N25423,N25424,N25425,N25426,N25427,N25428,
N25429,N25430,N25431,N25432,N25433,N25434,N25435,N25436,N25437,N25438,
N25439,N25440,N25441,N25442,N25443,N25444,N25445,N25446,N25447,N25448,
N25449,N25450,N25451,N25452,N25453,N25454,N25455,N25456,N25457,N25458,
N25459,N25460,N25461,N25462,N25463,N25464,N25465,N25466,N25467,N25468,
N25469,N25470,N25471,N25472,N25473,N25474,N25475,N25476,N25477,N25478,
N25479,N25480,N25481,N25482,N25483,N25484,N25485,N25486,N25487,N25488,
N25489,N25490,N25491,N25492,N25493,N25494,N25495,N25496,N25497,N25498,
N25499,N25500,N25501,N25502,N25503,N25504,N25505,N25506,N25507,N25508,
N25509,N25510,N25511,N25512,N25513,N25514,N25515,N25516,N25517,N25518,
N25519,N25520,N25521,N25522,N25523,N25524,N25525,N25526,N25527,N25528,
N25529,N25530,N25531,N25532,N25533,N25534,N25535,N25536,N25537,N25538,
N25539,N25540,N25541,N25542,N25543,N25544,N25545,N25546,N25547,N25548,
N25549,N25550,N25551,N25552,N25553,N25554,N25555,N25556,N25557,N25558,
N25559,N25560,N25561,N25562,N25563,N25564,N25565,N25566,N25567,N25568,
N25569,N25570,N25571,N25572,N25573,N25574,N25575,N25576,N25577,N25578,
N25579,N25580,N25581,N25582,N25583,N25584,N25585,N25586,N25587,N25588,
N25589,N25590,N25591,N25592,N25593,N25594,N25595,N25596,N25597,N25598,
N25599,N25600,N25601,N25602,N25603,N25604,N25605,N25606,N25607,N25608,
N25609,N25610,N25611,N25612,N25613,N25614,N25615,N25616,N25617,N25618,
N25619,N25620,N25621,N25622,N25623,N25624,N25625,N25626,N25627,N25628,
N25629,N25630,N25631,N25632,N25633,N25634,N25635,N25636,N25637,N25638,
N25639,N25640,N25641,N25642,N25643,N25644,N25645,N25646,N25647,N25648,
N25649,N25650,N25651,N25652,N25653,N25654,N25655,N25656,N25657,N25658,
N25659,N25660,N25661,N25662,N25663,N25664,N25665,N25666,N25667,N25668,
N25669,N25670,N25671,N25672,N25673,N25674,N25675,N25676,N25677,N25678,
N25679,N25680,N25681,N25682,N25683,N25684,N25685,N25686,N25687,N25688,
N25689,N25690,N25691,N25692,N25693,N25694,N25695,N25696,N25697,N25698,
N25699,N25700,N25701,N25702,N25703,N25704,N25705,N25706,N25707,N25708,
N25709,N25710,N25711,N25712,N25713,N25714,N25715,N25716,N25717,N25718,
N25719,N25720,N25721,N25722,N25723,N25724,N25725,N25726,N25727,N25728,
N25729,N25730,N25731,N25732,N25733,N25734,N25735,N25736,N25737,N25738,
N25739,N25740,N25741,N25742,N25743,N25744,N25745,N25746,N25747,N25748,
N25749,N25750,N25751,N25752,N25753,N25754,N25755,N25756,N25757,N25758,
N25759,N25760,N25761,N25762,N25763,N25764,N25765,N25766,N25767,N25768,
N25769,N25770,N25771,N25772,N25773,N25774,N25775,N25776,N25777,N25778,
N25779,N25780,N25781,N25782,N25783,N25784,N25785,N25786,N25787,N25788,
N25789,N25790,N25791,N25792,N25793,N25794,N25795,N25796,N25797,N25798,
N25799,N25800,N25801,N25802,N25803,N25804,N25805,N25806,N25807,N25808,
N25809,N25810,N25811,N25812,N25813,N25814,N25815,N25816,N25817,N25818,
N25819,N25820,N25821,N25822,N25823,N25824,N25825,N25826,N25827,N25828,
N25829,N25830,N25831,N25832,N25833,N25834,N25835,N25836,N25837,N25838,
N25839,N25840,N25841,N25842,N25843,N25844,N25845,N25846,N25847,N25848,
N25849,N25850,N25851,N25852,N25853,N25854,N25855,N25856,N25857,N25858,
N25859,N25860,N25861,N25862,N25863,N25864,N25865,N25866,N25867,N25868,
N25869,N25870,N25871,N25872,N25873,N25874,N25875,N25876,N25877,N25878,
N25879,N25880,N25881,N25882,N25883,N25884,N25885,N25886,N25887,N25888,
N25889,N25890,N25891,N25892,N25893,N25894,N25895,N25896,N25897,N25898,
N25899,N25900,N25901,N25902,N25903,N25904,N25905,N25906,N25907,N25908,
N25909,N25910,N25911,N25912,N25913,N25914,N25915,N25916,N25917,N25918,
N25919,N25920,N25921,N25922,N25923,N25924,N25925,N25926,N25927,N25928,
N25929,N25930,N25931,N25932,N25933,N25934,N25935,N25936,N25937,N25938,
N25939,N25940,N25941,N25942,N25943,N25944,N25945,N25946,N25947,N25948,
N25949,N25950,N25951,N25952,N25953,N25954,N25955,N25956,N25957,N25958,
N25959,N25960,N25961,N25962,N25963,N25964,N25965,N25966,N25967,N25968,
N25969,N25970,N25971,N25972,N25973,N25974,N25975,N25976,N25977,N25978,
N25979,N25980,N25981,N25982,N25983,N25984,N25985,N25986,N25987,N25988,
N25989,N25990,N25991,N25992,N25993,N25994,N25995,N25996,N25997,N25998,
N25999,N26000,N26001,N26002,N26003,N26004,N26005,N26006,N26007,N26008,
N26009,N26010,N26011,N26012,N26013,N26014,N26015,N26016,N26017,N26018,
N26019,N26020,N26021,N26022,N26023,N26024,N26025,N26026,N26027,N26028,
N26029,N26030,N26031,N26032,N26033,N26034,N26035,N26036,N26037,N26038,
N26039,N26040,N26041,N26042,N26043,N26044,N26045,N26046,N26047,N26048,
N26049,N26050,N26051,N26052,N26053,N26054,N26055,N26056,N26057,N26058,
N26059,N26060,N26061,N26062,N26063,N26064,N26065,N26066,N26067,N26068,
N26069,N26070,N26071,N26072,N26073,N26074,N26075,N26076,N26077,N26078,
N26079,N26080,N26081,N26082,N26083,N26084,N26085,N26086,N26087,N26088,
N26089,N26090,N26091,N26092,N26093,N26094,N26095,N26096,N26097,N26098,
N26099,N26100,N26101,N26102,N26103,N26104,N26105,N26106,N26107,N26108,
N26109,N26110,N26111,N26112,N26113,N26114,N26115,N26116,N26117,N26118,
N26119,N26120,N26121,N26122,N26123,N26124,N26125,N26126,N26127,N26128,
N26129,N26130,N26131,N26132,N26133,N26134,N26135,N26136,N26137,N26138,
N26139,N26140,N26141,N26142,N26143,N26144,N26145,N26146,N26147,N26148,
N26149,N26150,N26151,N26152,N26153,N26154,N26155,N26156,N26157,N26158,
N26159,N26160,N26161,N26162,N26163,N26164,N26165,N26166,N26167,N26168,
N26169,N26170,N26171,N26172,N26173,N26174,N26175,N26176,N26177,N26178,
N26179,N26180,N26181,N26182,N26183,N26184,N26185,N26186,N26187,N26188,
N26189,N26190,N26191,N26192,N26193,N26194,N26195,N26196,N26197,N26198,
N26199,N26200,N26201,N26202,N26203,N26204,N26205,N26206,N26207,N26208,
N26209,N26210,N26211,N26212,N26213,N26214,N26215,N26216,N26217,N26218,
N26219,N26220,N26221,N26222,N26223,N26224,N26225,N26226,N26227,N26228,
N26229,N26230,N26231,N26232,N26233,N26234,N26235,N26236,N26237,N26238,
N26239,N26240,N26241,N26242,N26243,N26244,N26245,N26246,N26247,N26248,
N26249,N26250,N26251,N26252,N26253,N26254,N26255,N26256,N26257,N26258,
N26259,N26260,N26261,N26262,N26263,N26264,N26265,N26266,N26267,N26268,
N26269,N26270,N26271,N26272,N26273,N26274,N26275,N26276,N26277,N26278,
N26279,N26280,N26281,N26282,N26283,N26284,N26285,N26286,N26287,N26288,
N26289,N26290,N26291,N26292,N26293,N26294,N26295,N26296,N26297,N26298,
N26299,N26300,N26301,N26302,N26303,N26304,N26305,N26306,N26307,N26308,
N26309,N26310,N26311,N26312,N26313,N26314,N26315,N26316,N26317,N26318,
N26319,N26320,N26321,N26322,N26323,N26324,N26325,N26326,N26327,N26328,
N26329,N26330,N26331,N26332,N26333,N26334,N26335,N26336,N26337,N26338,
N26339,N26340,N26341,N26342,N26343,N26344,N26345,N26346,N26347,N26348,
N26349,N26350,N26351,N26352,N26353,N26354,N26355,N26356,N26357,N26358,
N26359,N26360,N26361,N26362,N26363,N26364,N26365,N26366,N26367,N26368,
N26369,N26370,N26371,N26372,N26373,N26374,N26375,N26376,N26377,N26378,
N26379,N26380,N26381,N26382,N26383,N26384,N26385,N26386,N26387,N26388,
N26389,N26390,N26391,N26392,N26393,N26394,N26395,N26396,N26397,N26398,
N26399,N26400,N26401,N26402,N26403,N26404,N26405,N26406,N26407,N26408,
N26409,N26410,N26411,N26412,N26413,N26414,N26415,N26416,N26417,N26418,
N26419,N26420,N26421,N26422,N26423,N26424,N26425,N26426,N26427,N26428,
N26429,N26430,N26431,N26432,N26433,N26434,N26435,N26436,N26437,N26438,
N26439,N26440,N26441,N26442,N26443,N26444,N26445,N26446,N26447,N26448,
N26449,N26450,N26451,N26452,N26453,N26454,N26455,N26456,N26457,N26458,
N26459,N26460,N26461,N26462,N26463,N26464,N26465,N26466,N26467,N26468,
N26469,N26470,N26471,N26472,N26473,N26474,N26475,N26476,N26477,N26478,
N26479,N26480,N26481,N26482,N26483,N26484,N26485,N26486,N26487,N26488,
N26489,N26490,N26491,N26492,N26493,N26494,N26495,N26496,N26497,N26498,
N26499,N26500,N26501,N26502,N26503,N26504,N26505,N26506,N26507,N26508,
N26509,N26510,N26511,N26512,N26513,N26514,N26515,N26516,N26517,N26518,
N26519,N26520,N26521,N26522,N26523,N26524,N26525,N26526,N26527,N26528,
N26529,N26530,N26531,N26532,N26533,N26534,N26535,N26536,N26537,N26538,
N26539,N26540,N26541,N26542,N26543,N26544,N26545,N26546,N26547,N26548,
N26549,N26550,N26551,N26552,N26553,N26554,N26555,N26556,N26557,N26558,
N26559,N26560,N26561,N26562,N26563,N26564,N26565,N26566,N26567,N26568,
N26569,N26570,N26571,N26572,N26573,N26574,N26575,N26576,N26577,N26578,
N26579,N26580,N26581,N26582,N26583,N26584,N26585,N26586,N26587,N26588,
N26589,N26590,N26591,N26592,N26593,N26594,N26595,N26596,N26597,N26598,
N26599,N26600,N26601,N26602,N26603,N26604,N26605,N26606,N26607,N26608,
N26609,N26610,N26611,N26612,N26613,N26614,N26615,N26616,N26617,N26618,
N26619,N26620,N26621,N26622,N26623,N26624,N26625,N26626,N26627,N26628,
N26629,N26630,N26631,N26632,N26633,N26634,N26635,N26636,N26637,N26638,
N26639,N26640,N26641,N26642,N26643,N26644,N26645,N26646,N26647,N26648,
N26649,N26650,N26651,N26652,N26653,N26654,N26655,N26656,N26657,N26658,
N26659,N26660,N26661,N26662,N26663,N26664,N26665,N26666,N26667,N26668,
N26669,N26670,N26671,N26672,N26673,N26674,N26675,N26676,N26677,N26678,
N26679,N26680,N26681,N26682,N26683,N26684,N26685,N26686,N26687,N26688,
N26689,N26690,N26691,N26692,N26693,N26694,N26695,N26696,N26697,N26698,
N26699,N26700,N26701,N26702,N26703,N26704,N26705,N26706,N26707,N26708,
N26709,N26710,N26711,N26712,N26713,N26714,N26715,N26716,N26717,N26718,
N26719,N26720,N26721,N26722,N26723,N26724,N26725,N26726,N26727,N26728,
N26729,N26730,N26731,N26732,N26733,N26734,N26735,N26736,N26737,N26738,
N26739,N26740,N26741,N26742,N26743,N26744,N26745,N26746,N26747,N26748,
N26749,N26750,N26751,N26752,N26753,N26754,N26755,N26756,N26757,N26758,
N26759,N26760,N26761,N26762,N26763,N26764,N26765,N26766,N26767,N26768,
N26769,N26770,N26771,N26772,N26773,N26774,N26775,N26776,N26777,N26778,
N26779,N26780,N26781,N26782,N26783,N26784,N26785,N26786,N26787,N26788,
N26789,N26790,N26791,N26792,N26793,N26794,N26795,N26796,N26797,N26798,
N26799,N26800,N26801,N26802,N26803,N26804,N26805,N26806,N26807,N26808,
N26809,N26810,N26811,N26812,N26813,N26814,N26815,N26816,N26817,N26818,
N26819,N26820,N26821,N26822,N26823,N26824,N26825,N26826,N26827,N26828,
N26829,N26830,N26831,N26832,N26833,N26834,N26835,N26836,N26837,N26838,
N26839,N26840,N26841,N26842,N26843,N26844,N26845,N26846,N26847,N26848,
N26849,N26850,N26851,N26852,N26853,N26854,N26855,N26856,N26857,N26858,
N26859,N26860,N26861,N26862,N26863,N26864,N26865,N26866,N26867,N26868,
N26869,N26870,N26871,N26872,N26873,N26874,N26875,N26876,N26877,N26878,
N26879,N26880,N26881,N26882,N26883,N26884,N26885,N26886,N26887,N26888,
N26889,N26890,N26891,N26892,N26893,N26894,N26895,N26896,N26897,N26898,
N26899,N26900,N26901,N26902,N26903,N26904,N26905,N26906,N26907,N26908,
N26909,N26910,N26911,N26912,N26913,N26914,N26915,N26916,N26917,N26918,
N26919,N26920,N26921,N26922,N26923,N26924,N26925,N26926,N26927,N26928,
N26929,N26930,N26931,N26932,N26933,N26934,N26935,N26936,N26937,N26938,
N26939,N26940,N26941,N26942,N26943,N26944,N26945,N26946,N26947,N26948,
N26949,N26950,N26951,N26952,N26953,N26954,N26955,N26956,N26957,N26958,
N26959,N26960,N26961,N26962,N26963,N26964,N26965,N26966,N26967,N26968,
N26969,N26970,N26971,N26972,N26973,N26974,N26975,N26976,N26977,N26978,
N26979,N26980,N26981,N26982,N26983,N26984,N26985,N26986,N26987,N26988,
N26989,N26990,N26991,N26992,N26993,N26994,N26995,N26996,N26997,N26998,
N26999,N27000,N27001,N27002,N27003,N27004,N27005,N27006,N27007,N27008,
N27009,N27010,N27011,N27012,N27013,N27014,N27015,N27016,N27017,N27018,
N27019,N27020,N27021,N27022,N27023,N27024,N27025,N27026,N27027,N27028,
N27029,N27030,N27031,N27032,N27033,N27034,N27035,N27036,N27037,N27038,
N27039,N27040,N27041,N27042,N27043,N27044,N27045,N27046,N27047,N27048,
N27049,N27050,N27051,N27052,N27053,N27054,N27055,N27056,N27057,N27058,
N27059,N27060,N27061,N27062,N27063,N27064,N27065,N27066,N27067,N27068,
N27069,N27070,N27071,N27072,N27073,N27074,N27075,N27076,N27077,N27078,
N27079,N27080,N27081,N27082,N27083,N27084,N27085,N27086,N27087,N27088,
N27089,N27090,N27091,N27092,N27093,N27094,N27095,N27096,N27097,N27098,
N27099,N27100,N27101,N27102,N27103,N27104,N27105,N27106,N27107,N27108,
N27109,N27110,N27111,N27112,N27113,N27114,N27115,N27116,N27117,N27118,
N27119,N27120,N27121,N27122,N27123,N27124,N27125,N27126,N27127,N27128,
N27129,N27130,N27131,N27132,N27133,N27134,N27135,N27136,N27137,N27138,
N27139,N27140,N27141,N27142,N27143,N27144,N27145,N27146,N27147,N27148,
N27149,N27150,N27151,N27152,N27153,N27154,N27155,N27156,N27157,N27158,
N27159,N27160,N27161,N27162,N27163,N27164,N27165,N27166,N27167,N27168,
N27169,N27170,N27171,N27172,N27173,N27174,N27175,N27176,N27177,N27178,
N27179,N27180,N27181,N27182,N27183,N27184,N27185,N27186,N27187,N27188,
N27189,N27190,N27191,N27192,N27193,N27194,N27195,N27196,N27197,N27198,
N27199,N27200,N27201,N27202,N27203,N27204,N27205,N27206,N27207,N27208,
N27209,N27210,N27211,N27212,N27213,N27214,N27215,N27216,N27217,N27218,
N27219,N27220,N27221,N27222,N27223,N27224,N27225,N27226,N27227,N27228,
N27229,N27230,N27231,N27232,N27233,N27234,N27235,N27236,N27237,N27238,
N27239,N27240,N27241,N27242,N27243,N27244,N27245,N27246,N27247,N27248,
N27249,N27250,N27251,N27252,N27253,N27254,N27255,N27256,N27257,N27258,
N27259,N27260,N27261,N27262,N27263,N27264,N27265,N27266,N27267,N27268,
N27269,N27270,N27271,N27272,N27273,N27274,N27275,N27276,N27277,N27278,
N27279,N27280,N27281,N27282,N27283,N27284,N27285,N27286,N27287,N27288,
N27289,N27290,N27291,N27292,N27293,N27294,N27295,N27296,N27297,N27298,
N27299,N27300,N27301,N27302,N27303,N27304,N27305,N27306,N27307,N27308,
N27309,N27310,N27311,N27312,N27313,N27314,N27315,N27316,N27317,N27318,
N27319,N27320,N27321,N27322,N27323,N27324,N27325,N27326,N27327,N27328,
N27329,N27330,N27331,N27332,N27333,N27334,N27335,N27336,N27337,N27338,
N27339,N27340,N27341,N27342,N27343,N27344,N27345,N27346,N27347,N27348,
N27349,N27350,N27351,N27352,N27353,N27354,N27355,N27356,N27357,N27358,
N27359,N27360,N27361,N27362,N27363,N27364,N27365,N27366,N27367,N27368,
N27369,N27370,N27371,N27372,N27373,N27374,N27375,N27376,N27377,N27378,
N27379,N27380,N27381,N27382,N27383,N27384,N27385,N27386,N27387,N27388,
N27389,N27390,N27391,N27392,N27393,N27394,N27395,N27396,N27397,N27398,
N27399,N27400,N27401,N27402,N27403,N27404,N27405,N27406,N27407,N27408,
N27409,N27410,N27411,N27412,N27413,N27414,N27415,N27416,N27417,N27418,
N27419,N27420,N27421,N27422,N27423,N27424,N27425,N27426,N27427,N27428,
N27429,N27430,N27431,N27432,N27433,N27434,N27435,N27436,N27437,N27438,
N27439,N27440,N27441,N27442,N27443,N27444,N27445,N27446,N27447,N27448,
N27449,N27450,N27451,N27452,N27453,N27454,N27455,N27456,N27457,N27458,
N27459,N27460,N27461,N27462,N27463,N27464,N27465,N27466,N27467,N27468,
N27469,N27470,N27471,N27472,N27473,N27474,N27475,N27476,N27477,N27478,
N27479,N27480,N27481,N27482,N27483,N27484,N27485,N27486,N27487,N27488,
N27489,N27490,N27491,N27492,N27493,N27494,N27495,N27496,N27497,N27498,
N27499,N27500,N27501,N27502,N27503,N27504,N27505,N27506,N27507,N27508,
N27509,N27510,N27511,N27512,N27513,N27514,N27515,N27516,N27517,N27518,
N27519,N27520,N27521,N27522,N27523,N27524,N27525,N27526,N27527,N27528,
N27529,N27530,N27531,N27532,N27533,N27534,N27535,N27536,N27537,N27538,
N27539,N27540,N27541,N27542,N27543,N27544,N27545,N27546,N27547,N27548,
N27549,N27550,N27551,N27552,N27553,N27554,N27555,N27556,N27557,N27558,
N27559,N27560,N27561,N27562,N27563,N27564,N27565,N27566,N27567,N27568,
N27569,N27570,N27571,N27572,N27573,N27574,N27575,N27576,N27577,N27578,
N27579,N27580,N27581,N27582,N27583,N27584,N27585,N27586,N27587,N27588,
N27589,N27590,N27591,N27592,N27593,N27594,N27595,N27596,N27597,N27598,
N27599,N27600,N27601,N27602,N27603,N27604,N27605,N27606,N27607,N27608,
N27609,N27610,N27611,N27612,N27613,N27614,N27615,N27616,N27617,N27618,
N27619,N27620,N27621,N27622,N27623,N27624,N27625,N27626,N27627,N27628,
N27629,N27630,N27631,N27632,N27633,N27634,N27635,N27636,N27637,N27638,
N27639,N27640,N27641,N27642,N27643,N27644,N27645,N27646,N27647,N27648,
N27649,N27650,N27651,N27652,N27653,N27654,N27655,N27656,N27657,N27658,
N27659,N27660,N27661,N27662,N27663,N27664,N27665,N27666,N27667,N27668,
N27669,N27670,N27671,N27672,N27673,N27674,N27675,N27676,N27677,N27678,
N27679,N27680,N27681,N27682,N27683,N27684,N27685,N27686,N27687,N27688,
N27689,N27690,N27691,N27692,N27693,N27694,N27695,N27696,N27697,N27698,
N27699,N27700,N27701,N27702,N27703,N27704,N27705,N27706,N27707,N27708,
N27709,N27710,N27711,N27712,N27713,N27714,N27715,N27716,N27717,N27718,
N27719,N27720,N27721,N27722,N27723,N27724,N27725,N27726,N27727,N27728,
N27729,N27730,N27731,N27732,N27733,N27734,N27735,N27736,N27737,N27738,
N27739,N27740,N27741,N27742,N27743,N27744,N27745,N27746,N27747,N27748,
N27749,N27750,N27751,N27752,N27753,N27754,N27755,N27756,N27757,N27758,
N27759,N27760,N27761,N27762,N27763,N27764,N27765,N27766,N27767,N27768,
N27769,N27770,N27771,N27772,N27773,N27774,N27775,N27776,N27777,N27778,
N27779,N27780,N27781,N27782,N27783,N27784,N27785,N27786,N27787,N27788,
N27789,N27790,N27791,N27792,N27793,N27794,N27795,N27796,N27797,N27798,
N27799,N27800,N27801,N27802,N27803,N27804,N27805,N27806,N27807,N27808,
N27809,N27810,N27811,N27812,N27813,N27814,N27815,N27816,N27817,N27818,
N27819,N27820,N27821,N27822,N27823,N27824,N27825,N27826,N27827,N27828,
N27829,N27830,N27831,N27832,N27833,N27834,N27835,N27836,N27837,N27838,
N27839,N27840,N27841,N27842,N27843,N27844,N27845,N27846,N27847,N27848,
N27849,N27850,N27851,N27852,N27853,N27854,N27855,N27856,N27857,N27858,
N27859,N27860,N27861,N27862,N27863,N27864,N27865,N27866,N27867,N27868,
N27869,N27870,N27871,N27872,N27873,N27874,N27875,N27876,N27877,N27878,
N27879,N27880,N27881,N27882,N27883,N27884,N27885,N27886,N27887,N27888,
N27889,N27890,N27891,N27892,N27893,N27894,N27895,N27896,N27897,N27898,
N27899,N27900,N27901,N27902,N27903,N27904,N27905,N27906,N27907,N27908,
N27909,N27910,N27911,N27912,N27913,N27914,N27915,N27916,N27917,N27918,
N27919,N27920,N27921,N27922,N27923,N27924,N27925,N27926,N27927,N27928,
N27929,N27930,N27931,N27932,N27933,N27934,N27935,N27936,N27937,N27938,
N27939,N27940,N27941,N27942,N27943,N27944,N27945,N27946,N27947,N27948,
N27949,N27950,N27951,N27952,N27953,N27954,N27955,N27956,N27957,N27958,
N27959,N27960,N27961,N27962,N27963,N27964,N27965,N27966,N27967,N27968,
N27969,N27970,N27971,N27972,N27973,N27974,N27975,N27976,N27977,N27978,
N27979,N27980,N27981,N27982,N27983,N27984,N27985,N27986,N27987,N27988,
N27989,N27990,N27991,N27992,N27993,N27994,N27995,N27996,N27997,N27998,
N27999,N28000,N28001,N28002,N28003,N28004,N28005,N28006,N28007,N28008,
N28009,N28010,N28011,N28012,N28013,N28014,N28015,N28016,N28017,N28018,
N28019,N28020,N28021,N28022,N28023,N28024,N28025,N28026,N28027,N28028,
N28029,N28030,N28031,N28032,N28033,N28034,N28035,N28036,N28037,N28038,
N28039,N28040,N28041,N28042,N28043,N28044,N28045,N28046,N28047,N28048,
N28049,N28050,N28051,N28052,N28053,N28054,N28055,N28056,N28057,N28058,
N28059,N28060,N28061,N28062,N28063,N28064,N28065,N28066,N28067,N28068,
N28069,N28070,N28071,N28072,N28073,N28074,N28075,N28076,N28077,N28078,
N28079,N28080,N28081,N28082,N28083,N28084,N28085,N28086,N28087,N28088,
N28089,N28090,N28091,N28092,N28093,N28094,N28095,N28096,N28097,N28098,
N28099,N28100,N28101,N28102,N28103,N28104,N28105,N28106,N28107,N28108,
N28109,N28110,N28111,N28112,N28113,N28114,N28115,N28116,N28117,N28118,
N28119,N28120,N28121,N28122,N28123,N28124,N28125,N28126,N28127,N28128,
N28129,N28130,N28131,N28132,N28133,N28134,N28135,N28136,N28137,N28138,
N28139,N28140,N28141,N28142,N28143,N28144,N28145,N28146,N28147,N28148,
N28149,N28150,N28151,N28152,N28153,N28154,N28155,N28156,N28157,N28158,
N28159,N28160,N28161,N28162,N28163,N28164,N28165,N28166,N28167,N28168,
N28169,N28170,N28171,N28172,N28173,N28174,N28175,N28176,N28177,N28178,
N28179,N28180,N28181,N28182,N28183,N28184,N28185,N28186,N28187,N28188,
N28189,N28190,N28191,N28192,N28193,N28194,N28195,N28196,N28197,N28198,
N28199,N28200,N28201,N28202,N28203,N28204,N28205,N28206,N28207,N28208,
N28209,N28210,N28211,N28212,N28213,N28214,N28215,N28216,N28217,N28218,
N28219,N28220,N28221,N28222,N28223,N28224,N28225,N28226,N28227,N28228,
N28229,N28230,N28231,N28232,N28233,N28234,N28235,N28236,N28237,N28238,
N28239,N28240,N28241,N28242,N28243,N28244,N28245,N28246,N28247,N28248,
N28249,N28250,N28251,N28252,N28253,N28254,N28255,N28256,N28257,N28258,
N28259,N28260,N28261,N28262,N28263,N28264,N28265,N28266,N28267,N28268,
N28269,N28270,N28271,N28272,N28273,N28274,N28275,N28276,N28277,N28278,
N28279,N28280,N28281,N28282,N28283,N28284,N28285,N28286,N28287,N28288,
N28289,N28290,N28291,N28292,N28293,N28294,N28295,N28296,N28297,N28298,
N28299,N28300,N28301,N28302,N28303,N28304,N28305,N28306,N28307,N28308,
N28309,N28310,N28311,N28312,N28313,N28314,N28315,N28316,N28317,N28318,
N28319,N28320,N28321,N28322,N28323,N28324,N28325,N28326,N28327,N28328,
N28329,N28330,N28331,N28332,N28333,N28334,N28335,N28336,N28337,N28338,
N28339,N28340,N28341,N28342,N28343,N28344,N28345,N28346,N28347,N28348,
N28349,N28350,N28351,N28352,N28353,N28354,N28355,N28356,N28357,N28358,
N28359,N28360,N28361,N28362,N28363,N28364,N28365,N28366,N28367,N28368,
N28369,N28370,N28371,N28372,N28373,N28374,N28375,N28376,N28377,N28378,
N28379,N28380,N28381,N28382,N28383,N28384,N28385,N28386,N28387,N28388,
N28389,N28390,N28391,N28392,N28393,N28394,N28395,N28396,N28397,N28398,
N28399,N28400,N28401,N28402,N28403,N28404,N28405,N28406,N28407,N28408,
N28409,N28410,N28411,N28412,N28413,N28414,N28415,N28416,N28417,N28418,
N28419,N28420,N28421,N28422,N28423,N28424,N28425,N28426,N28427,N28428,
N28429,N28430,N28431,N28432,N28433,N28434,N28435,N28436,N28437,N28438,
N28439,N28440,N28441,N28442,N28443,N28444,N28445,N28446,N28447,N28448,
N28449,N28450,N28451,N28452,N28453,N28454,N28455,N28456,N28457,N28458,
N28459,N28460,N28461,N28462,N28463,N28464,N28465,N28466,N28467,N28468,
N28469,N28470,N28471,N28472,N28473,N28474,N28475,N28476,N28477,N28478,
N28479,N28480,N28481,N28482,N28483,N28484,N28485,N28486,N28487,N28488,
N28489,N28490,N28491,N28492,N28493,N28494,N28495,N28496,N28497,N28498,
N28499,N28500,N28501,N28502,N28503,N28504,N28505,N28506,N28507,N28508,
N28509,N28510,N28511,N28512,N28513,N28514,N28515,N28516,N28517,N28518,
N28519,N28520,N28521,N28522,N28523,N28524,N28525,N28526,N28527,N28528,
N28529,N28530,N28531,N28532,N28533,N28534,N28535,N28536,N28537,N28538,
N28539,N28540,N28541,N28542,N28543,N28544,N28545,N28546,N28547,N28548,
N28549,N28550,N28551,N28552,N28553,N28554,N28555,N28556,N28557,N28558,
N28559,N28560,N28561,N28562,N28563,N28564,N28565,N28566,N28567,N28568,
N28569,N28570,N28571,N28572,N28573,N28574,N28575,N28576,N28577,N28578,
N28579,N28580,N28581,N28582,N28583,N28584,N28585,N28586,N28587,N28588,
N28589,N28590,N28591,N28592,N28593,N28594,N28595,N28596,N28597,N28598,
N28599,N28600,N28601,N28602,N28603,N28604,N28605,N28606,N28607,N28608,
N28609,N28610,N28611,N28612,N28613,N28614,N28615,N28616,N28617,N28618,
N28619,N28620,N28621,N28622,N28623,N28624,N28625,N28626,N28627,N28628,
N28629,N28630,N28631,N28632,N28633,N28634,N28635,N28636,N28637,N28638,
N28639,N28640,N28641,N28642,N28643,N28644,N28645,N28646,N28647,N28648,
N28649,N28650,N28651,N28652,N28653,N28654,N28655,N28656,N28657,N28658,
N28659,N28660,N28661,N28662,N28663,N28664,N28665,N28666,N28667,N28668,
N28669,N28670,N28671,N28672,N28673,N28674,N28675,N28676,N28677,N28678,
N28679,N28680,N28681,N28682,N28683,N28684,N28685,N28686,N28687,N28688,
N28689,N28690,N28691,N28692,N28693,N28694,N28695,N28696,N28697,N28698,
N28699,N28700,N28701,N28702,N28703,N28704,N28705,N28706,N28707,N28708,
N28709,N28710,N28711,N28712,N28713,N28714,N28715,N28716,N28717,N28718,
N28719,N28720,N28721,N28722,N28723,N28724,N28725,N28726,N28727,N28728,
N28729,N28730,N28731,N28732,N28733,N28734,N28735,N28736,N28737,N28738,
N28739,N28740,N28741,N28742,N28743,N28744,N28745,N28746,N28747,N28748,
N28749,N28750,N28751,N28752,N28753,N28754,N28755,N28756,N28757,N28758,
N28759,N28760,N28761,N28762,N28763,N28764,N28765,N28766,N28767,N28768,
N28769,N28770,N28771,N28772,N28773,N28774,N28775,N28776,N28777,N28778,
N28779,N28780,N28781,N28782,N28783,N28784,N28785,N28786,N28787,N28788,
N28789,N28790,N28791,N28792,N28793,N28794,N28795,N28796,N28797,N28798,
N28799,N28800,N28801,N28802,N28803,N28804,N28805,N28806,N28807,N28808,
N28809,N28810,N28811,N28812,N28813,N28814,N28815,N28816,N28817,N28818,
N28819,N28820,N28821,N28822,N28823,N28824,N28825,N28826,N28827,N28828,
N28829,N28830,N28831,N28832,N28833,N28834,N28835,N28836,N28837,N28838,
N28839,N28840,N28841,N28842,N28843,N28844,N28845,N28846,N28847,N28848,
N28849,N28850,N28851,N28852,N28853,N28854,N28855,N28856,N28857,N28858,
N28859,N28860,N28861,N28862,N28863,N28864,N28865,N28866,N28867,N28868,
N28869,N28870,N28871,N28872,N28873,N28874,N28875,N28876,N28877,N28878,
N28879,N28880,N28881,N28882,N28883,N28884,N28885,N28886,N28887,N28888,
N28889,N28890,N28891,N28892,N28893,N28894,N28895,N28896,N28897,N28898,
N28899,N28900,N28901,N28902,N28903,N28904,N28905,N28906,N28907,N28908,
N28909,N28910,N28911,N28912,N28913,N28914,N28915,N28916,N28917,N28918,
N28919,N28920,N28921,N28922,N28923,N28924,N28925,N28926,N28927,N28928,
N28929,N28930,N28931,N28932,N28933,N28934,N28935,N28936,N28937,N28938,
N28939,N28940,N28941,N28942,N28943,N28944,N28945,N28946,N28947,N28948,
N28949,N28950,N28951,N28952,N28953,N28954,N28955,N28956,N28957,N28958,
N28959,N28960,N28961,N28962,N28963,N28964,N28965,N28966,N28967,N28968,
N28969,N28970,N28971,N28972,N28973,N28974,N28975,N28976,N28977,N28978,
N28979,N28980,N28981,N28982,N28983,N28984,N28985,N28986,N28987,N28988,
N28989,N28990,N28991,N28992,N28993,N28994,N28995,N28996,N28997,N28998,
N28999,N29000,N29001,N29002,N29003,N29004,N29005,N29006,N29007,N29008,
N29009,N29010,N29011,N29012,N29013,N29014,N29015,N29016,N29017,N29018,
N29019,N29020,N29021,N29022,N29023,N29024,N29025,N29026,N29027,N29028,
N29029,N29030,N29031,N29032,N29033,N29034,N29035,N29036,N29037,N29038,
N29039,N29040,N29041,N29042,N29043,N29044,N29045,N29046,N29047,N29048,
N29049,N29050,N29051,N29052,N29053,N29054,N29055,N29056,N29057,N29058,
N29059,N29060,N29061,N29062,N29063,N29064,N29065,N29066,N29067,N29068,
N29069,N29070,N29071,N29072,N29073,N29074,N29075,N29076,N29077,N29078,
N29079,N29080,N29081,N29082,N29083,N29084,N29085,N29086,N29087,N29088,
N29089,N29090,N29091,N29092,N29093,N29094,N29095,N29096,N29097,N29098,
N29099,N29100,N29101,N29102,N29103,N29104,N29105,N29106,N29107,N29108,
N29109,N29110,N29111,N29112,N29113,N29114,N29115,N29116,N29117,N29118,
N29119,N29120,N29121,N29122,N29123,N29124,N29125,N29126,N29127,N29128,
N29129,N29130,N29131,N29132,N29133,N29134,N29135,N29136,N29137,N29138,
N29139,N29140,N29141,N29142,N29143,N29144,N29145,N29146,N29147,N29148,
N29149,N29150,N29151,N29152,N29153,N29154,N29155,N29156,N29157,N29158,
N29159,N29160,N29161,N29162,N29163,N29164,N29165,N29166,N29167,N29168,
N29169,N29170,N29171,N29172,N29173,N29174,N29175,N29176,N29177,N29178,
N29179,N29180,N29181,N29182,N29183,N29184,N29185,N29186,N29187,N29188,
N29189,N29190,N29191,N29192,N29193,N29194,N29195,N29196,N29197,N29198,
N29199,N29200,N29201,N29202,N29203,N29204,N29205,N29206,N29207,N29208,
N29209,N29210,N29211,N29212,N29213,N29214,N29215,N29216,N29217,N29218,
N29219,N29220,N29221,N29222,N29223,N29224,N29225,N29226,N29227,N29228,
N29229,N29230,N29231,N29232,N29233,N29234,N29235,N29236,N29237,N29238,
N29239,N29240,N29241,N29242,N29243,N29244,N29245,N29246,N29247,N29248,
N29249,N29250,N29251,N29252,N29253,N29254,N29255,N29256,N29257,N29258,
N29259,N29260,N29261,N29262,N29263,N29264,N29265,N29266,N29267,N29268,
N29269,N29270,N29271,N29272,N29273,N29274,N29275,N29276,N29277,N29278,
N29279,N29280,N29281,N29282,N29283,N29284,N29285,N29286,N29287,N29288,
N29289,N29290,N29291,N29292,N29293,N29294,N29295,N29296,N29297,N29298,
N29299,N29300,N29301,N29302,N29303,N29304,N29305,N29306,N29307,N29308,
N29309,N29310,N29311,N29312,N29313,N29314,N29315,N29316,N29317,N29318,
N29319,N29320,N29321,N29322,N29323,N29324,N29325,N29326,N29327,N29328,
N29329,N29330,N29331,N29332,N29333,N29334,N29335,N29336,N29337,N29338,
N29339,N29340,N29341,N29342,N29343,N29344,N29345,N29346,N29347,N29348,
N29349,N29350,N29351,N29352,N29353,N29354,N29355,N29356,N29357,N29358,
N29359,N29360,N29361,N29362,N29363,N29364,N29365,N29366,N29367,N29368,
N29369,N29370,N29371,N29372,N29373,N29374,N29375,N29376,N29377,N29378,
N29379,N29380,N29381,N29382,N29383,N29384,N29385,N29386,N29387,N29388,
N29389,N29390,N29391,N29392,N29393,N29394,N29395,N29396,N29397,N29398,
N29399,N29400,N29401,N29402,N29403,N29404,N29405,N29406,N29407,N29408,
N29409,N29410,N29411,N29412,N29413,N29414,N29415,N29416,N29417,N29418,
N29419,N29420,N29421,N29422,N29423,N29424,N29425,N29426,N29427,N29428,
N29429,N29430,N29431,N29432,N29433,N29434,N29435,N29436,N29437,N29438,
N29439,N29440,N29441,N29442,N29443,N29444,N29445,N29446,N29447,N29448,
N29449,N29450,N29451,N29452,N29453,N29454,N29455,N29456,N29457,N29458,
N29459,N29460,N29461,N29462,N29463,N29464,N29465,N29466,N29467,N29468,
N29469,N29470,N29471,N29472,N29473,N29474,N29475,N29476,N29477,N29478,
N29479,N29480,N29481,N29482,N29483,N29484,N29485,N29486,N29487,N29488,
N29489,N29490,N29491,N29492,N29493,N29494,N29495,N29496,N29497,N29498,
N29499,N29500,N29501,N29502,N29503,N29504,N29505,N29506,N29507,N29508,
N29509,N29510,N29511,N29512,N29513,N29514,N29515,N29516,N29517,N29518,
N29519,N29520,N29521,N29522,N29523,N29524,N29525,N29526,N29527,N29528,
N29529,N29530,N29531,N29532,N29533,N29534,N29535,N29536,N29537,N29538,
N29539,N29540,N29541,N29542,N29543,N29544,N29545,N29546,N29547,N29548,
N29549,N29550,N29551,N29552,N29553,N29554,N29555,N29556,N29557,N29558,
N29559,N29560,N29561,N29562,N29563,N29564,N29565,N29566,N29567,N29568,
N29569,N29570,N29571,N29572,N29573,N29574,N29575,N29576,N29577,N29578,
N29579,N29580,N29581,N29582,N29583,N29584,N29585,N29586,N29587,N29588,
N29589,N29590,N29591,N29592,N29593,N29594,N29595,N29596,N29597,N29598,
N29599,N29600,N29601,N29602,N29603,N29604,N29605,N29606,N29607,N29608,
N29609,N29610,N29611,N29612,N29613,N29614,N29615,N29616,N29617,N29618,
N29619,N29620,N29621,N29622,N29623,N29624,N29625,N29626,N29627,N29628,
N29629,N29630,N29631,N29632,N29633,N29634,N29635,N29636,N29637,N29638,
N29639,N29640,N29641,N29642,N29643,N29644,N29645,N29646,N29647,N29648,
N29649,N29650,N29651,N29652,N29653,N29654,N29655,N29656,N29657,N29658,
N29659,N29660,N29661,N29662,N29663,N29664,N29665,N29666,N29667,N29668,
N29669,N29670,N29671,N29672,N29673,N29674,N29675,N29676,N29677,N29678,
N29679,N29680,N29681,N29682,N29683,N29684,N29685,N29686,N29687,N29688,
N29689,N29690,N29691,N29692,N29693,N29694,N29695,N29696,N29697,N29698,
N29699,N29700,N29701,N29702,N29703,N29704,N29705,N29706,N29707,N29708,
N29709,N29710,N29711,N29712,N29713,N29714,N29715,N29716,N29717,N29718,
N29719,N29720,N29721,N29722,N29723,N29724,N29725,N29726,N29727,N29728,
N29729,N29730,N29731,N29732,N29733,N29734,N29735,N29736,N29737,N29738,
N29739,N29740,N29741,N29742,N29743,N29744,N29745,N29746,N29747,N29748,
N29749,N29750,N29751,N29752,N29753,N29754,N29755,N29756,N29757,N29758,
N29759,N29760,N29761,N29762,N29763,N29764,N29765,N29766,N29767,N29768,
N29769,N29770,N29771,N29772,N29773,N29774,N29775,N29776,N29777,N29778,
N29779,N29780,N29781,N29782,N29783,N29784,N29785,N29786,N29787,N29788,
N29789,N29790,N29791,N29792,N29793,N29794,N29795,N29796,N29797,N29798,
N29799,N29800,N29801,N29802,N29803,N29804,N29805,N29806,N29807,N29808,
N29809,N29810,N29811,N29812,N29813,N29814,N29815,N29816,N29817,N29818,
N29819,N29820,N29821,N29822,N29823,N29824,N29825,N29826,N29827,N29828,
N29829,N29830,N29831,N29832,N29833,N29834,N29835,N29836,N29837,N29838,
N29839,N29840,N29841,N29842,N29843,N29844,N29845,N29846,N29847,N29848,
N29849,N29850,N29851,N29852,N29853,N29854,N29855,N29856,N29857,N29858,
N29859,N29860,N29861,N29862,N29863,N29864,N29865,N29866,N29867,N29868,
N29869,N29870,N29871,N29872,N29873,N29874,N29875,N29876,N29877,N29878,
N29879,N29880,N29881,N29882,N29883,N29884,N29885,N29886,N29887,N29888,
N29889,N29890,N29891,N29892,N29893,N29894,N29895,N29896,N29897,N29898,
N29899,N29900,N29901,N29902,N29903,N29904,N29905,N29906,N29907,N29908,
N29909,N29910,N29911,N29912,N29913,N29914,N29915,N29916,N29917,N29918,
N29919,N29920,N29921,N29922,N29923,N29924,N29925,N29926,N29927,N29928,
N29929,N29930,N29931,N29932,N29933,N29934,N29935,N29936,N29937,N29938,
N29939,N29940,N29941,N29942,N29943,N29944,N29945,N29946,N29947,N29948,
N29949,N29950,N29951,N29952,N29953,N29954,N29955,N29956,N29957,N29958,
N29959,N29960,N29961,N29962,N29963,N29964,N29965,N29966,N29967,N29968,
N29969,N29970,N29971,N29972,N29973,N29974,N29975,N29976,N29977,N29978,
N29979,N29980,N29981,N29982,N29983,N29984,N29985,N29986,N29987,N29988,
N29989,N29990,N29991,N29992,N29993,N29994,N29995,N29996,N29997,N29998,
N29999,N30000,N30001,N30002,N30003,N30004,N30005,N30006,N30007,N30008,
N30009,N30010,N30011,N30012,N30013,N30014,N30015,N30016,N30017,N30018,
N30019,N30020,N30021,N30022,N30023,N30024,N30025,N30026,N30027,N30028,
N30029,N30030,N30031,N30032,N30033,N30034,N30035,N30036,N30037,N30038,
N30039,N30040,N30041,N30042,N30043,N30044,N30045,N30046,N30047,N30048,
N30049,N30050,N30051,N30052,N30053,N30054,N30055,N30056,N30057,N30058,
N30059,N30060,N30061,N30062,N30063,N30064,N30065,N30066,N30067,N30068,
N30069,N30070,N30071,N30072,N30073,N30074,N30075,N30076,N30077,N30078,
N30079,N30080,N30081,N30082,N30083,N30084,N30085,N30086,N30087,N30088,
N30089,N30090,N30091,N30092,N30093,N30094,N30095,N30096,N30097,N30098,
N30099,N30100,N30101,N30102,N30103,N30104,N30105,N30106,N30107,N30108,
N30109,N30110,N30111,N30112,N30113,N30114,N30115,N30116,N30117,N30118,
N30119,N30120,N30121,N30122,N30123,N30124,N30125,N30126,N30127,N30128,
N30129,N30130,N30131,N30132,N30133,N30134,N30135,N30136,N30137,N30138,
N30139,N30140,N30141,N30142,N30143,N30144,N30145,N30146,N30147,N30148,
N30149,N30150,N30151,N30152,N30153,N30154,N30155,N30156,N30157,N30158,
N30159,N30160,N30161,N30162,N30163,N30164,N30165,N30166,N30167,N30168,
N30169,N30170,N30171,N30172,N30173,N30174,N30175,N30176,N30177,N30178,
N30179,N30180,N30181,N30182,N30183,N30184,N30185,N30186,N30187,N30188,
N30189,N30190,N30191,N30192,N30193,N30194,N30195,N30196,N30197,N30198,
N30199,N30200,N30201,N30202,N30203,N30204,N30205,N30206,N30207,N30208,
N30209,N30210,N30211,N30212,N30213,N30214,N30215,N30216,N30217,N30218,
N30219,N30220,N30221,N30222,N30223,N30224,N30225,N30226,N30227,N30228,
N30229,N30230,N30231,N30232,N30233,N30234,N30235,N30236,N30237,N30238,
N30239,N30240,N30241,N30242,N30243,N30244,N30245,N30246,N30247,N30248,
N30249,N30250,N30251,N30252,N30253,N30254,N30255,N30256,N30257,N30258,
N30259,N30260,N30261,N30262,N30263,N30264,N30265,N30266,N30267,N30268,
N30269,N30270,N30271,N30272,N30273,N30274,N30275,N30276,N30277,N30278,
N30279,N30280,N30281,N30282,N30283,N30284,N30285,N30286,N30287,N30288,
N30289,N30290,N30291,N30292,N30293,N30294,N30295,N30296,N30297,N30298,
N30299,N30300,N30301,N30302,N30303,N30304,N30305,N30306,N30307,N30308,
N30309,N30310,N30311,N30312,N30313,N30314,N30315,N30316,N30317,N30318,
N30319,N30320,N30321,N30322,N30323,N30324,N30325,N30326,N30327,N30328,
N30329,N30330,N30331,N30332,N30333,N30334,N30335,N30336,N30337,N30338,
N30339,N30340,N30341,N30342,N30343,N30344,N30345,N30346,N30347,N30348,
N30349,N30350,N30351,N30352,N30353,N30354,N30355,N30356,N30357,N30358,
N30359,N30360,N30361,N30362,N30363,N30364,N30365,N30366,N30367,N30368,
N30369,N30370,N30371,N30372,N30373,N30374,N30375,N30376,N30377,N30378,
N30379,N30380,N30381,N30382,N30383,N30384,N30385,N30386,N30387,N30388,
N30389,N30390,N30391,N30392,N30393,N30394,N30395,N30396,N30397,N30398,
N30399,N30400,N30401,N30402,N30403,N30404,N30405,N30406,N30407,N30408,
N30409,N30410,N30411,N30412,N30413,N30414,N30415,N30416,N30417,N30418,
N30419,N30420,N30421,N30422,N30423,N30424,N30425,N30426,N30427,N30428,
N30429,N30430,N30431,N30432,N30433,N30434,N30435,N30436,N30437,N30438,
N30439,N30440,N30441,N30442,N30443,N30444,N30445,N30446,N30447,N30448,
N30449,N30450,N30451,N30452,N30453,N30454,N30455,N30456,N30457,N30458,
N30459,N30460,N30461,N30462,N30463,N30464,N30465,N30466,N30467,N30468,
N30469,N30470,N30471,N30472,N30473,N30474,N30475,N30476,N30477,N30478,
N30479,N30480,N30481,N30482,N30483,N30484,N30485,N30486,N30487,N30488,
N30489,N30490,N30491,N30492,N30493,N30494,N30495,N30496,N30497,N30498,
N30499,N30500,N30501,N30502,N30503,N30504,N30505,N30506,N30507,N30508,
N30509,N30510,N30511,N30512,N30513,N30514,N30515,N30516,N30517,N30518,
N30519,N30520,N30521,N30522,N30523,N30524,N30525,N30526,N30527,N30528,
N30529,N30530,N30531,N30532,N30533,N30534,N30535,N30536,N30537,N30538,
N30539,N30540,N30541,N30542,N30543,N30544,N30545,N30546,N30547,N30548,
N30549,N30550,N30551,N30552,N30553,N30554,N30555,N30556,N30557,N30558,
N30559,N30560,N30561,N30562,N30563,N30564,N30565,N30566,N30567,N30568,
N30569,N30570,N30571,N30572,N30573,N30574,N30575,N30576,N30577,N30578,
N30579,N30580,N30581,N30582,N30583,N30584,N30585,N30586,N30587,N30588,
N30589,N30590,N30591,N30592,N30593,N30594,N30595,N30596,N30597,N30598,
N30599,N30600,N30601,N30602,N30603,N30604,N30605,N30606,N30607,N30608,
N30609,N30610,N30611,N30612,N30613,N30614,N30615,N30616,N30617,N30618,
N30619,N30620,N30621,N30622,N30623,N30624,N30625,N30626,N30627,N30628,
N30629,N30630,N30631,N30632,N30633,N30634,N30635,N30636,N30637,N30638,
N30639,N30640,N30641,N30642,N30643,N30644,N30645,N30646,N30647,N30648,
N30649,N30650,N30651,N30652,N30653,N30654,N30655,N30656,N30657,N30658,
N30659,N30660,N30661,N30662,N30663,N30664,N30665,N30666,N30667,N30668,
N30669,N30670,N30671,N30672,N30673,N30674,N30675,N30676,N30677,N30678,
N30679,N30680,N30681,N30682,N30683,N30684,N30685,N30686,N30687,N30688,
N30689,N30690,N30691,N30692,N30693,N30694,N30695,N30696,N30697,N30698,
N30699,N30700,N30701,N30702,N30703,N30704,N30705,N30706,N30707,N30708,
N30709,N30710,N30711,N30712,N30713,N30714,N30715,N30716,N30717,N30718,
N30719,N30720,N30721,N30722,N30723,N30724,N30725,N30726,N30727,N30728,
N30729,N30730,N30731,N30732,N30733,N30734,N30735,N30736,N30737,N30738,
N30739,N30740,N30741,N30742,N30743,N30744,N30745,N30746,N30747,N30748,
N30749,N30750,N30751,N30752,N30753,N30754,N30755,N30756,N30757,N30758,
N30759,N30760,N30761,N30762,N30763,N30764,N30765,N30766,N30767,N30768,
N30769,N30770,N30771,N30772,N30773,N30774,N30775,N30776,N30777,N30778,
N30779,N30780,N30781,N30782,N30783,N30784,N30785,N30786,N30787,N30788,
N30789,N30790,N30791,N30792,N30793,N30794,N30795,N30796,N30797,N30798,
N30799,N30800,N30801,N30802,N30803,N30804,N30805,N30806,N30807,N30808,
N30809,N30810,N30811,N30812,N30813,N30814,N30815,N30816,N30817,N30818,
N30819,N30820,N30821,N30822,N30823,N30824,N30825,N30826,N30827,N30828,
N30829,N30830,N30831,N30832,N30833,N30834,N30835,N30836,N30837,N30838,
N30839,N30840,N30841,N30842,N30843,N30844,N30845,N30846,N30847,N30848,
N30849,N30850,N30851,N30852,N30853,N30854,N30855,N30856,N30857,N30858,
N30859,N30860,N30861,N30862,N30863,N30864,N30865,N30866,N30867,N30868,
N30869,N30870,N30871,N30872,N30873,N30874,N30875,N30876,N30877,N30878,
N30879,N30880,N30881,N30882,N30883,N30884,N30885,N30886,N30887,N30888,
N30889,N30890,N30891,N30892,N30893,N30894,N30895,N30896,N30897,N30898,
N30899,N30900,N30901,N30902,N30903,N30904,N30905,N30906,N30907,N30908,
N30909,N30910,N30911,N30912,N30913,N30914,N30915,N30916,N30917,N30918,
N30919,N30920,N30921,N30922,N30923,N30924,N30925,N30926,N30927,N30928,
N30929,N30930,N30931,N30932,N30933,N30934,N30935,N30936,N30937,N30938,
N30939,N30940,N30941,N30942,N30943,N30944,N30945,N30946,N30947,N30948,
N30949,N30950,N30951,N30952,N30953,N30954,N30955,N30956,N30957,N30958,
N30959,N30960,N30961,N30962,N30963,N30964,N30965,N30966,N30967,N30968,
N30969,N30970,N30971,N30972,N30973,N30974,N30975,N30976,N30977,N30978,
N30979,N30980,N30981,N30982,N30983,N30984,N30985,N30986,N30987,N30988,
N30989,N30990,N30991,N30992,N30993,N30994,N30995,N30996,N30997,N30998,
N30999,N31000,N31001,N31002,N31003,N31004,N31005,N31006,N31007,N31008,
N31009,N31010,N31011,N31012,N31013,N31014,N31015,N31016,N31017,N31018,
N31019,N31020,N31021,N31022,N31023,N31024,N31025,N31026,N31027,N31028,
N31029,N31030,N31031,N31032,N31033,N31034,N31035,N31036,N31037,N31038,
N31039,N31040,N31041,N31042,N31043,N31044,N31045,N31046,N31047,N31048,
N31049,N31050,N31051,N31052,N31053,N31054,N31055,N31056,N31057,N31058,
N31059,N31060,N31061,N31062,N31063,N31064,N31065,N31066,N31067,N31068,
N31069,N31070,N31071,N31072,N31073,N31074,N31075,N31076,N31077,N31078,
N31079,N31080,N31081,N31082,N31083,N31084,N31085,N31086,N31087,N31088,
N31089,N31090,N31091,N31092,N31093,N31094,N31095,N31096,N31097,N31098,
N31099,N31100,N31101,N31102,N31103,N31104,N31105,N31106,N31107,N31108,
N31109,N31110,N31111,N31112,N31113,N31114,N31115,N31116,N31117,N31118,
N31119,N31120,N31121,N31122,N31123,N31124,N31125,N31126,N31127,N31128,
N31129,N31130,N31131,N31132,N31133,N31134,N31135,N31136,N31137,N31138,
N31139,N31140,N31141,N31142,N31143,N31144,N31145,N31146,N31147,N31148,
N31149,N31150,N31151,N31152,N31153,N31154,N31155,N31156,N31157,N31158,
N31159,N31160,N31161,N31162,N31163,N31164,N31165,N31166,N31167,N31168,
N31169,N31170,N31171,N31172,N31173,N31174,N31175,N31176,N31177,N31178,
N31179,N31180,N31181,N31182,N31183,N31184,N31185,N31186,N31187,N31188,
N31189,N31190,N31191,N31192,N31193,N31194,N31195,N31196,N31197,N31198,
N31199,N31200,N31201,N31202,N31203,N31204,N31205,N31206,N31207,N31208,
N31209,N31210,N31211,N31212,N31213,N31214,N31215,N31216,N31217,N31218,
N31219,N31220,N31221,N31222,N31223,N31224,N31225,N31226,N31227,N31228,
N31229,N31230,N31231,N31232,N31233,N31234,N31235,N31236,N31237,N31238,
N31239,N31240,N31241,N31242,N31243,N31244,N31245,N31246,N31247,N31248,
N31249,N31250,N31251,N31252,N31253,N31254,N31255,N31256,N31257,N31258,
N31259,N31260,N31261,N31262,N31263,N31264,N31265,N31266,N31267,N31268,
N31269,N31270,N31271,N31272,N31273,N31274,N31275,N31276,N31277,N31278,
N31279,N31280,N31281,N31282,N31283,N31284,N31285,N31286,N31287,N31288,
N31289,N31290,N31291,N31292,N31293,N31294,N31295,N31296,N31297,N31298,
N31299,N31300,N31301,N31302,N31303,N31304,N31305,N31306,N31307,N31308,
N31309,N31310,N31311,N31312,N31313,N31314,N31315,N31316,N31317,N31318,
N31319,N31320,N31321,N31322,N31323,N31324,N31325,N31326,N31327,N31328,
N31329,N31330,N31331,N31332,N31333,N31334,N31335,N31336,N31337,N31338,
N31339,N31340,N31341,N31342,N31343,N31344,N31345,N31346,N31347,N31348,
N31349,N31350,N31351,N31352,N31353,N31354,N31355,N31356,N31357,N31358,
N31359,N31360,N31361,N31362,N31363,N31364,N31365,N31366,N31367,N31368,
N31369,N31370,N31371,N31372,N31373,N31374,N31375,N31376,N31377,N31378,
N31379,N31380,N31381,N31382,N31383,N31384,N31385,N31386,N31387,N31388,
N31389,N31390,N31391,N31392,N31393,N31394,N31395,N31396,N31397,N31398,
N31399,N31400,N31401,N31402,N31403,N31404,N31405,N31406,N31407,N31408,
N31409,N31410,N31411,N31412,N31413,N31414,N31415,N31416,N31417,N31418,
N31419,N31420,N31421,N31422,N31423,N31424,N31425,N31426,N31427,N31428,
N31429,N31430,N31431,N31432,N31433,N31434,N31435,N31436,N31437,N31438,
N31439,N31440,N31441,N31442,N31443,N31444,N31445,N31446,N31447,N31448,
N31449,N31450,N31451,N31452,N31453,N31454,N31455,N31456,N31457,N31458,
N31459,N31460,N31461,N31462,N31463,N31464,N31465,N31466,N31467,N31468,
N31469,N31470,N31471,N31472,N31473,N31474,N31475,N31476,N31477,N31478,
N31479,N31480,N31481,N31482,N31483,N31484,N31485,N31486,N31487,N31488,
N31489,N31490,N31491,N31492,N31493,N31494,N31495,N31496,N31497,N31498,
N31499,N31500,N31501,N31502,N31503,N31504,N31505,N31506,N31507,N31508,
N31509,N31510,N31511,N31512,N31513,N31514,N31515,N31516,N31517,N31518,
N31519,N31520,N31521,N31522,N31523,N31524,N31525,N31526,N31527,N31528,
N31529,N31530,N31531,N31532,N31533,N31534,N31535,N31536,N31537,N31538,
N31539,N31540,N31541,N31542,N31543,N31544,N31545,N31546,N31547,N31548,
N31549,N31550,N31551,N31552,N31553,N31554,N31555,N31556,N31557,N31558,
N31559,N31560,N31561,N31562,N31563,N31564,N31565,N31566,N31567,N31568,
N31569,N31570,N31571,N31572,N31573,N31574,N31575,N31576,N31577,N31578,
N31579,N31580,N31581,N31582,N31583,N31584,N31585,N31586,N31587,N31588,
N31589,N31590,N31591,N31592,N31593,N31594,N31595,N31596,N31597,N31598,
N31599,N31600,N31601,N31602,N31603,N31604,N31605,N31606,N31607,N31608,
N31609,N31610,N31611,N31612,N31613,N31614,N31615,N31616,N31617,N31618,
N31619,N31620,N31621,N31622,N31623,N31624,N31625,N31626,N31627,N31628,
N31629,N31630,N31631,N31632,N31633,N31634,N31635,N31636,N31637,N31638,
N31639,N31640,N31641,N31642,N31643,N31644,N31645,N31646,N31647,N31648,
N31649,N31650,N31651,N31652,N31653,N31654,N31655,N31656,N31657,N31658,
N31659,N31660,N31661,N31662,N31663,N31664,N31665,N31666,N31667,N31668,
N31669,N31670,N31671,N31672,N31673,N31674,N31675,N31676,N31677,N31678,
N31679,N31680,N31681,N31682,N31683,N31684,N31685,N31686,N31687,N31688,
N31689,N31690,N31691,N31692,N31693,N31694,N31695,N31696,N31697,N31698,
N31699,N31700,N31701,N31702,N31703,N31704,N31705,N31706,N31707,N31708,
N31709,N31710,N31711,N31712,N31713,N31714,N31715,N31716,N31717,N31718,
N31719,N31720,N31721,N31722,N31723,N31724,N31725,N31726,N31727,N31728,
N31729,N31730,N31731,N31732,N31733,N31734,N31735,N31736,N31737,N31738,
N31739,N31740,N31741,N31742,N31743,N31744,N31745,N31746,N31747,N31748,
N31749,N31750,N31751,N31752,N31753,N31754,N31755,N31756,N31757,N31758,
N31759,N31760,N31761,N31762,N31763,N31764,N31765,N31766,N31767,N31768,
N31769,N31770,N31771,N31772,N31773,N31774,N31775,N31776,N31777,N31778,
N31779,N31780,N31781,N31782,N31783,N31784,N31785,N31786,N31787,N31788,
N31789,N31790,N31791,N31792,N31793,N31794,N31795,N31796,N31797,N31798,
N31799,N31800,N31801,N31802,N31803,N31804,N31805,N31806,N31807,N31808,
N31809,N31810,N31811,N31812,N31813,N31814,N31815,N31816,N31817,N31818,
N31819,N31820,N31821,N31822,N31823,N31824,N31825,N31826,N31827,N31828,
N31829,N31830,N31831,N31832,N31833,N31834,N31835,N31836,N31837,N31838,
N31839,N31840,N31841,N31842,N31843,N31844,N31845,N31846,N31847,N31848,
N31849,N31850,N31851,N31852,N31853,N31854,N31855,N31856,N31857,N31858,
N31859,N31860,N31861,N31862,N31863,N31864,N31865,N31866,N31867,N31868,
N31869,N31870,N31871,N31872,N31873,N31874,N31875,N31876,N31877,N31878,
N31879,N31880,N31881,N31882,N31883,N31884,N31885,N31886,N31887,N31888,
N31889,N31890,N31891,N31892,N31893,N31894,N31895,N31896,N31897,N31898,
N31899,N31900,N31901,N31902,N31903,N31904,N31905,N31906,N31907,N31908,
N31909,N31910,N31911,N31912,N31913,N31914,N31915,N31916,N31917,N31918,
N31919,N31920,N31921,N31922,N31923,N31924,N31925,N31926,N31927,N31928,
N31929,N31930,N31931,N31932,N31933,N31934,N31935,N31936,N31937,N31938,
N31939,N31940,N31941,N31942,N31943,N31944,N31945,N31946,N31947,N31948,
N31949,N31950,N31951,N31952,N31953,N31954,N31955,N31956,N31957,N31958,
N31959,N31960,N31961,N31962,N31963,N31964,N31965,N31966,N31967,N31968,
N31969,N31970,N31971,N31972,N31973,N31974,N31975,N31976,N31977,N31978,
N31979,N31980,N31981,N31982,N31983,N31984,N31985,N31986,N31987,N31988,
N31989,N31990,N31991,N31992,N31993,N31994,N31995,N31996,N31997,N31998,
N31999,N32000,N32001,N32002,N32003,N32004,N32005,N32006,N32007,N32008,
N32009,N32010,N32011,N32012,N32013,N32014,N32015,N32016,N32017,N32018,
N32019,N32020,N32021,N32022,N32023,N32024,N32025,N32026,N32027,N32028,
N32029,N32030,N32031,N32032,N32033,N32034,N32035,N32036,N32037,N32038,
N32039,N32040,N32041,N32042,N32043,N32044,N32045,N32046,N32047,N32048,
N32049,N32050,N32051,N32052,N32053,N32054,N32055,N32056,N32057,N32058,
N32059,N32060,N32061,N32062,N32063,N32064,N32065,N32066,N32067,N32068,
N32069,N32070,N32071,N32072,N32073,N32074,N32075,N32076,N32077,N32078,
N32079,N32080,N32081,N32082,N32083,N32084,N32085,N32086,N32087,N32088,
N32089,N32090,N32091,N32092,N32093,N32094,N32095,N32096,N32097,N32098,
N32099,N32100,N32101,N32102,N32103,N32104,N32105,N32106,N32107,N32108,
N32109,N32110,N32111,N32112,N32113,N32114,N32115,N32116,N32117,N32118,
N32119,N32120,N32121,N32122,N32123,N32124,N32125,N32126,N32127,N32128,
N32129,N32130,N32131,N32132,N32133,N32134,N32135,N32136,N32137,N32138,
N32139,N32140,N32141,N32142,N32143,N32144,N32145,N32146,N32147,N32148,
N32149,N32150,N32151,N32152,N32153,N32154,N32155,N32156,N32157,N32158,
N32159,N32160,N32161,N32162,N32163,N32164,N32165,N32166,N32167,N32168,
N32169,N32170,N32171,N32172,N32173,N32174,N32175,N32176,N32177,N32178,
N32179,N32180,N32181,N32182,N32183,N32184,N32185,N32186,N32187,N32188,
N32189,N32190,N32191,N32192,N32193,N32194,N32195,N32196,N32197,N32198,
N32199,N32200,N32201,N32202,N32203,N32204,N32205,N32206,N32207,N32208,
N32209,N32210,N32211,N32212,N32213,N32214,N32215,N32216,N32217,N32218,
N32219,N32220,N32221,N32222,N32223,N32224,N32225,N32226,N32227,N32228,
N32229,N32230,N32231,N32232,N32233,N32234,N32235,N32236,N32237,N32238,
N32239,N32240,N32241,N32242,N32243,N32244,N32245,N32246,N32247,N32248,
N32249,N32250,N32251,N32252,N32253,N32254,N32255,N32256,N32257,N32258,
N32259,N32260,N32261,N32262,N32263,N32264,N32265,N32266,N32267,N32268,
N32269,N32270,N32271,N32272,N32273,N32274,N32275,N32276,N32277,N32278,
N32279,N32280,N32281,N32282,N32283,N32284,N32285,N32286,N32287,N32288,
N32289,N32290,N32291,N32292,N32293,N32294,N32295,N32296,N32297,N32298,
N32299,N32300,N32301,N32302,N32303,N32304,N32305,N32306,N32307,N32308,
N32309,N32310,N32311,N32312,N32313,N32314,N32315,N32316,N32317,N32318,
N32319,N32320,N32321,N32322,N32323,N32324,N32325,N32326,N32327,N32328,
N32329,N32330,N32331,N32332,N32333,N32334,N32335,N32336,N32337,N32338,
N32339,N32340,N32341,N32342,N32343,N32344,N32345,N32346,N32347,N32348,
N32349,N32350,N32351,N32352,N32353,N32354,N32355,N32356,N32357,N32358,
N32359,N32360,N32361,N32362,N32363,N32364,N32365,N32366,N32367,N32368,
N32369,N32370,N32371,N32372,N32373,N32374,N32375,N32376,N32377,N32378,
N32379,N32380,N32381,N32382,N32383,N32384,N32385,N32386,N32387,N32388,
N32389,N32390,N32391,N32392,N32393,N32394,N32395,N32396,N32397,N32398,
N32399,N32400,N32401,N32402,N32403,N32404,N32405,N32406,N32407,N32408,
N32409,N32410,N32411,N32412,N32413,N32414,N32415,N32416,N32417,N32418,
N32419,N32420,N32421,N32422,N32423,N32424,N32425,N32426,N32427,N32428,
N32429,N32430,N32431,N32432,N32433,N32434,N32435,N32436,N32437,N32438,
N32439,N32440,N32441,N32442,N32443,N32444,N32445,N32446,N32447,N32448,
N32449,N32450,N32451,N32452,N32453,N32454,N32455,N32456,N32457,N32458,
N32459,N32460,N32461,N32462,N32463,N32464,N32465,N32466,N32467,N32468,
N32469,N32470,N32471,N32472,N32473,N32474,N32475,N32476,N32477,N32478,
N32479,N32480,N32481,N32482,N32483,N32484,N32485,N32486,N32487,N32488,
N32489,N32490,N32491,N32492,N32493,N32494,N32495,N32496,N32497,N32498,
N32499,N32500,N32501,N32502,N32503,N32504,N32505,N32506,N32507,N32508,
N32509,N32510,N32511,N32512,N32513,N32514,N32515,N32516,N32517,N32518,
N32519,N32520,N32521,N32522,N32523,N32524,N32525,N32526,N32527,N32528,
N32529,N32530,N32531,N32532,N32533,N32534,N32535,N32536,N32537,N32538,
N32539,N32540,N32541,N32542,N32543,N32544,N32545,N32546,N32547,N32548,
N32549,N32550,N32551,N32552,N32553,N32554,N32555,N32556,N32557,N32558,
N32559,N32560,N32561,N32562,N32563,N32564,N32565,N32566,N32567,N32568,
N32569,N32570,N32571,N32572,N32573,N32574,N32575,N32576,N32577,N32578,
N32579,N32580,N32581,N32582,N32583,N32584,N32585,N32586,N32587,N32588,
N32589,N32590,N32591,N32592,N32593,N32594,N32595,N32596,N32597,N32598,
N32599,N32600,N32601,N32602,N32603,N32604,N32605,N32606,N32607,N32608,
N32609,N32610,N32611,N32612,N32613,N32614,N32615,N32616,N32617,N32618,
N32619,N32620,N32621,N32622,N32623,N32624,N32625,N32626,N32627,N32628,
N32629,N32630,N32631,N32632,N32633,N32634,N32635,N32636,N32637,N32638,
N32639,N32640,N32641,N32642,N32643,N32644,N32645,N32646,N32647,N32648,
N32649,N32650,N32651,N32652,N32653,N32654,N32655,N32656,N32657,N32658,
N32659,N32660,N32661,N32662,N32663,N32664,N32665,N32666,N32667,N32668,
N32669,N32670,N32671,N32672,N32673,N32674,N32675,N32676,N32677,N32678,
N32679,N32680,N32681,N32682,N32683,N32684,N32685,N32686,N32687,N32688,
N32689,N32690,N32691,N32692,N32693,N32694,N32695,N32696,N32697,N32698,
N32699,N32700,N32701,N32702,N32703,N32704,N32705,N32706,N32707,N32708,
N32709,N32710,N32711,N32712,N32713,N32714,N32715,N32716,N32717,N32718,
N32719,N32720,N32721,N32722,N32723,N32724,N32725,N32726,N32727,N32728,
N32729,N32730,N32731,N32732,N32733,N32734,N32735,N32736,N32737,N32738,
N32739,N32740,N32741,N32742,N32743,N32744,N32745,N32746,N32747,N32748,
N32749,N32750,N32751,N32752,N32753,N32754,N32755,N32756,N32757,N32758,
N32759,N32760,N32761,N32762,N32763,N32764,N32765,N32766,N32767,N32768,
N32769,N32770,N32771,N32772,N32773,N32774,N32775,N32776,N32777,N32778,
N32779,N32780,N32781,N32782,N32783,N32784,N32785,N32786,N32787,N32788,
N32789,N32790,N32791,N32792,N32793,N32794,N32795,N32796,N32797,N32798,
N32799,N32800,N32801,N32802,N32803,N32804,N32805,N32806,N32807,N32808,
N32809,N32810,N32811,N32812,N32813,N32814,N32815,N32816,N32817,N32818,
N32819,N32820,N32821,N32822,N32823,N32824,N32825,N32826,N32827,N32828,
N32829,N32830,N32831,N32832,N32833,N32834,N32835,N32836,N32837,N32838,
N32839,N32840,N32841,N32842,N32843,N32844,N32845,N32846,N32847,N32848,
N32849,N32850,N32851,N32852,N32853,N32854,N32855,N32856,N32857,N32858,
N32859,N32860,N32861,N32862,N32863,N32864,N32865,N32866,N32867,N32868,
N32869,N32870,N32871,N32872,N32873,N32874,N32875,N32876,N32877,N32878,
N32879,N32880,N32881,N32882,N32883,N32884,N32885,N32886,N32887,N32888,
N32889,N32890,N32891,N32892,N32893,N32894,N32895,N32896,N32897,N32898,
N32899,N32900,N32901,N32902,N32903,N32904,N32905,N32906,N32907,N32908,
N32909,N32910,N32911,N32912,N32913,N32914,N32915,N32916,N32917,N32918,
N32919,N32920,N32921,N32922,N32923,N32924,N32925,N32926,N32927,N32928,
N32929,N32930,N32931,N32932,N32933,N32934,N32935,N32936,N32937,N32938,
N32939,N32940,N32941,N32942,N32943,N32944,N32945,N32946,N32947,N32948,
N32949,N32950,N32951,N32952,N32953,N32954,N32955,N32956,N32957,N32958,
N32959,N32960,N32961,N32962,N32963,N32964,N32965,N32966,N32967,N32968,
N32969,N32970,N32971,N32972,N32973,N32974,N32975,N32976,N32977,N32978,
N32979,N32980,N32981,N32982,N32983,N32984,N32985,N32986,N32987,N32988,
N32989,N32990,N32991,N32992,N32993,N32994,N32995,N32996,N32997,N32998,
N32999,N33000,N33001,N33002,N33003,N33004,N33005,N33006,N33007,N33008,
N33009,N33010,N33011,N33012,N33013,N33014,N33015,N33016,N33017,N33018,
N33019,N33020,N33021,N33022,N33023,N33024,N33025,N33026,N33027,N33028,
N33029,N33030,N33031,N33032,N33033,N33034,N33035,N33036,N33037,N33038,
N33039,N33040,N33041,N33042,N33043,N33044,N33045,N33046,N33047,N33048,
N33049,N33050,N33051,N33052,N33053,N33054,N33055,N33056,N33057,N33058,
N33059,N33060,N33061,N33062,N33063,N33064,N33065,N33066,N33067,N33068,
N33069,N33070,N33071,N33072,N33073,N33074,N33075,N33076,N33077,N33078,
N33079,N33080,N33081,N33082,N33083,N33084,N33085,N33086,N33087,N33088,
N33089,N33090,N33091,N33092,N33093,N33094,N33095,N33096,N33097,N33098,
N33099,N33100,N33101,N33102,N33103,N33104,N33105,N33106,N33107,N33108,
N33109,N33110,N33111,N33112,N33113,N33114,N33115,N33116,N33117,N33118,
N33119,N33120,N33121,N33122,N33123,N33124,N33125,N33126,N33127,N33128,
N33129,N33130,N33131,N33132,N33133,N33134,N33135,N33136,N33137,N33138,
N33139,N33140,N33141,N33142,N33143,N33144,N33145,N33146,N33147,N33148,
N33149,N33150,N33151,N33152,N33153,N33154,N33155,N33156,N33157,N33158,
N33159,N33160,N33161,N33162,N33163,N33164,N33165,N33166,N33167,N33168,
N33169,N33170,N33171,N33172,N33173,N33174,N33175,N33176,N33177,N33178,
N33179,N33180,N33181,N33182,N33183,N33184,N33185,N33186,N33187,N33188,
N33189,N33190,N33191,N33192,N33193,N33194,N33195,N33196,N33197,N33198,
N33199,N33200,N33201,N33202,N33203,N33204,N33205,N33206,N33207,N33208,
N33209,N33210,N33211,N33212,N33213,N33214,N33215,N33216,N33217,N33218,
N33219,N33220,N33221,N33222,N33223,N33224,N33225,N33226,N33227,N33228,
N33229,N33230,N33231,N33232,N33233,N33234,N33235,N33236,N33237,N33238,
N33239,N33240,N33241,N33242,N33243,N33244,N33245,N33246,N33247,N33248,
N33249,N33250,N33251,N33252,N33253,N33254,N33255,N33256,N33257,N33258,
N33259,N33260,N33261,N33262,N33263,N33264,N33265,N33266,N33267,N33268,
N33269,N33270,N33271,N33272,N33273,N33274,N33275,N33276,N33277,N33278,
N33279,N33280,N33281,N33282,N33283,N33284,N33285,N33286,N33287,N33288,
N33289,N33290,N33291,N33292,N33293,N33294,N33295,N33296,N33297,N33298,
N33299,N33300,N33301,N33302,N33303,N33304,N33305,N33306,N33307,N33308,
N33309,N33310,N33311,N33312,N33313,N33314,N33315,N33316,N33317,N33318,
N33319,N33320,N33321,N33322,N33323,N33324,N33325,N33326,N33327,N33328,
N33329,N33330,N33331,N33332,N33333,N33334,N33335,N33336,N33337,N33338,
N33339,N33340,N33341,N33342,N33343,N33344,N33345,N33346,N33347,N33348,
N33349,N33350,N33351,N33352,N33353,N33354,N33355,N33356,N33357,N33358,
N33359,N33360,N33361,N33362,N33363,N33364,N33365,N33366,N33367,N33368,
N33369,N33370,N33371,N33372,N33373,N33374,N33375,N33376,N33377,N33378,
N33379,N33380,N33381,N33382,N33383,N33384,N33385,N33386,N33387,N33388,
N33389,N33390,N33391,N33392,N33393,N33394,N33395,N33396,N33397,N33398,
N33399,N33400,N33401,N33402,N33403,N33404,N33405,N33406,N33407,N33408,
N33409,N33410,N33411,N33412,N33413,N33414,N33415,N33416,N33417,N33418,
N33419,N33420,N33421,N33422,N33423,N33424,N33425,N33426,N33427,N33428,
N33429,N33430,N33431,N33432,N33433,N33434,N33435,N33436,N33437,N33438,
N33439,N33440,N33441,N33442,N33443,N33444,N33445,N33446,N33447,N33448,
N33449,N33450,N33451,N33452,N33453,N33454,N33455,N33456,N33457,N33458,
N33459,N33460,N33461,N33462,N33463,N33464,N33465,N33466,N33467,N33468,
N33469,N33470,N33471,N33472,N33473,N33474,N33475,N33476,N33477,N33478,
N33479,N33480,N33481,N33482,N33483,N33484,N33485,N33486,N33487,N33488,
N33489,N33490,N33491,N33492,N33493,N33494,N33495,N33496,N33497,N33498,
N33499,N33500,N33501,N33502,N33503,N33504,N33505,N33506,N33507,N33508,
N33509,N33510,N33511,N33512,N33513,N33514,N33515,N33516,N33517,N33518,
N33519,N33520,N33521,N33522,N33523,N33524,N33525,N33526,N33527,N33528,
N33529,N33530,N33531,N33532,N33533,N33534,N33535,N33536,N33537,N33538,
N33539,N33540,N33541,N33542,N33543,N33544,N33545,N33546,N33547,N33548,
N33549,N33550,N33551,N33552,N33553,N33554,N33555,N33556,N33557,N33558,
N33559,N33560,N33561,N33562,N33563,N33564,N33565,N33566,N33567,N33568,
N33569,N33570,N33571,N33572,N33573,N33574,N33575,N33576,N33577,N33578,
N33579,N33580,N33581,N33582,N33583,N33584,N33585,N33586,N33587,N33588,
N33589,N33590,N33591,N33592,N33593,N33594,N33595,N33596,N33597,N33598,
N33599,N33600,N33601,N33602,N33603,N33604,N33605,N33606,N33607,N33608,
N33609,N33610,N33611,N33612,N33613,N33614,N33615,N33616,N33617,N33618,
N33619,N33620,N33621,N33622,N33623,N33624,N33625,N33626,N33627,N33628,
N33629,N33630,N33631,N33632,N33633,N33634,N33635,N33636,N33637,N33638,
N33639,N33640,N33641,N33642,N33643,N33644,N33645,N33646,N33647,N33648,
N33649,N33650,N33651,N33652,N33653,N33654,N33655,N33656,N33657,N33658,
N33659,N33660,N33661,N33662,N33663,N33664,N33665,N33666,N33667,N33668,
N33669,N33670,N33671,N33672,N33673,N33674,N33675,N33676,N33677,N33678,
N33679,N33680,N33681,N33682,N33683,N33684,N33685,N33686,N33687,N33688,
N33689,N33690,N33691,N33692,N33693,N33694,N33695,N33696,N33697,N33698,
N33699,N33700,N33701,N33702,N33703,N33704,N33705,N33706,N33707,N33708,
N33709,N33710,N33711,N33712,N33713,N33714,N33715,N33716,N33717,N33718,
N33719,N33720,N33721,N33722,N33723,N33724,N33725,N33726,N33727,N33728,
N33729,N33730,N33731,N33732,N33733,N33734,N33735,N33736,N33737,N33738,
N33739,N33740,N33741,N33742,N33743,N33744,N33745,N33746,N33747,N33748,
N33749,N33750,N33751,N33752,N33753,N33754,N33755,N33756,N33757,N33758,
N33759,N33760,N33761,N33762,N33763,N33764,N33765,N33766,N33767,N33768,
N33769,N33770,N33771,N33772,N33773,N33774,N33775,N33776,N33777,N33778,
N33779,N33780,N33781,N33782,N33783,N33784,N33785,N33786,N33787,N33788,
N33789,N33790,N33791,N33792,N33793,N33794,N33795,N33796,N33797,N33798,
N33799,N33800,N33801,N33802,N33803,N33804,N33805,N33806,N33807,N33808,
N33809,N33810,N33811,N33812,N33813,N33814,N33815,N33816,N33817,N33818,
N33819,N33820,N33821,N33822,N33823,N33824,N33825,N33826,N33827,N33828,
N33829,N33830,N33831,N33832,N33833,N33834,N33835,N33836,N33837,N33838,
N33839,N33840,N33841,N33842,N33843,N33844,N33845,N33846,N33847,N33848,
N33849,N33850,N33851,N33852,N33853,N33854,N33855,N33856,N33857,N33858,
N33859,N33860,N33861,N33862,N33863,N33864,N33865,N33866,N33867,N33868,
N33869,N33870,N33871,N33872,N33873,N33874,N33875,N33876,N33877,N33878,
N33879,N33880,N33881,N33882,N33883,N33884,N33885,N33886,N33887,N33888,
N33889,N33890,N33891,N33892,N33893,N33894,N33895,N33896,N33897,N33898,
N33899,N33900,N33901,N33902,N33903,N33904,N33905,N33906,N33907,N33908,
N33909,N33910,N33911,N33912,N33913,N33914,N33915,N33916,N33917,N33918,
N33919,N33920,N33921,N33922,N33923,N33924,N33925,N33926,N33927,N33928,
N33929,N33930,N33931,N33932,N33933,N33934,N33935,N33936,N33937,N33938,
N33939,N33940,N33941,N33942,N33943,N33944,N33945,N33946,N33947,N33948,
N33949,N33950,N33951,N33952,N33953,N33954,N33955,N33956,N33957,N33958,
N33959,N33960,N33961,N33962,N33963,N33964,N33965,N33966,N33967,N33968,
N33969,N33970,N33971,N33972,N33973,N33974,N33975,N33976,N33977,N33978,
N33979,N33980,N33981,N33982,N33983,N33984,N33985,N33986,N33987,N33988,
N33989,N33990,N33991,N33992,N33993,N33994,N33995,N33996,N33997,N33998,
N33999,N34000,N34001,N34002,N34003,N34004,N34005,N34006,N34007,N34008,
N34009,N34010,N34011,N34012,N34013,N34014,N34015,N34016,N34017,N34018,
N34019,N34020,N34021,N34022,N34023,N34024,N34025,N34026,N34027,N34028,
N34029,N34030,N34031,N34032,N34033,N34034,N34035,N34036,N34037,N34038,
N34039,N34040,N34041,N34042,N34043,N34044,N34045,N34046,N34047,N34048,
N34049,N34050,N34051,N34052,N34053,N34054,N34055,N34056,N34057,N34058,
N34059,N34060,N34061,N34062,N34063,N34064,N34065,N34066,N34067,N34068,
N34069,N34070,N34071,N34072,N34073,N34074,N34075,N34076,N34077,N34078,
N34079,N34080,N34081,N34082,N34083,N34084,N34085,N34086,N34087,N34088,
N34089,N34090,N34091,N34092,N34093,N34094,N34095,N34096,N34097,N34098,
N34099,N34100,N34101,N34102,N34103,N34104,N34105,N34106,N34107,N34108,
N34109,N34110,N34111,N34112,N34113,N34114,N34115,N34116,N34117,N34118,
N34119,N34120,N34121,N34122,N34123,N34124,N34125,N34126,N34127,N34128,
N34129,N34130,N34131,N34132,N34133,N34134,N34135,N34136,N34137,N34138,
N34139,N34140,N34141,N34142,N34143,N34144,N34145,N34146,N34147,N34148,
N34149,N34150,N34151,N34152,N34153,N34154,N34155,N34156,N34157,N34158,
N34159,N34160,N34161,N34162,N34163,N34164,N34165,N34166,N34167,N34168,
N34169,N34170,N34171,N34172,N34173,N34174,N34175,N34176,N34177,N34178,
N34179,N34180,N34181,N34182,N34183,N34184,N34185,N34186,N34187,N34188,
N34189,N34190,N34191,N34192,N34193,N34194,N34195,N34196,N34197,N34198,
N34199,N34200,N34201,N34202,N34203,N34204,N34205,N34206,N34207,N34208,
N34209,N34210,N34211,N34212,N34213,N34214,N34215,N34216,N34217,N34218,
N34219,N34220,N34221,N34222,N34223,N34224,N34225,N34226,N34227,N34228,
N34229,N34230,N34231,N34232,N34233,N34234,N34235,N34236,N34237,N34238,
N34239,N34240,N34241,N34242,N34243,N34244,N34245,N34246,N34247,N34248,
N34249,N34250,N34251,N34252,N34253,N34254,N34255,N34256,N34257,N34258,
N34259,N34260,N34261,N34262,N34263,N34264,N34265,N34266,N34267,N34268,
N34269,N34270,N34271,N34272,N34273,N34274,N34275,N34276,N34277,N34278,
N34279,N34280,N34281,N34282,N34283,N34284,N34285,N34286,N34287,N34288,
N34289,N34290,N34291,N34292,N34293,N34294,N34295,N34296,N34297,N34298,
N34299,N34300,N34301,N34302,N34303,N34304,N34305,N34306,N34307,N34308,
N34309,N34310,N34311,N34312,N34313,N34314,N34315,N34316,N34317,N34318,
N34319,N34320,N34321,N34322,N34323,N34324,N34325,N34326,N34327,N34328,
N34329,N34330,N34331,N34332,N34333,N34334,N34335,N34336,N34337,N34338,
N34339,N34340,N34341,N34342,N34343,N34344,N34345,N34346,N34347,N34348,
N34349,N34350,N34351,N34352,N34353,N34354,N34355,N34356,N34357,N34358,
N34359,N34360,N34361,N34362,N34363,N34364,N34365,N34366,N34367,N34368,
N34369,N34370,N34371,N34372,N34373,N34374,N34375,N34376,N34377,N34378,
N34379,N34380,N34381,N34382,N34383,N34384,N34385,N34386,N34387,N34388,
N34389,N34390,N34391,N34392,N34393,N34394,N34395,N34396,N34397,N34398,
N34399,N34400,N34401,N34402,N34403,N34404,N34405,N34406,N34407,N34408,
N34409,N34410,N34411,N34412,N34413,N34414,N34415,N34416,N34417,N34418,
N34419,N34420,N34421,N34422,N34423,N34424,N34425,N34426,N34427,N34428,
N34429,N34430,N34431,N34432,N34433,N34434,N34435,N34436,N34437,N34438,
N34439,N34440,N34441,N34442,N34443,N34444,N34445,N34446,N34447,N34448,
N34449,N34450,N34451,N34452,N34453,N34454,N34455,N34456,N34457,N34458,
N34459,N34460,N34461,N34462,N34463,N34464,N34465,N34466,N34467,N34468,
N34469,N34470,N34471,N34472,N34473,N34474,N34475,N34476,N34477,N34478,
N34479,N34480,N34481,N34482,N34483,N34484,N34485,N34486,N34487,N34488,
N34489,N34490,N34491,N34492,N34493,N34494,N34495,N34496,N34497,N34498,
N34499,N34500,N34501,N34502,N34503,N34504,N34505,N34506,N34507,N34508,
N34509,N34510,N34511,N34512,N34513,N34514,N34515,N34516,N34517,N34518,
N34519,N34520,N34521,N34522,N34523,N34524,N34525,N34526,N34527,N34528,
N34529,N34530,N34531,N34532,N34533,N34534,N34535,N34536,N34537,N34538,
N34539,N34540,N34541,N34542,N34543,N34544,N34545,N34546,N34547,N34548,
N34549,N34550,N34551,N34552,N34553,N34554,N34555,N34556,N34557,N34558,
N34559,N34560,N34561,N34562,N34563,N34564,N34565,N34566,N34567,N34568,
N34569,N34570,N34571,N34572,N34573,N34574,N34575,N34576,N34577,N34578,
N34579,N34580,N34581,N34582,N34583,N34584,N34585,N34586,N34587,N34588,
N34589,N34590,N34591,N34592,N34593,N34594,N34595,N34596,N34597,N34598,
N34599,N34600,N34601,N34602,N34603,N34604,N34605,N34606,N34607,N34608,
N34609,N34610,N34611,N34612,N34613,N34614,N34615,N34616,N34617,N34618,
N34619,N34620,N34621,N34622,N34623,N34624,N34625,N34626,N34627,N34628,
N34629,N34630,N34631,N34632,N34633,N34634,N34635,N34636,N34637,N34638,
N34639,N34640,N34641,N34642,N34643,N34644,N34645,N34646,N34647,N34648,
N34649,N34650,N34651,N34652,N34653,N34654,N34655,N34656,N34657,N34658,
N34659,N34660,N34661,N34662,N34663,N34664,N34665,N34666,N34667,N34668,
N34669,N34670,N34671,N34672,N34673,N34674,N34675,N34676,N34677,N34678,
N34679,N34680,N34681,N34682,N34683,N34684,N34685,N34686,N34687,N34688,
N34689,N34690,N34691,N34692,N34693,N34694,N34695,N34696,N34697,N34698,
N34699,N34700,N34701,N34702,N34703,N34704,N34705,N34706,N34707,N34708,
N34709,N34710,N34711,N34712,N34713,N34714,N34715,N34716,N34717,N34718,
N34719,N34720,N34721,N34722,N34723,N34724,N34725,N34726,N34727,N34728,
N34729,N34730,N34731,N34732,N34733,N34734,N34735,N34736,N34737,N34738,
N34739,N34740,N34741,N34742,N34743,N34744,N34745,N34746,N34747,N34748,
N34749,N34750,N34751,N34752,N34753,N34754,N34755,N34756,N34757,N34758,
N34759,N34760,N34761,N34762,N34763,N34764,N34765,N34766,N34767,N34768,
N34769,N34770,N34771,N34772,N34773,N34774,N34775,N34776,N34777,N34778,
N34779,N34780,N34781,N34782,N34783,N34784,N34785,N34786,N34787,N34788,
N34789,N34790,N34791,N34792,N34793,N34794,N34795,N34796,N34797,N34798,
N34799,N34800,N34801,N34802,N34803,N34804,N34805,N34806,N34807,N34808,
N34809,N34810,N34811,N34812,N34813,N34814,N34815,N34816,N34817,N34818,
N34819,N34820,N34821,N34822,N34823,N34824,N34825,N34826,N34827,N34828,
N34829,N34830,N34831,N34832,N34833,N34834,N34835,N34836,N34837,N34838,
N34839,N34840,N34841,N34842,N34843,N34844,N34845,N34846,N34847,N34848,
N34849,N34850,N34851,N34852,N34853,N34854,N34855,N34856,N34857,N34858,
N34859,N34860,N34861,N34862,N34863,N34864,N34865,N34866,N34867,N34868,
N34869,N34870,N34871,N34872,N34873,N34874,N34875,N34876,N34877,N34878,
N34879,N34880,N34881,N34882,N34883,N34884,N34885,N34886,N34887,N34888,
N34889,N34890,N34891,N34892,N34893,N34894,N34895,N34896,N34897,N34898,
N34899,N34900,N34901,N34902,N34903,N34904,N34905,N34906,N34907,N34908,
N34909,N34910,N34911,N34912,N34913,N34914,N34915,N34916,N34917,N34918,
N34919,N34920,N34921,N34922,N34923,N34924,N34925,N34926,N34927,N34928,
N34929,N34930,N34931,N34932,N34933,N34934,N34935,N34936,N34937,N34938,
N34939,N34940,N34941,N34942,N34943,N34944,N34945,N34946,N34947,N34948,
N34949,N34950,N34951,N34952,N34953,N34954,N34955,N34956,N34957,N34958,
N34959,N34960,N34961,N34962,N34963,N34964,N34965,N34966,N34967,N34968,
N34969,N34970,N34971,N34972,N34973,N34974,N34975,N34976,N34977,N34978,
N34979,N34980,N34981,N34982,N34983,N34984,N34985,N34986,N34987,N34988,
N34989,N34990,N34991,N34992,N34993,N34994,N34995,N34996,N34997,N34998,
N34999,N35000,N35001,N35002,N35003,N35004,N35005,N35006,N35007,N35008,
N35009,N35010,N35011,N35012,N35013,N35014,N35015,N35016,N35017,N35018,
N35019,N35020,N35021,N35022,N35023,N35024,N35025,N35026,N35027,N35028,
N35029,N35030,N35031,N35032,N35033,N35034,N35035,N35036,N35037,N35038,
N35039,N35040,N35041,N35042,N35043,N35044,N35045,N35046,N35047,N35048,
N35049,N35050,N35051,N35052,N35053,N35054,N35055,N35056,N35057,N35058,
N35059,N35060,N35061,N35062,N35063,N35064,N35065,N35066,N35067,N35068,
N35069,N35070,N35071,N35072,N35073,N35074,N35075,N35076,N35077,N35078,
N35079,N35080,N35081,N35082,N35083,N35084,N35085,N35086,N35087,N35088,
N35089,N35090,N35091,N35092,N35093,N35094,N35095,N35096,N35097,N35098,
N35099,N35100,N35101,N35102,N35103,N35104,N35105,N35106,N35107,N35108,
N35109,N35110,N35111,N35112,N35113,N35114,N35115,N35116,N35117,N35118,
N35119,N35120,N35121,N35122,N35123,N35124,N35125,N35126,N35127,N35128,
N35129,N35130,N35131,N35132,N35133,N35134,N35135,N35136,N35137,N35138,
N35139,N35140,N35141,N35142,N35143,N35144,N35145,N35146,N35147,N35148,
N35149,N35150,N35151,N35152,N35153,N35154,N35155,N35156,N35157,N35158,
N35159,N35160,N35161,N35162,N35163,N35164,N35165,N35166,N35167,N35168,
N35169,N35170,N35171,N35172,N35173,N35174,N35175,N35176,N35177,N35178,
N35179,N35180,N35181,N35182,N35183,N35184,N35185,N35186,N35187,N35188,
N35189,N35190,N35191,N35192,N35193,N35194,N35195,N35196,N35197,N35198,
N35199,N35200,N35201,N35202,N35203,N35204,N35205,N35206,N35207,N35208,
N35209,N35210,N35211,N35212,N35213,N35214,N35215,N35216,N35217,N35218,
N35219,N35220,N35221,N35222,N35223,N35224,N35225,N35226,N35227,N35228,
N35229,N35230,N35231,N35232,N35233,N35234,N35235,N35236,N35237,N35238,
N35239,N35240,N35241,N35242,N35243,N35244,N35245,N35246,N35247,N35248,
N35249,N35250,N35251,N35252,N35253,N35254,N35255,N35256,N35257,N35258,
N35259,N35260,N35261,N35262,N35263,N35264,N35265,N35266,N35267,N35268,
N35269,N35270,N35271,N35272,N35273,N35274,N35275,N35276,N35277,N35278,
N35279,N35280,N35281,N35282,N35283,N35284,N35285,N35286,N35287,N35288,
N35289,N35290,N35291,N35292,N35293,N35294,N35295,N35296,N35297,N35298,
N35299,N35300,N35301,N35302,N35303,N35304,N35305,N35306,N35307,N35308,
N35309,N35310,N35311,N35312,N35313,N35314,N35315,N35316,N35317,N35318,
N35319,N35320,N35321,N35322,N35323,N35324,N35325,N35326,N35327,N35328,
N35329,N35330,N35331,N35332,N35333,N35334,N35335,N35336,N35337,N35338,
N35339,N35340,N35341,N35342,N35343,N35344,N35345,N35346,N35347,N35348,
N35349,N35350,N35351,N35352,N35353,N35354,N35355,N35356,N35357,N35358,
N35359,N35360,N35361,N35362,N35363,N35364,N35365,N35366,N35367,N35368,
N35369,N35370,N35371,N35372,N35373,N35374,N35375,N35376,N35377,N35378,
N35379,N35380,N35381,N35382,N35383,N35384,N35385,N35386,N35387,N35388,
N35389,N35390,N35391,N35392,N35393,N35394,N35395,N35396,N35397,N35398,
N35399,N35400,N35401,N35402,N35403,N35404,N35405,N35406,N35407,N35408,
N35409,N35410,N35411,N35412,N35413,N35414,N35415,N35416,N35417,N35418,
N35419,N35420,N35421,N35422,N35423,N35424,N35425,N35426,N35427,N35428,
N35429,N35430,N35431,N35432,N35433,N35434,N35435,N35436,N35437,N35438,
N35439,N35440,N35441,N35442,N35443,N35444,N35445,N35446,N35447,N35448,
N35449,N35450,N35451,N35452,N35453,N35454,N35455,N35456,N35457,N35458,
N35459,N35460,N35461,N35462,N35463,N35464,N35465,N35466,N35467,N35468,
N35469,N35470,N35471,N35472,N35473,N35474,N35475,N35476,N35477,N35478,
N35479,N35480,N35481,N35482,N35483,N35484,N35485,N35486,N35487,N35488,
N35489,N35490,N35491,N35492,N35493,N35494,N35495,N35496,N35497,N35498,
N35499,N35500,N35501,N35502,N35503,N35504,N35505,N35506,N35507,N35508,
N35509,N35510,N35511,N35512,N35513,N35514,N35515,N35516,N35517,N35518,
N35519,N35520,N35521,N35522,N35523,N35524,N35525,N35526,N35527,N35528,
N35529,N35530,N35531,N35532,N35533,N35534,N35535,N35536,N35537,N35538,
N35539,N35540,N35541,N35542,N35543,N35544,N35545,N35546,N35547,N35548,
N35549,N35550,N35551,N35552,N35553,N35554,N35555,N35556,N35557,N35558,
N35559,N35560,N35561,N35562,N35563,N35564,N35565,N35566,N35567,N35568,
N35569,N35570,N35571,N35572,N35573,N35574,N35575,N35576,N35577,N35578,
N35579,N35580,N35581,N35582,N35583,N35584,N35585,N35586,N35587,N35588,
N35589,N35590,N35591,N35592,N35593,N35594,N35595,N35596,N35597,N35598,
N35599,N35600,N35601,N35602,N35603,N35604,N35605,N35606,N35607,N35608,
N35609,N35610,N35611,N35612,N35613,N35614,N35615,N35616,N35617,N35618,
N35619,N35620,N35621,N35622,N35623,N35624,N35625,N35626,N35627,N35628,
N35629,N35630,N35631,N35632,N35633,N35634,N35635,N35636,N35637,N35638,
N35639,N35640,N35641,N35642,N35643,N35644,N35645,N35646,N35647,N35648,
N35649,N35650,N35651,N35652,N35653,N35654,N35655,N35656,N35657,N35658,
N35659,N35660,N35661,N35662,N35663,N35664,N35665,N35666,N35667,N35668,
N35669,N35670,N35671,N35672,N35673,N35674,N35675,N35676,N35677,N35678,
N35679,N35680,N35681,N35682,N35683,N35684,N35685,N35686,N35687,N35688,
N35689,N35690,N35691,N35692,N35693,N35694,N35695,N35696,N35697,N35698,
N35699,N35700,N35701,N35702,N35703,N35704,N35705,N35706,N35707,N35708,
N35709,N35710,N35711,N35712,N35713,N35714,N35715,N35716,N35717,N35718,
N35719,N35720,N35721,N35722,N35723,N35724,N35725,N35726,N35727,N35728,
N35729,N35730,N35731,N35732,N35733,N35734,N35735,N35736,N35737,N35738,
N35739,N35740,N35741,N35742,N35743,N35744,N35745,N35746,N35747,N35748,
N35749,N35750,N35751,N35752,N35753,N35754,N35755,N35756,N35757,N35758,
N35759,N35760,N35761,N35762,N35763,N35764,N35765,N35766,N35767,N35768,
N35769,N35770,N35771,N35772,N35773,N35774,N35775,N35776,N35777,N35778,
N35779,N35780,N35781,N35782,N35783,N35784,N35785,N35786,N35787,N35788,
N35789,N35790,N35791,N35792,N35793,N35794,N35795,N35796,N35797,N35798,
N35799,N35800,N35801,N35802,N35803,N35804,N35805,N35806,N35807,N35808,
N35809,N35810,N35811,N35812,N35813,N35814,N35815,N35816,N35817,N35818,
N35819,N35820,N35821,N35822,N35823,N35824,N35825,N35826,N35827,N35828,
N35829,N35830,N35831,N35832,N35833,N35834,N35835,N35836,N35837,N35838,
N35839,N35840,N35841,N35842,N35843,N35844,N35845,N35846,N35847,N35848,
N35849,N35850,N35851,N35852,N35853,N35854,N35855,N35856,N35857,N35858,
N35859,N35860,N35861,N35862,N35863,N35864,N35865,N35866,N35867,N35868,
N35869,N35870,N35871,N35872,N35873,N35874,N35875,N35876,N35877,N35878,
N35879,N35880,N35881,N35882,N35883,N35884,N35885,N35886,N35887,N35888,
N35889,N35890,N35891,N35892,N35893,N35894,N35895,N35896,N35897,N35898,
N35899,N35900,N35901,N35902,N35903,N35904,N35905,N35906,N35907,N35908,
N35909,N35910,N35911,N35912,N35913,N35914,N35915,N35916,N35917,N35918,
N35919,N35920,N35921,N35922,N35923,N35924,N35925,N35926,N35927,N35928,
N35929,N35930,N35931,N35932,N35933,N35934,N35935,N35936,N35937,N35938,
N35939,N35940,N35941,N35942,N35943,N35944,N35945,N35946,N35947,N35948,
N35949,N35950,N35951,N35952,N35953,N35954,N35955,N35956,N35957,N35958,
N35959,N35960,N35961,N35962,N35963,N35964,N35965,N35966,N35967,N35968,
N35969,N35970,N35971,N35972,N35973,N35974,N35975,N35976,N35977,N35978,
N35979,N35980,N35981,N35982,N35983,N35984,N35985,N35986,N35987,N35988,
N35989,N35990,N35991,N35992,N35993,N35994,N35995,N35996,N35997,N35998,
N35999,N36000,N36001,N36002,N36003,N36004,N36005,N36006,N36007,N36008,
N36009,N36010,N36011,N36012,N36013,N36014,N36015,N36016,N36017,N36018,
N36019,N36020,N36021,N36022,N36023,N36024,N36025,N36026,N36027,N36028,
N36029,N36030,N36031,N36032,N36033,N36034,N36035,N36036,N36037,N36038,
N36039,N36040,N36041,N36042,N36043,N36044,N36045,N36046,N36047,N36048,
N36049,N36050,N36051,N36052,N36053,N36054,N36055,N36056,N36057,N36058,
N36059,N36060,N36061,N36062,N36063,N36064,N36065,N36066,N36067,N36068,
N36069,N36070,N36071,N36072,N36073,N36074,N36075,N36076,N36077,N36078,
N36079,N36080,N36081,N36082,N36083,N36084,N36085,N36086,N36087,N36088,
N36089,N36090,N36091,N36092,N36093,N36094,N36095,N36096,N36097,N36098,
N36099,N36100,N36101,N36102,N36103,N36104,N36105,N36106,N36107,N36108,
N36109,N36110,N36111,N36112,N36113,N36114,N36115,N36116,N36117,N36118,
N36119,N36120,N36121,N36122,N36123,N36124,N36125,N36126,N36127,N36128,
N36129,N36130,N36131,N36132,N36133,N36134,N36135,N36136,N36137,N36138,
N36139,N36140,N36141,N36142,N36143,N36144,N36145,N36146,N36147,N36148,
N36149,N36150,N36151,N36152,N36153,N36154,N36155,N36156,N36157,N36158,
N36159,N36160,N36161,N36162,N36163,N36164,N36165,N36166,N36167,N36168,
N36169,N36170,N36171,N36172,N36173,N36174,N36175,N36176,N36177,N36178,
N36179,N36180,N36181,N36182,N36183,N36184,N36185,N36186,N36187,N36188,
N36189,N36190,N36191,N36192,N36193,N36194,N36195,N36196,N36197,N36198,
N36199,N36200,N36201,N36202,N36203,N36204,N36205,N36206,N36207,N36208,
N36209,N36210,N36211,N36212,N36213,N36214,N36215,N36216,N36217,N36218,
N36219,N36220,N36221,N36222,N36223,N36224,N36225,N36226,N36227,N36228,
N36229,N36230,N36231,N36232,N36233,N36234,N36235,N36236,N36237,N36238,
N36239,N36240,N36241,N36242,N36243,N36244,N36245,N36246,N36247,N36248,
N36249,N36250,N36251,N36252,N36253,N36254,N36255,N36256,N36257,N36258,
N36259,N36260,N36261,N36262,N36263,N36264,N36265,N36266,N36267,N36268,
N36269,N36270,N36271,N36272,N36273,N36274,N36275,N36276,N36277,N36278,
N36279,N36280,N36281,N36282,N36283,N36284,N36285,N36286,N36287,N36288,
N36289,N36290,N36291,N36292,N36293,N36294,N36295,N36296,N36297,N36298,
N36299,N36300,N36301,N36302,N36303,N36304,N36305,N36306,N36307,N36308,
N36309,N36310,N36311,N36312,N36313,N36314,N36315,N36316,N36317,N36318,
N36319,N36320,N36321,N36322,N36323,N36324,N36325,N36326,N36327,N36328,
N36329,N36330,N36331,N36332,N36333,N36334,N36335,N36336,N36337,N36338,
N36339,N36340,N36341,N36342,N36343,N36344,N36345,N36346,N36347,N36348,
N36349,N36350,N36351,N36352,N36353,N36354,N36355,N36356,N36357,N36358,
N36359,N36360,N36361,N36362,N36363,N36364,N36365,N36366,N36367,N36368,
N36369,N36370,N36371,N36372,N36373,N36374,N36375,N36376,N36377,N36378,
N36379,N36380,N36381,N36382,N36383,N36384,N36385,N36386,N36387,N36388,
N36389,N36390,N36391,N36392,N36393,N36394,N36395,N36396,N36397,N36398,
N36399,N36400,N36401,N36402,N36403,N36404,N36405,N36406,N36407,N36408,
N36409,N36410,N36411,N36412,N36413,N36414,N36415,N36416,N36417,N36418,
N36419,N36420,N36421,N36422,N36423,N36424,N36425,N36426,N36427,N36428,
N36429,N36430,N36431,N36432,N36433,N36434,N36435,N36436,N36437,N36438,
N36439,N36440,N36441,N36442,N36443,N36444,N36445,N36446,N36447,N36448,
N36449,N36450,N36451,N36452,N36453,N36454,N36455,N36456,N36457,N36458,
N36459,N36460,N36461,N36462,N36463,N36464,N36465,N36466,N36467,N36468,
N36469,N36470,N36471,N36472,N36473,N36474,N36475,N36476,N36477,N36478,
N36479,N36480,N36481,N36482,N36483,N36484,N36485,N36486,N36487,N36488,
N36489,N36490,N36491,N36492,N36493,N36494,N36495,N36496,N36497,N36498,
N36499,N36500,N36501,N36502,N36503,N36504,N36505,N36506,N36507,N36508,
N36509,N36510,N36511,N36512,N36513,N36514,N36515,N36516,N36517,N36518,
N36519,N36520,N36521,N36522,N36523,N36524,N36525,N36526,N36527,N36528,
N36529,N36530,N36531,N36532,N36533,N36534,N36535,N36536,N36537,N36538,
N36539,N36540,N36541,N36542,N36543,N36544,N36545,N36546,N36547,N36548,
N36549,N36550,N36551,N36552,N36553,N36554,N36555,N36556,N36557,N36558,
N36559,N36560,N36561,N36562,N36563,N36564,N36565,N36566,N36567,N36568,
N36569,N36570,N36571,N36572,N36573,N36574,N36575,N36576,N36577,N36578,
N36579,N36580,N36581,N36582,N36583,N36584,N36585,N36586,N36587,N36588,
N36589,N36590,N36591,N36592,N36593,N36594,N36595,N36596,N36597,N36598,
N36599,N36600,N36601,N36602,N36603,N36604,N36605,N36606,N36607,N36608,
N36609,N36610,N36611,N36612,N36613,N36614,N36615,N36616,N36617,N36618,
N36619,N36620,N36621,N36622,N36623,N36624,N36625,N36626,N36627,N36628,
N36629,N36630,N36631,N36632,N36633,N36634,N36635,N36636,N36637,N36638,
N36639,N36640,N36641,N36642,N36643,N36644,N36645,N36646,N36647,N36648,
N36649,N36650,N36651,N36652,N36653,N36654,N36655,N36656,N36657,N36658,
N36659,N36660,N36661,N36662,N36663,N36664,N36665,N36666,N36667,N36668,
N36669,N36670,N36671,N36672,N36673,N36674,N36675,N36676,N36677,N36678,
N36679,N36680,N36681,N36682,N36683,N36684,N36685,N36686,N36687,N36688,
N36689,N36690,N36691,N36692,N36693,N36694,N36695,N36696,N36697,N36698,
N36699,N36700,N36701,N36702,N36703,N36704,N36705,N36706,N36707,N36708,
N36709,N36710,N36711,N36712,N36713,N36714,N36715,N36716,N36717,N36718,
N36719,N36720,N36721,N36722,N36723,N36724,N36725,N36726,N36727,N36728,
N36729,N36730,N36731,N36732,N36733,N36734,N36735,N36736,N36737,N36738,
N36739,N36740,N36741,N36742,N36743,N36744,N36745,N36746,N36747,N36748,
N36749,N36750,N36751,N36752,N36753,N36754,N36755,N36756,N36757,N36758,
N36759,N36760,N36761,N36762,N36763,N36764,N36765,N36766,N36767,N36768,
N36769,N36770,N36771,N36772,N36773,N36774,N36775,N36776,N36777,N36778,
N36779,N36780,N36781,N36782,N36783,N36784,N36785,N36786,N36787,N36788,
N36789,N36790,N36791,N36792,N36793,N36794,N36795,N36796,N36797,N36798,
N36799,N36800,N36801,N36802,N36803,N36804,N36805,N36806,N36807,N36808,
N36809,N36810,N36811,N36812,N36813,N36814,N36815,N36816,N36817,N36818,
N36819,N36820,N36821,N36822,N36823,N36824,N36825,N36826,N36827,N36828,
N36829,N36830,N36831,N36832,N36833,N36834,N36835,N36836,N36837,N36838,
N36839,N36840,N36841,N36842,N36843,N36844,N36845,N36846,N36847,N36848,
N36849,N36850,N36851,N36852,N36853,N36854,N36855,N36856,N36857,N36858,
N36859,N36860,N36861,N36862,N36863,N36864,N36865,N36866,N36867,N36868,
N36869,N36870,N36871,N36872,N36873,N36874,N36875,N36876,N36877,N36878,
N36879,N36880,N36881,N36882,N36883,N36884,N36885,N36886,N36887,N36888,
N36889,N36890,N36891,N36892,N36893,N36894,N36895,N36896,N36897,N36898,
N36899,N36900,N36901,N36902,N36903,N36904,N36905,N36906,N36907,N36908,
N36909,N36910,N36911,N36912,N36913,N36914,N36915,N36916,N36917,N36918,
N36919,N36920,N36921,N36922,N36923,N36924,N36925,N36926,N36927,N36928,
N36929,N36930,N36931,N36932,N36933,N36934,N36935,N36936,N36937,N36938,
N36939,N36940,N36941,N36942,N36943,N36944,N36945,N36946,N36947,N36948,
N36949,N36950,N36951,N36952,N36953,N36954,N36955,N36956,N36957,N36958,
N36959,N36960,N36961,N36962,N36963,N36964,N36965,N36966,N36967,N36968,
N36969,N36970,N36971,N36972,N36973,N36974,N36975,N36976,N36977,N36978,
N36979,N36980,N36981,N36982,N36983,N36984,N36985,N36986,N36987,N36988,
N36989,N36990,N36991,N36992,N36993,N36994,N36995,N36996,N36997,N36998,
N36999,N37000,N37001,N37002,N37003,N37004,N37005,N37006,N37007,N37008,
N37009,N37010,N37011,N37012,N37013,N37014,N37015,N37016,N37017,N37018,
N37019,N37020,N37021,N37022,N37023,N37024,N37025,N37026,N37027,N37028,
N37029,N37030,N37031,N37032,N37033,N37034,N37035,N37036,N37037,N37038,
N37039,N37040,N37041,N37042,N37043,N37044,N37045,N37046,N37047,N37048,
N37049,N37050,N37051,N37052,N37053,N37054,N37055,N37056,N37057,N37058,
N37059,N37060,N37061,N37062,N37063,N37064,N37065,N37066,N37067,N37068,
N37069,N37070,N37071,N37072,N37073,N37074,N37075,N37076,N37077,N37078,
N37079,N37080,N37081,N37082,N37083,N37084,N37085,N37086,N37087,N37088,
N37089,N37090,N37091,N37092,N37093,N37094,N37095,N37096,N37097,N37098,
N37099,N37100,N37101,N37102,N37103,N37104,N37105,N37106,N37107,N37108,
N37109,N37110,N37111,N37112,N37113,N37114,N37115,N37116,N37117,N37118,
N37119,N37120,N37121,N37122,N37123,N37124,N37125,N37126,N37127,N37128,
N37129,N37130,N37131,N37132,N37133,N37134,N37135,N37136,N37137,N37138,
N37139,N37140,N37141,N37142,N37143,N37144,N37145,N37146,N37147,N37148,
N37149,N37150,N37151,N37152,N37153,N37154,N37155,N37156,N37157,N37158,
N37159,N37160,N37161,N37162,N37163,N37164,N37165,N37166,N37167,N37168,
N37169,N37170,N37171,N37172,N37173,N37174,N37175,N37176,N37177,N37178,
N37179,N37180,N37181,N37182,N37183,N37184,N37185,N37186,N37187,N37188,
N37189,N37190,N37191,N37192,N37193,N37194,N37195,N37196,N37197,N37198,
N37199,N37200,N37201,N37202,N37203,N37204,N37205,N37206,N37207,N37208,
N37209,N37210,N37211,N37212,N37213,N37214,N37215,N37216,N37217,N37218,
N37219,N37220,N37221,N37222,N37223,N37224,N37225,N37226,N37227,N37228,
N37229,N37230,N37231,N37232,N37233,N37234,N37235,N37236,N37237,N37238,
N37239,N37240,N37241,N37242,N37243,N37244,N37245,N37246,N37247,N37248,
N37249,N37250,N37251,N37252,N37253,N37254,N37255,N37256,N37257,N37258,
N37259,N37260,N37261,N37262,N37263,N37264,N37265,N37266,N37267,N37268,
N37269,N37270,N37271,N37272,N37273,N37274,N37275,N37276,N37277,N37278,
N37279,N37280,N37281,N37282,N37283,N37284,N37285,N37286,N37287,N37288,
N37289,N37290,N37291,N37292,N37293,N37294,N37295,N37296,N37297,N37298,
N37299,N37300,N37301,N37302,N37303,N37304,N37305,N37306,N37307,N37308,
N37309,N37310,N37311,N37312,N37313,N37314,N37315,N37316,N37317,N37318,
N37319,N37320,N37321,N37322,N37323,N37324,N37325,N37326,N37327,N37328,
N37329,N37330,N37331,N37332,N37333,N37334,N37335,N37336,N37337,N37338,
N37339,N37340,N37341,N37342,N37343,N37344,N37345,N37346,N37347,N37348,
N37349,N37350,N37351,N37352,N37353,N37354,N37355,N37356,N37357,N37358,
N37359,N37360,N37361,N37362,N37363,N37364,N37365,N37366,N37367,N37368,
N37369,N37370,N37371,N37372,N37373,N37374,N37375,N37376,N37377,N37378,
N37379,N37380,N37381,N37382,N37383,N37384,N37385,N37386,N37387,N37388,
N37389,N37390,N37391,N37392,N37393,N37394,N37395,N37396,N37397,N37398,
N37399,N37400,N37401,N37402,N37403,N37404,N37405,N37406,N37407,N37408,
N37409,N37410,N37411,N37412,N37413,N37414,N37415,N37416,N37417,N37418,
N37419,N37420,N37421,N37422,N37423,N37424,N37425,N37426,N37427,N37428,
N37429,N37430,N37431,N37432,N37433,N37434,N37435,N37436,N37437,N37438,
N37439,N37440,N37441,N37442,N37443,N37444,N37445,N37446,N37447,N37448,
N37449,N37450,N37451,N37452,N37453,N37454,N37455,N37456,N37457,N37458,
N37459,N37460,N37461,N37462,N37463,N37464,N37465,N37466,N37467,N37468,
N37469,N37470,N37471,N37472,N37473,N37474,N37475,N37476,N37477,N37478,
N37479,N37480,N37481,N37482,N37483,N37484,N37485,N37486,N37487,N37488,
N37489,N37490,N37491,N37492,N37493,N37494,N37495,N37496,N37497,N37498,
N37499,N37500,N37501,N37502,N37503,N37504,N37505,N37506,N37507,N37508,
N37509,N37510,N37511,N37512,N37513,N37514,N37515,N37516,N37517,N37518,
N37519,N37520,N37521,N37522,N37523,N37524,N37525,N37526,N37527,N37528,
N37529,N37530,N37531,N37532,N37533,N37534,N37535,N37536,N37537,N37538,
N37539,N37540,N37541,N37542,N37543,N37544,N37545,N37546,N37547,N37548,
N37549,N37550,N37551,N37552,N37553,N37554,N37555,N37556,N37557,N37558,
N37559,N37560,N37561,N37562,N37563,N37564,N37565,N37566,N37567,N37568,
N37569,N37570,N37571,N37572,N37573,N37574,N37575,N37576,N37577,N37578,
N37579,N37580,N37581,N37582,N37583,N37584,N37585,N37586,N37587,N37588,
N37589,N37590,N37591,N37592,N37593,N37594,N37595,N37596,N37597,N37598,
N37599,N37600,N37601,N37602,N37603,N37604,N37605,N37606,N37607,N37608,
N37609,N37610,N37611,N37612,N37613,N37614,N37615,N37616,N37617,N37618,
N37619,N37620,N37621,N37622,N37623,N37624,N37625,N37626,N37627,N37628,
N37629,N37630,N37631,N37632,N37633,N37634,N37635,N37636,N37637,N37638,
N37639,N37640,N37641,N37642,N37643,N37644,N37645,N37646,N37647,N37648,
N37649,N37650,N37651,N37652,N37653,N37654,N37655,N37656,N37657,N37658,
N37659,N37660,N37661,N37662,N37663,N37664,N37665,N37666,N37667,N37668,
N37669,N37670,N37671,N37672,N37673,N37674,N37675,N37676,N37677,N37678,
N37679,N37680,N37681,N37682,N37683,N37684,N37685,N37686,N37687,N37688,
N37689,N37690,N37691,N37692,N37693,N37694,N37695,N37696,N37697,N37698,
N37699,N37700,N37701,N37702,N37703,N37704,N37705,N37706,N37707,N37708,
N37709,N37710,N37711,N37712,N37713,N37714,N37715,N37716,N37717,N37718,
N37719,N37720,N37721,N37722,N37723,N37724,N37725,N37726,N37727,N37728,
N37729,N37730,N37731,N37732,N37733,N37734,N37735,N37736,N37737,N37738,
N37739,N37740,N37741,N37742,N37743,N37744,N37745,N37746,N37747,N37748,
N37749,N37750,N37751,N37752,N37753,N37754,N37755,N37756,N37757,N37758,
N37759,N37760,N37761,N37762,N37763,N37764,N37765,N37766,N37767,N37768,
N37769,N37770,N37771,N37772,N37773,N37774,N37775,N37776,N37777,N37778,
N37779,N37780,N37781,N37782,N37783,N37784,N37785,N37786,N37787,N37788,
N37789,N37790,N37791,N37792,N37793,N37794,N37795,N37796,N37797,N37798,
N37799,N37800,N37801,N37802,N37803,N37804,N37805,N37806,N37807,N37808,
N37809,N37810,N37811,N37812,N37813,N37814,N37815,N37816,N37817,N37818,
N37819,N37820,N37821,N37822,N37823,N37824,N37825,N37826,N37827,N37828,
N37829,N37830,N37831,N37832,N37833,N37834,N37835,N37836,N37837,N37838,
N37839,N37840,N37841,N37842,N37843,N37844,N37845,N37846,N37847,N37848,
N37849,N37850,N37851,N37852,N37853,N37854,N37855,N37856,N37857,N37858,
N37859,N37860,N37861,N37862,N37863,N37864,N37865,N37866,N37867,N37868,
N37869,N37870,N37871,N37872,N37873,N37874,N37875,N37876,N37877,N37878,
N37879,N37880,N37881,N37882,N37883,N37884,N37885,N37886,N37887,N37888,
N37889,N37890,N37891,N37892,N37893,N37894,N37895,N37896,N37897,N37898,
N37899,N37900,N37901,N37902,N37903,N37904,N37905,N37906,N37907,N37908,
N37909,N37910,N37911,N37912,N37913,N37914,N37915,N37916,N37917,N37918,
N37919,N37920,N37921,N37922,N37923,N37924,N37925,N37926,N37927,N37928,
N37929,N37930,N37931,N37932,N37933,N37934,N37935,N37936,N37937,N37938,
N37939,N37940,N37941,N37942,N37943,N37944,N37945,N37946,N37947,N37948,
N37949,N37950,N37951,N37952,N37953,N37954,N37955,N37956,N37957,N37958,
N37959,N37960,N37961,N37962,N37963,N37964,N37965,N37966,N37967,N37968,
N37969,N37970,N37971,N37972,N37973,N37974,N37975,N37976,N37977,N37978,
N37979,N37980,N37981,N37982,N37983,N37984,N37985,N37986,N37987,N37988,
N37989,N37990,N37991,N37992,N37993,N37994,N37995,N37996,N37997,N37998,
N37999,N38000,N38001,N38002,N38003,N38004,N38005,N38006,N38007,N38008,
N38009,N38010,N38011,N38012,N38013,N38014,N38015,N38016,N38017,N38018,
N38019,N38020,N38021,N38022,N38023,N38024,N38025,N38026,N38027,N38028,
N38029,N38030,N38031,N38032,N38033,N38034,N38035,N38036,N38037,N38038,
N38039,N38040,N38041,N38042,N38043,N38044,N38045,N38046,N38047,N38048,
N38049,N38050,N38051,N38052,N38053,N38054,N38055,N38056,N38057,N38058,
N38059,N38060,N38061,N38062,N38063,N38064,N38065,N38066,N38067,N38068,
N38069,N38070,N38071,N38072,N38073,N38074,N38075,N38076,N38077,N38078,
N38079,N38080,N38081,N38082,N38083,N38084,N38085,N38086,N38087,N38088,
N38089,N38090,N38091,N38092,N38093,N38094,N38095,N38096,N38097,N38098,
N38099,N38100,N38101,N38102,N38103,N38104,N38105,N38106,N38107,N38108,
N38109,N38110,N38111,N38112,N38113,N38114,N38115,N38116,N38117,N38118,
N38119,N38120,N38121,N38122,N38123,N38124,N38125,N38126,N38127,N38128,
N38129,N38130,N38131,N38132,N38133,N38134,N38135,N38136,N38137,N38138,
N38139,N38140,N38141,N38142,N38143,N38144,N38145,N38146,N38147,N38148,
N38149,N38150,N38151,N38152,N38153,N38154,N38155,N38156,N38157,N38158,
N38159,N38160,N38161,N38162,N38163,N38164,N38165,N38166,N38167,N38168,
N38169,N38170,N38171,N38172,N38173,N38174,N38175,N38176,N38177,N38178,
N38179,N38180,N38181,N38182,N38183,N38184,N38185,N38186,N38187,N38188,
N38189,N38190,N38191,N38192,N38193,N38194,N38195,N38196,N38197,N38198,
N38199,N38200,N38201,N38202,N38203,N38204,N38205,N38206,N38207,N38208,
N38209,N38210,N38211,N38212,N38213,N38214,N38215,N38216,N38217,N38218,
N38219,N38220,N38221,N38222,N38223,N38224,N38225,N38226,N38227,N38228,
N38229,N38230,N38231,N38232,N38233,N38234,N38235,N38236,N38237,N38238,
N38239,N38240,N38241,N38242,N38243,N38244,N38245,N38246,N38247,N38248,
N38249,N38250,N38251,N38252,N38253,N38254,N38255,N38256,N38257,N38258,
N38259,N38260,N38261,N38262,N38263,N38264,N38265,N38266,N38267,N38268,
N38269,N38270,N38271,N38272,N38273,N38274,N38275,N38276,N38277,N38278,
N38279,N38280,N38281,N38282,N38283,N38284,N38285,N38286,N38287,N38288,
N38289,N38290,N38291,N38292,N38293,N38294,N38295,N38296,N38297,N38298,
N38299,N38300,N38301,N38302,N38303,N38304,N38305,N38306,N38307,N38308,
N38309,N38310,N38311,N38312,N38313,N38314,N38315,N38316,N38317,N38318,
N38319,N38320,N38321,N38322,N38323,N38324,N38325,N38326,N38327,N38328,
N38329,N38330,N38331,N38332,N38333,N38334,N38335,N38336,N38337,N38338,
N38339,N38340,N38341,N38342,N38343,N38344,N38345,N38346,N38347,N38348,
N38349,N38350,N38351,N38352,N38353,N38354,N38355,N38356,N38357,N38358,
N38359,N38360,N38361,N38362,N38363,N38364,N38365,N38366,N38367,N38368,
N38369,N38370,N38371,N38372,N38373,N38374,N38375,N38376,N38377,N38378,
N38379,N38380,N38381,N38382,N38383,N38384,N38385,N38386,N38387,N38388,
N38389,N38390,N38391,N38392,N38393,N38394,N38395,N38396,N38397,N38398,
N38399,N38400,N38401,N38402,N38403,N38404,N38405,N38406,N38407,N38408,
N38409,N38410,N38411,N38412,N38413,N38414,N38415,N38416,N38417,N38418,
N38419,N38420,N38421,N38422,N38423,N38424,N38425,N38426,N38427,N38428,
N38429,N38430,N38431,N38432,N38433,N38434,N38435,N38436,N38437,N38438,
N38439,N38440,N38441,N38442,N38443,N38444,N38445,N38446,N38447,N38448,
N38449,N38450,N38451,N38452,N38453,N38454,N38455,N38456,N38457,N38458,
N38459,N38460,N38461,N38462,N38463,N38464,N38465,N38466,N38467,N38468,
N38469,N38470,N38471,N38472,N38473,N38474,N38475,N38476,N38477,N38478,
N38479,N38480,N38481,N38482,N38483,N38484,N38485,N38486,N38487,N38488,
N38489,N38490,N38491,N38492,N38493,N38494,N38495,N38496,N38497,N38498,
N38499,N38500,N38501,N38502,N38503,N38504,N38505,N38506,N38507,N38508,
N38509,N38510,N38511,N38512,N38513,N38514,N38515,N38516,N38517,N38518,
N38519,N38520,N38521,N38522,N38523,N38524,N38525,N38526,N38527,N38528,
N38529,N38530,N38531,N38532,N38533,N38534,N38535,N38536,N38537,N38538,
N38539,N38540,N38541,N38542,N38543,N38544,N38545,N38546,N38547,N38548,
N38549,N38550,N38551,N38552,N38553,N38554,N38555,N38556,N38557,N38558,
N38559,N38560,N38561,N38562,N38563,N38564,N38565,N38566,N38567,N38568,
N38569,N38570,N38571,N38572,N38573,N38574,N38575,N38576,N38577,N38578,
N38579,N38580,N38581,N38582,N38583,N38584,N38585,N38586,N38587,N38588,
N38589,N38590,N38591,N38592,N38593,N38594,N38595,N38596,N38597,N38598,
N38599,N38600,N38601,N38602,N38603,N38604,N38605,N38606,N38607,N38608,
N38609,N38610,N38611,N38612,N38613,N38614,N38615,N38616,N38617,N38618,
N38619,N38620,N38621,N38622,N38623,N38624,N38625,N38626,N38627,N38628,
N38629,N38630,N38631,N38632,N38633,N38634,N38635,N38636,N38637,N38638,
N38639,N38640,N38641,N38642,N38643,N38644,N38645,N38646,N38647,N38648,
N38649,N38650,N38651,N38652,N38653,N38654,N38655,N38656,N38657,N38658,
N38659,N38660,N38661,N38662,N38663,N38664,N38665,N38666,N38667,N38668,
N38669,N38670,N38671,N38672,N38673,N38674,N38675,N38676,N38677,N38678,
N38679,N38680,N38681,N38682,N38683,N38684,N38685,N38686,N38687,N38688,
N38689,N38690,N38691,N38692,N38693,N38694,N38695,N38696,N38697,N38698,
N38699,N38700,N38701,N38702,N38703,N38704,N38705,N38706,N38707,N38708,
N38709,N38710,N38711,N38712,N38713,N38714,N38715,N38716,N38717,N38718,
N38719,N38720,N38721,N38722,N38723,N38724,N38725,N38726,N38727,N38728,
N38729,N38730,N38731,N38732,N38733,N38734,N38735,N38736,N38737,N38738,
N38739,N38740,N38741,N38742,N38743,N38744,N38745,N38746,N38747,N38748,
N38749,N38750,N38751,N38752,N38753,N38754,N38755,N38756,N38757,N38758,
N38759,N38760,N38761,N38762,N38763,N38764,N38765,N38766,N38767,N38768,
N38769,N38770,N38771,N38772,N38773,N38774,N38775,N38776,N38777,N38778,
N38779,N38780,N38781,N38782,N38783,N38784,N38785,N38786,N38787,N38788,
N38789,N38790,N38791,N38792,N38793,N38794,N38795,N38796,N38797,N38798,
N38799,N38800,N38801,N38802,N38803,N38804,N38805,N38806,N38807,N38808,
N38809,N38810,N38811,N38812,N38813,N38814,N38815,N38816,N38817,N38818,
N38819,N38820,N38821,N38822,N38823,N38824,N38825,N38826,N38827,N38828,
N38829,N38830,N38831,N38832,N38833,N38834,N38835,N38836,N38837,N38838,
N38839,N38840,N38841,N38842,N38843,N38844,N38845,N38846,N38847,N38848,
N38849,N38850,N38851,N38852,N38853,N38854,N38855,N38856,N38857,N38858,
N38859,N38860,N38861,N38862,N38863,N38864,N38865,N38866,N38867,N38868,
N38869,N38870,N38871,N38872,N38873,N38874,N38875,N38876,N38877,N38878,
N38879,N38880,N38881,N38882,N38883,N38884,N38885,N38886,N38887,N38888,
N38889,N38890,N38891,N38892,N38893,N38894,N38895,N38896,N38897,N38898,
N38899,N38900,N38901,N38902,N38903,N38904,N38905,N38906,N38907,N38908,
N38909,N38910,N38911,N38912,N38913,N38914,N38915,N38916,N38917,N38918,
N38919,N38920,N38921,N38922,N38923,N38924,N38925,N38926,N38927,N38928,
N38929,N38930,N38931,N38932,N38933,N38934,N38935,N38936,N38937,N38938,
N38939,N38940,N38941,N38942,N38943,N38944,N38945,N38946,N38947,N38948,
N38949,N38950,N38951,N38952,N38953,N38954,N38955,N38956,N38957,N38958,
N38959,N38960,N38961,N38962,N38963,N38964,N38965,N38966,N38967,N38968,
N38969,N38970,N38971,N38972,N38973,N38974,N38975,N38976,N38977,N38978,
N38979,N38980,N38981,N38982,N38983,N38984,N38985,N38986,N38987,N38988,
N38989,N38990,N38991,N38992,N38993,N38994,N38995,N38996,N38997,N38998,
N38999,N39000,N39001,N39002,N39003,N39004,N39005,N39006,N39007,N39008,
N39009,N39010,N39011,N39012,N39013,N39014,N39015,N39016,N39017,N39018,
N39019,N39020,N39021,N39022,N39023,N39024,N39025,N39026,N39027,N39028,
N39029,N39030,N39031,N39032,N39033,N39034,N39035,N39036,N39037,N39038,
N39039,N39040,N39041,N39042,N39043,N39044,N39045,N39046,N39047,N39048,
N39049,N39050,N39051,N39052,N39053,N39054,N39055,N39056,N39057,N39058,
N39059,N39060,N39061,N39062,N39063,N39064,N39065,N39066,N39067,N39068,
N39069,N39070,N39071,N39072,N39073,N39074,N39075,N39076,N39077,N39078,
N39079,N39080,N39081,N39082,N39083,N39084,N39085,N39086,N39087,N39088,
N39089,N39090,N39091,N39092,N39093,N39094,N39095,N39096,N39097,N39098,
N39099,N39100,N39101,N39102,N39103,N39104,N39105,N39106,N39107,N39108,
N39109,N39110,N39111,N39112,N39113,N39114,N39115,N39116,N39117,N39118,
N39119,N39120,N39121,N39122,N39123,N39124,N39125,N39126,N39127,N39128,
N39129,N39130,N39131,N39132,N39133,N39134,N39135,N39136,N39137,N39138,
N39139,N39140,N39141,N39142,N39143,N39144,N39145,N39146,N39147,N39148,
N39149,N39150,N39151,N39152,N39153,N39154,N39155,N39156,N39157,N39158,
N39159,N39160,N39161,N39162,N39163,N39164,N39165,N39166,N39167,N39168,
N39169,N39170,N39171,N39172,N39173,N39174,N39175,N39176,N39177,N39178,
N39179,N39180,N39181,N39182,N39183,N39184,N39185,N39186,N39187,N39188,
N39189,N39190,N39191,N39192,N39193,N39194,N39195,N39196,N39197,N39198,
N39199,N39200,N39201,N39202,N39203,N39204,N39205,N39206,N39207,N39208,
N39209,N39210,N39211,N39212,N39213,N39214,N39215,N39216,N39217,N39218,
N39219,N39220,N39221,N39222,N39223,N39224,N39225,N39226,N39227,N39228,
N39229,N39230,N39231,N39232,N39233,N39234,N39235,N39236,N39237,N39238,
N39239,N39240,N39241,N39242,N39243,N39244,N39245,N39246,N39247,N39248,
N39249,N39250,N39251,N39252,N39253,N39254,N39255,N39256,N39257,N39258,
N39259,N39260,N39261,N39262,N39263,N39264,N39265,N39266,N39267,N39268,
N39269,N39270,N39271,N39272,N39273,N39274,N39275,N39276,N39277,N39278,
N39279,N39280,N39281,N39282,N39283,N39284,N39285,N39286,N39287,N39288,
N39289,N39290,N39291,N39292,N39293,N39294,N39295,N39296,N39297,N39298,
N39299,N39300,N39301,N39302,N39303,N39304,N39305,N39306,N39307,N39308,
N39309,N39310,N39311,N39312,N39313,N39314,N39315,N39316,N39317,N39318,
N39319,N39320,N39321,N39322,N39323,N39324,N39325,N39326,N39327,N39328,
N39329,N39330,N39331,N39332,N39333,N39334,N39335,N39336,N39337,N39338,
N39339,N39340,N39341,N39342,N39343,N39344,N39345,N39346,N39347,N39348,
N39349,N39350,N39351,N39352,N39353,N39354,N39355,N39356,N39357,N39358,
N39359,N39360,N39361,N39362,N39363,N39364,N39365,N39366,N39367,N39368,
N39369,N39370,N39371,N39372,N39373,N39374,N39375,N39376,N39377,N39378,
N39379,N39380,N39381,N39382,N39383,N39384,N39385,N39386,N39387,N39388,
N39389,N39390,N39391,N39392,N39393,N39394,N39395,N39396,N39397,N39398,
N39399,N39400,N39401,N39402,N39403,N39404,N39405,N39406,N39407,N39408,
N39409,N39410,N39411,N39412,N39413,N39414,N39415,N39416,N39417,N39418,
N39419,N39420,N39421,N39422,N39423,N39424,N39425,N39426,N39427,N39428,
N39429,N39430,N39431,N39432,N39433,N39434,N39435,N39436,N39437,N39438,
N39439,N39440,N39441,N39442,N39443,N39444,N39445,N39446,N39447,N39448,
N39449,N39450,N39451,N39452,N39453,N39454,N39455,N39456,N39457,N39458,
N39459,N39460,N39461,N39462,N39463,N39464,N39465,N39466,N39467,N39468,
N39469,N39470,N39471,N39472,N39473,N39474,N39475,N39476,N39477,N39478,
N39479,N39480,N39481,N39482,N39483,N39484,N39485,N39486,N39487,N39488,
N39489,N39490,N39491,N39492,N39493,N39494,N39495,N39496,N39497,N39498,
N39499,N39500,N39501,N39502,N39503,N39504,N39505,N39506,N39507,N39508,
N39509,N39510,N39511,N39512,N39513,N39514,N39515,N39516,N39517,N39518,
N39519,N39520,N39521,N39522,N39523,N39524,N39525,clk,rst;

reg R0,R1,R2,R3,R4,R5,R6,R7,O0,O1,O2,O3,O4,O5;

always@(posedge clk or negedge rst)
 if(!rst)
   R0 <= N0;
   else
   R0= 1'b0;

always@(posedge clk or negedge rst)
 if(!rst)
   R1 <= N5497;
   else
   R1= 1'b0;

always@(posedge clk or negedge rst)
 if(!rst)
   R2 <= N11430;
   else
   R2= 1'b0;

always@(posedge clk or negedge rst)
 if(!rst)
   R3 <= N17644;
   else
   R3= 1'b0;

always@(posedge clk or negedge rst)
 if(!rst)
   R4 <= N24056;
   else
   R4= 1'b0;

always@(posedge clk or negedge rst)
 if(!rst)
   R5 <= N29273;
   else
   R5= 1'b0;

always@(posedge clk or negedge rst)
 if(!rst)
   R6 <= N31740;
   else
   R6= 1'b0;

always@(posedge clk or negedge rst)
 if(!rst)
   R7 <= N34392;
   else
   R7= 1'b0;

always@(posedge clk or negedge rst)
  if(!rst)
   O0 <= N37264;
  else
       O0=1'b0;
always@(posedge clk or negedge rst)
  if(!rst)
   O1 <= N37882;
  else
       O1=1'b0;
always@(posedge clk or negedge rst)
  if(!rst)
   O2 <= N38213;
  else
       O2=1'b0;
always@(posedge clk or negedge rst)
  if(!rst)
   O3 <= N38364;
  else
       O3=1'b0;
always@(posedge clk or negedge rst)
  if(!rst)
   O4 <= N38772;
  else
       O4=1'b0;
always@(posedge clk or negedge rst)
  if(!rst)
   O5 <= N39035;
  else
       O5=1'b0;

and and0(N388,N389,N390);
and and9(N405,N406,N407);
and and18(N422,N423,N424);
and and27(N439,N440,N441);
and and36(N456,N457,N458);
and and45(N473,N474,N475);
and and54(N489,N490,N491);
and and63(N505,N506,N507);
and and72(N521,N522,N523);
and and81(N537,N538,N539);
and and90(N553,N554,N555);
and and99(N569,N570,N571);
and and108(N585,N586,N587);
and and117(N601,N602,N603);
and and126(N617,N618,N619);
and and135(N633,N634,N635);
and and144(N649,N650,N651);
and and153(N665,N666,N667);
and and162(N681,N682,N683);
and and171(N697,N698,N699);
and and180(N713,N714,N715);
and and189(N729,N730,N731);
and and198(N745,N746,N747);
and and207(N761,N762,N763);
and and216(N777,N778,N779);
and and225(N793,N794,N795);
and and234(N809,N810,N811);
and and243(N824,N825,N826);
and and252(N839,N840,N841);
and and261(N854,N855,N856);
and and270(N869,N870,N871);
and and279(N884,N885,N886);
and and288(N899,N900,N901);
and and297(N914,N915,N916);
and and306(N929,N930,N931);
and and315(N944,N945,N946);
and and324(N959,N960,N961);
and and333(N974,N975,N976);
and and342(N989,N990,N991);
and and351(N1004,N1005,N1006);
and and360(N1019,N1020,N1021);
and and369(N1034,N1035,N1036);
and and378(N1049,N1050,N1051);
and and387(N1064,N1065,N1066);
and and396(N1079,N1080,N1081);
and and405(N1094,N1095,N1096);
and and414(N1109,N1110,N1111);
and and423(N1124,N1125,N1126);
and and432(N1139,N1140,N1141);
and and441(N1154,N1155,N1156);
and and450(N1169,N1170,N1171);
and and459(N1184,N1185,N1186);
and and468(N1199,N1200,N1201);
and and477(N1214,N1215,N1216);
and and486(N1229,N1230,N1231);
and and495(N1244,N1245,N1246);
and and504(N1259,N1260,N1261);
and and513(N1274,N1275,N1276);
and and522(N1289,N1290,N1291);
and and531(N1304,N1305,N1306);
and and540(N1319,N1320,N1321);
and and549(N1334,N1335,N1336);
and and558(N1349,N1350,N1351);
and and567(N1364,N1365,N1366);
and and576(N1379,N1380,N1381);
and and585(N1394,N1395,N1396);
and and594(N1409,N1410,N1411);
and and603(N1424,N1425,N1426);
and and612(N1438,N1439,N1440);
and and621(N1452,N1453,N1454);
and and630(N1466,N1467,N1468);
and and639(N1480,N1481,N1482);
and and648(N1494,N1495,N1496);
and and657(N1508,N1509,N1510);
and and666(N1522,N1523,N1524);
and and675(N1536,N1537,N1538);
and and684(N1550,N1551,N1552);
and and693(N1564,N1565,N1566);
and and702(N1578,N1579,N1580);
and and711(N1592,N1593,N1594);
and and720(N1606,N1607,N1608);
and and729(N1620,N1621,N1622);
and and738(N1634,N1635,N1636);
and and747(N1648,N1649,N1650);
and and756(N1662,N1663,N1664);
and and765(N1676,N1677,N1678);
and and774(N1690,N1691,N1692);
and and783(N1704,N1705,N1706);
and and792(N1718,N1719,N1720);
and and801(N1732,N1733,N1734);
and and810(N1746,N1747,N1748);
and and819(N1760,N1761,N1762);
and and828(N1774,N1775,N1776);
and and837(N1788,N1789,N1790);
and and846(N1802,N1803,N1804);
and and855(N1816,N1817,N1818);
and and864(N1830,N1831,N1832);
and and873(N1844,N1845,N1846);
and and882(N1858,N1859,N1860);
and and891(N1872,N1873,N1874);
and and900(N1886,N1887,N1888);
and and909(N1900,N1901,N1902);
and and918(N1914,N1915,N1916);
and and927(N1928,N1929,N1930);
and and936(N1942,N1943,N1944);
and and945(N1956,N1957,N1958);
and and954(N1970,N1971,N1972);
and and963(N1984,N1985,N1986);
and and972(N1998,N1999,N2000);
and and981(N2012,N2013,N2014);
and and990(N2026,N2027,N2028);
and and999(N2040,N2041,N2042);
and and1008(N2054,N2055,N2056);
and and1017(N2068,N2069,N2070);
and and1026(N2082,N2083,N2084);
and and1035(N2096,N2097,N2098);
and and1044(N2110,N2111,N2112);
and and1053(N2123,N2124,N2125);
and and1062(N2136,N2137,N2138);
and and1071(N2149,N2150,N2151);
and and1080(N2162,N2163,N2164);
and and1089(N2175,N2176,N2177);
and and1098(N2188,N2189,N2190);
and and1107(N2201,N2202,N2203);
and and1116(N2214,N2215,N2216);
and and1125(N2227,N2228,N2229);
and and1134(N2240,N2241,N2242);
and and1143(N2253,N2254,N2255);
and and1152(N2266,N2267,N2268);
and and1161(N2279,N2280,N2281);
and and1170(N2292,N2293,N2294);
and and1179(N2305,N2306,N2307);
and and1188(N2318,N2319,N2320);
and and1197(N2331,N2332,N2333);
and and1206(N2344,N2345,N2346);
and and1215(N2357,N2358,N2359);
and and1224(N2370,N2371,N2372);
and and1233(N2383,N2384,N2385);
and and1242(N2396,N2397,N2398);
and and1251(N2409,N2410,N2411);
and and1260(N2422,N2423,N2424);
and and1269(N2435,N2436,N2437);
and and1278(N2448,N2449,N2450);
and and1287(N2461,N2462,N2463);
and and1296(N2474,N2475,N2476);
and and1305(N2487,N2488,N2489);
and and1314(N2500,N2501,N2502);
and and1323(N2513,N2514,N2515);
and and1332(N2526,N2527,N2528);
and and1341(N2539,N2540,N2541);
and and1350(N2552,N2553,N2554);
and and1359(N2565,N2566,N2567);
and and1368(N2578,N2579,N2580);
and and1377(N2591,N2592,N2593);
and and1386(N2604,N2605,N2606);
and and1395(N2616,N2617,N2618);
and and1404(N2628,N2629,N2630);
and and1413(N2640,N2641,N2642);
and and1422(N2652,N2653,N2654);
and and1431(N2664,N2665,N2666);
and and1440(N2676,N2677,N2678);
and and1449(N2688,N2689,N2690);
and and1458(N2700,N2701,N2702);
and and1467(N2712,N2713,N2714);
and and1476(N2724,N2725,N2726);
and and1485(N2736,N2737,N2738);
and and1494(N2748,N2749,N2750);
and and1503(N2760,N2761,N2762);
and and1512(N2772,N2773,N2774);
and and1521(N2784,N2785,N2786);
and and1530(N2796,N2797,N2798);
and and1539(N2808,N2809,N2810);
and and1548(N2820,N2821,N2822);
and and1557(N2832,N2833,N2834);
and and1566(N2844,N2845,N2846);
and and1575(N2856,N2857,N2858);
and and1584(N2868,N2869,N2870);
and and1593(N2880,N2881,N2882);
and and1602(N2892,N2893,N2894);
and and1611(N2904,N2905,N2906);
and and1620(N2916,N2917,N2918);
and and1629(N2928,N2929,N2930);
and and1638(N2940,N2941,N2942);
and and1647(N2952,N2953,N2954);
and and1656(N2964,N2965,N2966);
and and1665(N2976,N2977,N2978);
and and1674(N2988,N2989,N2990);
and and1683(N3000,N3001,N3002);
and and1692(N3012,N3013,N3014);
and and1701(N3024,N3025,N3026);
and and1710(N3036,N3037,N3038);
and and1719(N3048,N3049,N3050);
and and1728(N3060,N3061,N3062);
and and1737(N3072,N3073,N3074);
and and1746(N3084,N3085,N3086);
and and1755(N3095,N3096,N3097);
and and1764(N3106,N3107,N3108);
and and1773(N3117,N3118,N3119);
and and1782(N3128,N3129,N3130);
and and1791(N3139,N3140,N3141);
and and1800(N3150,N3151,N3152);
and and1809(N3161,N3162,N3163);
and and1818(N3172,N3173,N3174);
and and1827(N3183,N3184,N3185);
and and1836(N3194,N3195,N3196);
and and1845(N3205,N3206,N3207);
and and1854(N3216,N3217,N3218);
and and1863(N3227,N3228,N3229);
and and1872(N3237,N3238,N3239);
and and1881(N3247,N3248,N3249);
and and1890(N3256,N3257,N3258);
and and1898(N3272,N3273,N3274);
and and1906(N3288,N3289,N3290);
and and1914(N3304,N3305,N3306);
and and1922(N3320,N3321,N3322);
and and1930(N3336,N3337,N3338);
and and1938(N3352,N3353,N3354);
and and1946(N3368,N3369,N3370);
and and1954(N3383,N3384,N3385);
and and1962(N3398,N3399,N3400);
and and1970(N3413,N3414,N3415);
and and1978(N3428,N3429,N3430);
and and1986(N3443,N3444,N3445);
and and1994(N3458,N3459,N3460);
and and2002(N3473,N3474,N3475);
and and2010(N3488,N3489,N3490);
and and2018(N3503,N3504,N3505);
and and2026(N3518,N3519,N3520);
and and2034(N3532,N3533,N3534);
and and2042(N3546,N3547,N3548);
and and2050(N3560,N3561,N3562);
and and2058(N3574,N3575,N3576);
and and2066(N3588,N3589,N3590);
and and2074(N3602,N3603,N3604);
and and2082(N3616,N3617,N3618);
and and2090(N3630,N3631,N3632);
and and2098(N3644,N3645,N3646);
and and2106(N3658,N3659,N3660);
and and2114(N3672,N3673,N3674);
and and2122(N3686,N3687,N3688);
and and2130(N3700,N3701,N3702);
and and2138(N3714,N3715,N3716);
and and2146(N3728,N3729,N3730);
and and2154(N3742,N3743,N3744);
and and2162(N3756,N3757,N3758);
and and2170(N3770,N3771,N3772);
and and2178(N3784,N3785,N3786);
and and2186(N3798,N3799,N3800);
and and2194(N3812,N3813,N3814);
and and2202(N3826,N3827,N3828);
and and2210(N3840,N3841,N3842);
and and2218(N3854,N3855,N3856);
and and2226(N3868,N3869,N3870);
and and2234(N3882,N3883,N3884);
and and2242(N3895,N3896,N3897);
and and2250(N3908,N3909,N3910);
and and2258(N3921,N3922,N3923);
and and2266(N3934,N3935,N3936);
and and2274(N3947,N3948,N3949);
and and2282(N3960,N3961,N3962);
and and2290(N3973,N3974,N3975);
and and2298(N3986,N3987,N3988);
and and2306(N3999,N4000,N4001);
and and2314(N4012,N4013,N4014);
and and2322(N4025,N4026,N4027);
and and2330(N4038,N4039,N4040);
and and2338(N4051,N4052,N4053);
and and2346(N4064,N4065,N4066);
and and2354(N4077,N4078,N4079);
and and2362(N4090,N4091,N4092);
and and2370(N4103,N4104,N4105);
and and2378(N4116,N4117,N4118);
and and2386(N4129,N4130,N4131);
and and2394(N4142,N4143,N4144);
and and2402(N4155,N4156,N4157);
and and2410(N4168,N4169,N4170);
and and2418(N4181,N4182,N4183);
and and2426(N4194,N4195,N4196);
and and2434(N4207,N4208,N4209);
and and2442(N4220,N4221,N4222);
and and2450(N4233,N4234,N4235);
and and2458(N4246,N4247,N4248);
and and2466(N4259,N4260,N4261);
and and2474(N4272,N4273,N4274);
and and2482(N4285,N4286,N4287);
and and2490(N4298,N4299,N4300);
and and2498(N4311,N4312,N4313);
and and2506(N4324,N4325,N4326);
and and2514(N4337,N4338,N4339);
and and2522(N4350,N4351,N4352);
and and2530(N4363,N4364,N4365);
and and2538(N4376,N4377,N4378);
and and2546(N4389,N4390,N4391);
and and2554(N4402,N4403,N4404);
and and2562(N4415,N4416,N4417);
and and2570(N4428,N4429,N4430);
and and2578(N4441,N4442,N4443);
and and2586(N4454,N4455,N4456);
and and2594(N4467,N4468,N4469);
and and2602(N4480,N4481,N4482);
and and2610(N4493,N4494,N4495);
and and2618(N4505,N4506,N4507);
and and2626(N4517,N4518,N4519);
and and2634(N4529,N4530,N4531);
and and2642(N4541,N4542,N4543);
and and2650(N4553,N4554,N4555);
and and2658(N4565,N4566,N4567);
and and2666(N4577,N4578,N4579);
and and2674(N4589,N4590,N4591);
and and2682(N4601,N4602,N4603);
and and2690(N4613,N4614,N4615);
and and2698(N4625,N4626,N4627);
and and2706(N4637,N4638,N4639);
and and2714(N4649,N4650,N4651);
and and2722(N4661,N4662,N4663);
and and2730(N4673,N4674,N4675);
and and2738(N4685,N4686,N4687);
and and2746(N4697,N4698,N4699);
and and2754(N4709,N4710,N4711);
and and2762(N4721,N4722,N4723);
and and2770(N4733,N4734,N4735);
and and2778(N4745,N4746,N4747);
and and2786(N4757,N4758,N4759);
and and2794(N4769,N4770,N4771);
and and2802(N4781,N4782,N4783);
and and2810(N4793,N4794,N4795);
and and2818(N4805,N4806,N4807);
and and2826(N4817,N4818,N4819);
and and2834(N4829,N4830,N4831);
and and2842(N4841,N4842,N4843);
and and2850(N4853,N4854,N4855);
and and2858(N4865,N4866,N4867);
and and2866(N4877,N4878,N4879);
and and2874(N4889,N4890,N4891);
and and2882(N4901,N4902,N4903);
and and2890(N4913,N4914,N4915);
and and2898(N4925,N4926,N4927);
and and2906(N4937,N4938,N4939);
and and2914(N4949,N4950,N4951);
and and2922(N4961,N4962,N4963);
and and2930(N4973,N4974,N4975);
and and2938(N4984,N4985,N4986);
and and2946(N4995,N4996,N4997);
and and2954(N5006,N5007,N5008);
and and2962(N5017,N5018,N5019);
and and2970(N5028,N5029,N5030);
and and2978(N5039,N5040,N5041);
and and2986(N5050,N5051,N5052);
and and2994(N5061,N5062,N5063);
and and3002(N5072,N5073,N5074);
and and3010(N5083,N5084,N5085);
and and3018(N5094,N5095,N5096);
and and3026(N5105,N5106,N5107);
and and3034(N5116,N5117,N5118);
and and3042(N5127,N5128,N5129);
and and3050(N5138,N5139,N5140);
and and3058(N5149,N5150,N5151);
and and3066(N5160,N5161,N5162);
and and3074(N5171,N5172,N5173);
and and3082(N5182,N5183,N5184);
and and3090(N5192,N5193,N5194);
and and3098(N5202,N5203,N5204);
and and3106(N5212,N5213,N5214);
and and3114(N5222,N5223,N5224);
and and3122(N5232,N5233,N5234);
and and3130(N5242,N5243,N5244);
and and3138(N5252,N5253,N5254);
and and3146(N5261,N5262,N5263);
and and3154(N5270,N5271,N5272);
and and3162(N5279,N5280,N5281);
and and3169(N5293,N5294,N5295);
and and3176(N5306,N5307,N5308);
and and3183(N5319,N5320,N5321);
and and3190(N5331,N5332,N5333);
and and3197(N5343,N5344,N5345);
and and3204(N5355,N5356,N5357);
and and3211(N5367,N5368,N5369);
and and3218(N5378,N5379,N5380);
and and3225(N5389,N5390,N5391);
and and3232(N5400,N5401,N5402);
and and3239(N5411,N5412,N5413);
and and3246(N5422,N5423,N5424);
and and3253(N5432,N5433,N5434);
and and3260(N5442,N5443,N5444);
and and3267(N5452,N5453,N5454);
and and3274(N5462,N5463,N5464);
and and3281(N5471,N5472,N5473);
and and3288(N5480,N5481,N5482);
and and3295(N5489,N5490,N5491);
and and1(N389,N391,N392);
and and2(N390,N393,N394);
and and10(N406,N408,N409);
and and11(N407,N410,N411);
and and19(N423,N425,N426);
and and20(N424,N427,N428);
and and28(N440,N442,N443);
and and29(N441,N444,N445);
and and37(N457,N459,N460);
and and38(N458,N461,N462);
and and46(N474,N476,N477);
and and47(N475,N478,N479);
and and55(N490,N492,N493);
and and56(N491,N494,N495);
and and64(N506,N508,N509);
and and65(N507,N510,N511);
and and73(N522,N524,N525);
and and74(N523,N526,N527);
and and82(N538,N540,N541);
and and83(N539,N542,N543);
and and91(N554,N556,N557);
and and92(N555,N558,N559);
and and100(N570,N572,N573);
and and101(N571,N574,N575);
and and109(N586,N588,N589);
and and110(N587,N590,N591);
and and118(N602,N604,N605);
and and119(N603,N606,N607);
and and127(N618,N620,N621);
and and128(N619,N622,N623);
and and136(N634,N636,N637);
and and137(N635,N638,N639);
and and145(N650,N652,N653);
and and146(N651,N654,N655);
and and154(N666,N668,N669);
and and155(N667,N670,N671);
and and163(N682,N684,N685);
and and164(N683,N686,N687);
and and172(N698,N700,N701);
and and173(N699,N702,N703);
and and181(N714,N716,N717);
and and182(N715,N718,N719);
and and190(N730,N732,N733);
and and191(N731,N734,N735);
and and199(N746,N748,N749);
and and200(N747,N750,N751);
and and208(N762,N764,N765);
and and209(N763,N766,N767);
and and217(N778,N780,N781);
and and218(N779,N782,N783);
and and226(N794,N796,N797);
and and227(N795,N798,N799);
and and235(N810,N812,N813);
and and236(N811,N814,N815);
and and244(N825,N827,N828);
and and245(N826,N829,N830);
and and253(N840,N842,N843);
and and254(N841,N844,N845);
and and262(N855,N857,N858);
and and263(N856,N859,N860);
and and271(N870,N872,N873);
and and272(N871,N874,N875);
and and280(N885,N887,N888);
and and281(N886,N889,N890);
and and289(N900,N902,N903);
and and290(N901,N904,N905);
and and298(N915,N917,N918);
and and299(N916,N919,N920);
and and307(N930,N932,N933);
and and308(N931,N934,N935);
and and316(N945,N947,N948);
and and317(N946,N949,N950);
and and325(N960,N962,N963);
and and326(N961,N964,N965);
and and334(N975,N977,N978);
and and335(N976,N979,N980);
and and343(N990,N992,N993);
and and344(N991,N994,N995);
and and352(N1005,N1007,N1008);
and and353(N1006,N1009,N1010);
and and361(N1020,N1022,N1023);
and and362(N1021,N1024,N1025);
and and370(N1035,N1037,N1038);
and and371(N1036,N1039,N1040);
and and379(N1050,N1052,N1053);
and and380(N1051,N1054,N1055);
and and388(N1065,N1067,N1068);
and and389(N1066,N1069,N1070);
and and397(N1080,N1082,N1083);
and and398(N1081,N1084,N1085);
and and406(N1095,N1097,N1098);
and and407(N1096,N1099,N1100);
and and415(N1110,N1112,N1113);
and and416(N1111,N1114,N1115);
and and424(N1125,N1127,N1128);
and and425(N1126,N1129,N1130);
and and433(N1140,N1142,N1143);
and and434(N1141,N1144,N1145);
and and442(N1155,N1157,N1158);
and and443(N1156,N1159,N1160);
and and451(N1170,N1172,N1173);
and and452(N1171,N1174,N1175);
and and460(N1185,N1187,N1188);
and and461(N1186,N1189,N1190);
and and469(N1200,N1202,N1203);
and and470(N1201,N1204,N1205);
and and478(N1215,N1217,N1218);
and and479(N1216,N1219,N1220);
and and487(N1230,N1232,N1233);
and and488(N1231,N1234,N1235);
and and496(N1245,N1247,N1248);
and and497(N1246,N1249,N1250);
and and505(N1260,N1262,N1263);
and and506(N1261,N1264,N1265);
and and514(N1275,N1277,N1278);
and and515(N1276,N1279,N1280);
and and523(N1290,N1292,N1293);
and and524(N1291,N1294,N1295);
and and532(N1305,N1307,N1308);
and and533(N1306,N1309,N1310);
and and541(N1320,N1322,N1323);
and and542(N1321,N1324,N1325);
and and550(N1335,N1337,N1338);
and and551(N1336,N1339,N1340);
and and559(N1350,N1352,N1353);
and and560(N1351,N1354,N1355);
and and568(N1365,N1367,N1368);
and and569(N1366,N1369,N1370);
and and577(N1380,N1382,N1383);
and and578(N1381,N1384,N1385);
and and586(N1395,N1397,N1398);
and and587(N1396,N1399,N1400);
and and595(N1410,N1412,N1413);
and and596(N1411,N1414,N1415);
and and604(N1425,N1427,N1428);
and and605(N1426,N1429,N1430);
and and613(N1439,N1441,N1442);
and and614(N1440,N1443,N1444);
and and622(N1453,N1455,N1456);
and and623(N1454,N1457,N1458);
and and631(N1467,N1469,N1470);
and and632(N1468,N1471,N1472);
and and640(N1481,N1483,N1484);
and and641(N1482,N1485,N1486);
and and649(N1495,N1497,N1498);
and and650(N1496,N1499,N1500);
and and658(N1509,N1511,N1512);
and and659(N1510,N1513,N1514);
and and667(N1523,N1525,N1526);
and and668(N1524,N1527,N1528);
and and676(N1537,N1539,N1540);
and and677(N1538,N1541,N1542);
and and685(N1551,N1553,N1554);
and and686(N1552,N1555,N1556);
and and694(N1565,N1567,N1568);
and and695(N1566,N1569,N1570);
and and703(N1579,N1581,N1582);
and and704(N1580,N1583,N1584);
and and712(N1593,N1595,N1596);
and and713(N1594,N1597,N1598);
and and721(N1607,N1609,N1610);
and and722(N1608,N1611,N1612);
and and730(N1621,N1623,N1624);
and and731(N1622,N1625,N1626);
and and739(N1635,N1637,N1638);
and and740(N1636,N1639,N1640);
and and748(N1649,N1651,N1652);
and and749(N1650,N1653,N1654);
and and757(N1663,N1665,N1666);
and and758(N1664,N1667,N1668);
and and766(N1677,N1679,N1680);
and and767(N1678,N1681,N1682);
and and775(N1691,N1693,N1694);
and and776(N1692,N1695,N1696);
and and784(N1705,N1707,N1708);
and and785(N1706,N1709,N1710);
and and793(N1719,N1721,N1722);
and and794(N1720,N1723,N1724);
and and802(N1733,N1735,N1736);
and and803(N1734,N1737,N1738);
and and811(N1747,N1749,N1750);
and and812(N1748,N1751,N1752);
and and820(N1761,N1763,N1764);
and and821(N1762,N1765,N1766);
and and829(N1775,N1777,N1778);
and and830(N1776,N1779,N1780);
and and838(N1789,N1791,N1792);
and and839(N1790,N1793,N1794);
and and847(N1803,N1805,N1806);
and and848(N1804,N1807,N1808);
and and856(N1817,N1819,N1820);
and and857(N1818,N1821,N1822);
and and865(N1831,N1833,N1834);
and and866(N1832,N1835,N1836);
and and874(N1845,N1847,N1848);
and and875(N1846,N1849,N1850);
and and883(N1859,N1861,N1862);
and and884(N1860,N1863,N1864);
and and892(N1873,N1875,N1876);
and and893(N1874,N1877,N1878);
and and901(N1887,N1889,N1890);
and and902(N1888,N1891,N1892);
and and910(N1901,N1903,N1904);
and and911(N1902,N1905,N1906);
and and919(N1915,N1917,N1918);
and and920(N1916,N1919,N1920);
and and928(N1929,N1931,N1932);
and and929(N1930,N1933,N1934);
and and937(N1943,N1945,N1946);
and and938(N1944,N1947,N1948);
and and946(N1957,N1959,N1960);
and and947(N1958,N1961,N1962);
and and955(N1971,N1973,N1974);
and and956(N1972,N1975,N1976);
and and964(N1985,N1987,N1988);
and and965(N1986,N1989,N1990);
and and973(N1999,N2001,N2002);
and and974(N2000,N2003,N2004);
and and982(N2013,N2015,N2016);
and and983(N2014,N2017,N2018);
and and991(N2027,N2029,N2030);
and and992(N2028,N2031,N2032);
and and1000(N2041,N2043,N2044);
and and1001(N2042,N2045,N2046);
and and1009(N2055,N2057,N2058);
and and1010(N2056,N2059,N2060);
and and1018(N2069,N2071,N2072);
and and1019(N2070,N2073,N2074);
and and1027(N2083,N2085,N2086);
and and1028(N2084,N2087,N2088);
and and1036(N2097,N2099,N2100);
and and1037(N2098,N2101,N2102);
and and1045(N2111,N2113,N2114);
and and1046(N2112,N2115,N2116);
and and1054(N2124,N2126,N2127);
and and1055(N2125,N2128,N2129);
and and1063(N2137,N2139,N2140);
and and1064(N2138,N2141,N2142);
and and1072(N2150,N2152,N2153);
and and1073(N2151,N2154,N2155);
and and1081(N2163,N2165,N2166);
and and1082(N2164,N2167,N2168);
and and1090(N2176,N2178,N2179);
and and1091(N2177,N2180,N2181);
and and1099(N2189,N2191,N2192);
and and1100(N2190,N2193,N2194);
and and1108(N2202,N2204,N2205);
and and1109(N2203,N2206,N2207);
and and1117(N2215,N2217,N2218);
and and1118(N2216,N2219,N2220);
and and1126(N2228,N2230,N2231);
and and1127(N2229,N2232,N2233);
and and1135(N2241,N2243,N2244);
and and1136(N2242,N2245,N2246);
and and1144(N2254,N2256,N2257);
and and1145(N2255,N2258,N2259);
and and1153(N2267,N2269,N2270);
and and1154(N2268,N2271,N2272);
and and1162(N2280,N2282,N2283);
and and1163(N2281,N2284,N2285);
and and1171(N2293,N2295,N2296);
and and1172(N2294,N2297,N2298);
and and1180(N2306,N2308,N2309);
and and1181(N2307,N2310,N2311);
and and1189(N2319,N2321,N2322);
and and1190(N2320,N2323,N2324);
and and1198(N2332,N2334,N2335);
and and1199(N2333,N2336,N2337);
and and1207(N2345,N2347,N2348);
and and1208(N2346,N2349,N2350);
and and1216(N2358,N2360,N2361);
and and1217(N2359,N2362,N2363);
and and1225(N2371,N2373,N2374);
and and1226(N2372,N2375,N2376);
and and1234(N2384,N2386,N2387);
and and1235(N2385,N2388,N2389);
and and1243(N2397,N2399,N2400);
and and1244(N2398,N2401,N2402);
and and1252(N2410,N2412,N2413);
and and1253(N2411,N2414,N2415);
and and1261(N2423,N2425,N2426);
and and1262(N2424,N2427,N2428);
and and1270(N2436,N2438,N2439);
and and1271(N2437,N2440,N2441);
and and1279(N2449,N2451,N2452);
and and1280(N2450,N2453,N2454);
and and1288(N2462,N2464,N2465);
and and1289(N2463,N2466,N2467);
and and1297(N2475,N2477,N2478);
and and1298(N2476,N2479,N2480);
and and1306(N2488,N2490,N2491);
and and1307(N2489,N2492,N2493);
and and1315(N2501,N2503,N2504);
and and1316(N2502,N2505,N2506);
and and1324(N2514,N2516,N2517);
and and1325(N2515,N2518,N2519);
and and1333(N2527,N2529,N2530);
and and1334(N2528,N2531,N2532);
and and1342(N2540,N2542,N2543);
and and1343(N2541,N2544,N2545);
and and1351(N2553,N2555,N2556);
and and1352(N2554,N2557,N2558);
and and1360(N2566,N2568,N2569);
and and1361(N2567,N2570,N2571);
and and1369(N2579,N2581,N2582);
and and1370(N2580,N2583,N2584);
and and1378(N2592,N2594,N2595);
and and1379(N2593,N2596,N2597);
and and1387(N2605,N2607,N2608);
and and1388(N2606,N2609,N2610);
and and1396(N2617,N2619,N2620);
and and1397(N2618,N2621,N2622);
and and1405(N2629,N2631,N2632);
and and1406(N2630,N2633,N2634);
and and1414(N2641,N2643,N2644);
and and1415(N2642,N2645,N2646);
and and1423(N2653,N2655,N2656);
and and1424(N2654,N2657,N2658);
and and1432(N2665,N2667,N2668);
and and1433(N2666,N2669,N2670);
and and1441(N2677,N2679,N2680);
and and1442(N2678,N2681,N2682);
and and1450(N2689,N2691,N2692);
and and1451(N2690,N2693,N2694);
and and1459(N2701,N2703,N2704);
and and1460(N2702,N2705,N2706);
and and1468(N2713,N2715,N2716);
and and1469(N2714,N2717,N2718);
and and1477(N2725,N2727,N2728);
and and1478(N2726,N2729,N2730);
and and1486(N2737,N2739,N2740);
and and1487(N2738,N2741,N2742);
and and1495(N2749,N2751,N2752);
and and1496(N2750,N2753,N2754);
and and1504(N2761,N2763,N2764);
and and1505(N2762,N2765,N2766);
and and1513(N2773,N2775,N2776);
and and1514(N2774,N2777,N2778);
and and1522(N2785,N2787,N2788);
and and1523(N2786,N2789,N2790);
and and1531(N2797,N2799,N2800);
and and1532(N2798,N2801,N2802);
and and1540(N2809,N2811,N2812);
and and1541(N2810,N2813,N2814);
and and1549(N2821,N2823,N2824);
and and1550(N2822,N2825,N2826);
and and1558(N2833,N2835,N2836);
and and1559(N2834,N2837,N2838);
and and1567(N2845,N2847,N2848);
and and1568(N2846,N2849,N2850);
and and1576(N2857,N2859,N2860);
and and1577(N2858,N2861,N2862);
and and1585(N2869,N2871,N2872);
and and1586(N2870,N2873,N2874);
and and1594(N2881,N2883,N2884);
and and1595(N2882,N2885,N2886);
and and1603(N2893,N2895,N2896);
and and1604(N2894,N2897,N2898);
and and1612(N2905,N2907,N2908);
and and1613(N2906,N2909,N2910);
and and1621(N2917,N2919,N2920);
and and1622(N2918,N2921,N2922);
and and1630(N2929,N2931,N2932);
and and1631(N2930,N2933,N2934);
and and1639(N2941,N2943,N2944);
and and1640(N2942,N2945,N2946);
and and1648(N2953,N2955,N2956);
and and1649(N2954,N2957,N2958);
and and1657(N2965,N2967,N2968);
and and1658(N2966,N2969,N2970);
and and1666(N2977,N2979,N2980);
and and1667(N2978,N2981,N2982);
and and1675(N2989,N2991,N2992);
and and1676(N2990,N2993,N2994);
and and1684(N3001,N3003,N3004);
and and1685(N3002,N3005,N3006);
and and1693(N3013,N3015,N3016);
and and1694(N3014,N3017,N3018);
and and1702(N3025,N3027,N3028);
and and1703(N3026,N3029,N3030);
and and1711(N3037,N3039,N3040);
and and1712(N3038,N3041,N3042);
and and1720(N3049,N3051,N3052);
and and1721(N3050,N3053,N3054);
and and1729(N3061,N3063,N3064);
and and1730(N3062,N3065,N3066);
and and1738(N3073,N3075,N3076);
and and1739(N3074,N3077,N3078);
and and1747(N3085,N3087,N3088);
and and1748(N3086,N3089,N3090);
and and1756(N3096,N3098,N3099);
and and1757(N3097,N3100,N3101);
and and1765(N3107,N3109,N3110);
and and1766(N3108,N3111,N3112);
and and1774(N3118,N3120,N3121);
and and1775(N3119,N3122,N3123);
and and1783(N3129,N3131,N3132);
and and1784(N3130,N3133,N3134);
and and1792(N3140,N3142,N3143);
and and1793(N3141,N3144,N3145);
and and1801(N3151,N3153,N3154);
and and1802(N3152,N3155,N3156);
and and1810(N3162,N3164,N3165);
and and1811(N3163,N3166,N3167);
and and1819(N3173,N3175,N3176);
and and1820(N3174,N3177,N3178);
and and1828(N3184,N3186,N3187);
and and1829(N3185,N3188,N3189);
and and1837(N3195,N3197,N3198);
and and1838(N3196,N3199,N3200);
and and1846(N3206,N3208,N3209);
and and1847(N3207,N3210,N3211);
and and1855(N3217,N3219,N3220);
and and1856(N3218,N3221,N3222);
and and1864(N3228,N3230,N3231);
and and1865(N3229,N3232,N3233);
and and1873(N3238,N3240,N3241);
and and1874(N3239,N3242,N3243);
and and1882(N3248,N3250,N3251);
and and1883(N3249,N3252,N3253);
and and1891(N3257,N3259,N3260);
and and1892(N3258,N3261,N3262);
and and1899(N3273,N3275,N3276);
and and1900(N3274,N3277,N3278);
and and1907(N3289,N3291,N3292);
and and1908(N3290,N3293,N3294);
and and1915(N3305,N3307,N3308);
and and1916(N3306,N3309,N3310);
and and1923(N3321,N3323,N3324);
and and1924(N3322,N3325,N3326);
and and1931(N3337,N3339,N3340);
and and1932(N3338,N3341,N3342);
and and1939(N3353,N3355,N3356);
and and1940(N3354,N3357,N3358);
and and1947(N3369,N3371,N3372);
and and1948(N3370,N3373,N3374);
and and1955(N3384,N3386,N3387);
and and1956(N3385,N3388,N3389);
and and1963(N3399,N3401,N3402);
and and1964(N3400,N3403,N3404);
and and1971(N3414,N3416,N3417);
and and1972(N3415,N3418,N3419);
and and1979(N3429,N3431,N3432);
and and1980(N3430,N3433,N3434);
and and1987(N3444,N3446,N3447);
and and1988(N3445,N3448,N3449);
and and1995(N3459,N3461,N3462);
and and1996(N3460,N3463,N3464);
and and2003(N3474,N3476,N3477);
and and2004(N3475,N3478,N3479);
and and2011(N3489,N3491,N3492);
and and2012(N3490,N3493,N3494);
and and2019(N3504,N3506,N3507);
and and2020(N3505,N3508,N3509);
and and2027(N3519,N3521,N3522);
and and2028(N3520,N3523,N3524);
and and2035(N3533,N3535,N3536);
and and2036(N3534,N3537,N3538);
and and2043(N3547,N3549,N3550);
and and2044(N3548,N3551,N3552);
and and2051(N3561,N3563,N3564);
and and2052(N3562,N3565,N3566);
and and2059(N3575,N3577,N3578);
and and2060(N3576,N3579,N3580);
and and2067(N3589,N3591,N3592);
and and2068(N3590,N3593,N3594);
and and2075(N3603,N3605,N3606);
and and2076(N3604,N3607,N3608);
and and2083(N3617,N3619,N3620);
and and2084(N3618,N3621,N3622);
and and2091(N3631,N3633,N3634);
and and2092(N3632,N3635,N3636);
and and2099(N3645,N3647,N3648);
and and2100(N3646,N3649,N3650);
and and2107(N3659,N3661,N3662);
and and2108(N3660,N3663,N3664);
and and2115(N3673,N3675,N3676);
and and2116(N3674,N3677,N3678);
and and2123(N3687,N3689,N3690);
and and2124(N3688,N3691,N3692);
and and2131(N3701,N3703,N3704);
and and2132(N3702,N3705,N3706);
and and2139(N3715,N3717,N3718);
and and2140(N3716,N3719,N3720);
and and2147(N3729,N3731,N3732);
and and2148(N3730,N3733,N3734);
and and2155(N3743,N3745,N3746);
and and2156(N3744,N3747,N3748);
and and2163(N3757,N3759,N3760);
and and2164(N3758,N3761,N3762);
and and2171(N3771,N3773,N3774);
and and2172(N3772,N3775,N3776);
and and2179(N3785,N3787,N3788);
and and2180(N3786,N3789,N3790);
and and2187(N3799,N3801,N3802);
and and2188(N3800,N3803,N3804);
and and2195(N3813,N3815,N3816);
and and2196(N3814,N3817,N3818);
and and2203(N3827,N3829,N3830);
and and2204(N3828,N3831,N3832);
and and2211(N3841,N3843,N3844);
and and2212(N3842,N3845,N3846);
and and2219(N3855,N3857,N3858);
and and2220(N3856,N3859,N3860);
and and2227(N3869,N3871,N3872);
and and2228(N3870,N3873,N3874);
and and2235(N3883,N3885,N3886);
and and2236(N3884,N3887,N3888);
and and2243(N3896,N3898,N3899);
and and2244(N3897,N3900,N3901);
and and2251(N3909,N3911,N3912);
and and2252(N3910,N3913,N3914);
and and2259(N3922,N3924,N3925);
and and2260(N3923,N3926,N3927);
and and2267(N3935,N3937,N3938);
and and2268(N3936,N3939,N3940);
and and2275(N3948,N3950,N3951);
and and2276(N3949,N3952,N3953);
and and2283(N3961,N3963,N3964);
and and2284(N3962,N3965,N3966);
and and2291(N3974,N3976,N3977);
and and2292(N3975,N3978,N3979);
and and2299(N3987,N3989,N3990);
and and2300(N3988,N3991,N3992);
and and2307(N4000,N4002,N4003);
and and2308(N4001,N4004,N4005);
and and2315(N4013,N4015,N4016);
and and2316(N4014,N4017,N4018);
and and2323(N4026,N4028,N4029);
and and2324(N4027,N4030,N4031);
and and2331(N4039,N4041,N4042);
and and2332(N4040,N4043,N4044);
and and2339(N4052,N4054,N4055);
and and2340(N4053,N4056,N4057);
and and2347(N4065,N4067,N4068);
and and2348(N4066,N4069,N4070);
and and2355(N4078,N4080,N4081);
and and2356(N4079,N4082,N4083);
and and2363(N4091,N4093,N4094);
and and2364(N4092,N4095,N4096);
and and2371(N4104,N4106,N4107);
and and2372(N4105,N4108,N4109);
and and2379(N4117,N4119,N4120);
and and2380(N4118,N4121,N4122);
and and2387(N4130,N4132,N4133);
and and2388(N4131,N4134,N4135);
and and2395(N4143,N4145,N4146);
and and2396(N4144,N4147,N4148);
and and2403(N4156,N4158,N4159);
and and2404(N4157,N4160,N4161);
and and2411(N4169,N4171,N4172);
and and2412(N4170,N4173,N4174);
and and2419(N4182,N4184,N4185);
and and2420(N4183,N4186,N4187);
and and2427(N4195,N4197,N4198);
and and2428(N4196,N4199,N4200);
and and2435(N4208,N4210,N4211);
and and2436(N4209,N4212,N4213);
and and2443(N4221,N4223,N4224);
and and2444(N4222,N4225,N4226);
and and2451(N4234,N4236,N4237);
and and2452(N4235,N4238,N4239);
and and2459(N4247,N4249,N4250);
and and2460(N4248,N4251,N4252);
and and2467(N4260,N4262,N4263);
and and2468(N4261,N4264,N4265);
and and2475(N4273,N4275,N4276);
and and2476(N4274,N4277,N4278);
and and2483(N4286,N4288,N4289);
and and2484(N4287,N4290,N4291);
and and2491(N4299,N4301,N4302);
and and2492(N4300,N4303,N4304);
and and2499(N4312,N4314,N4315);
and and2500(N4313,N4316,N4317);
and and2507(N4325,N4327,N4328);
and and2508(N4326,N4329,N4330);
and and2515(N4338,N4340,N4341);
and and2516(N4339,N4342,N4343);
and and2523(N4351,N4353,N4354);
and and2524(N4352,N4355,N4356);
and and2531(N4364,N4366,N4367);
and and2532(N4365,N4368,N4369);
and and2539(N4377,N4379,N4380);
and and2540(N4378,N4381,N4382);
and and2547(N4390,N4392,N4393);
and and2548(N4391,N4394,N4395);
and and2555(N4403,N4405,N4406);
and and2556(N4404,N4407,N4408);
and and2563(N4416,N4418,N4419);
and and2564(N4417,N4420,N4421);
and and2571(N4429,N4431,N4432);
and and2572(N4430,N4433,N4434);
and and2579(N4442,N4444,N4445);
and and2580(N4443,N4446,N4447);
and and2587(N4455,N4457,N4458);
and and2588(N4456,N4459,N4460);
and and2595(N4468,N4470,N4471);
and and2596(N4469,N4472,N4473);
and and2603(N4481,N4483,N4484);
and and2604(N4482,N4485,N4486);
and and2611(N4494,N4496,N4497);
and and2612(N4495,N4498,N4499);
and and2619(N4506,N4508,N4509);
and and2620(N4507,N4510,N4511);
and and2627(N4518,N4520,N4521);
and and2628(N4519,N4522,N4523);
and and2635(N4530,N4532,N4533);
and and2636(N4531,N4534,N4535);
and and2643(N4542,N4544,N4545);
and and2644(N4543,N4546,N4547);
and and2651(N4554,N4556,N4557);
and and2652(N4555,N4558,N4559);
and and2659(N4566,N4568,N4569);
and and2660(N4567,N4570,N4571);
and and2667(N4578,N4580,N4581);
and and2668(N4579,N4582,N4583);
and and2675(N4590,N4592,N4593);
and and2676(N4591,N4594,N4595);
and and2683(N4602,N4604,N4605);
and and2684(N4603,N4606,N4607);
and and2691(N4614,N4616,N4617);
and and2692(N4615,N4618,N4619);
and and2699(N4626,N4628,N4629);
and and2700(N4627,N4630,N4631);
and and2707(N4638,N4640,N4641);
and and2708(N4639,N4642,N4643);
and and2715(N4650,N4652,N4653);
and and2716(N4651,N4654,N4655);
and and2723(N4662,N4664,N4665);
and and2724(N4663,N4666,N4667);
and and2731(N4674,N4676,N4677);
and and2732(N4675,N4678,N4679);
and and2739(N4686,N4688,N4689);
and and2740(N4687,N4690,N4691);
and and2747(N4698,N4700,N4701);
and and2748(N4699,N4702,N4703);
and and2755(N4710,N4712,N4713);
and and2756(N4711,N4714,N4715);
and and2763(N4722,N4724,N4725);
and and2764(N4723,N4726,N4727);
and and2771(N4734,N4736,N4737);
and and2772(N4735,N4738,N4739);
and and2779(N4746,N4748,N4749);
and and2780(N4747,N4750,N4751);
and and2787(N4758,N4760,N4761);
and and2788(N4759,N4762,N4763);
and and2795(N4770,N4772,N4773);
and and2796(N4771,N4774,N4775);
and and2803(N4782,N4784,N4785);
and and2804(N4783,N4786,N4787);
and and2811(N4794,N4796,N4797);
and and2812(N4795,N4798,N4799);
and and2819(N4806,N4808,N4809);
and and2820(N4807,N4810,N4811);
and and2827(N4818,N4820,N4821);
and and2828(N4819,N4822,N4823);
and and2835(N4830,N4832,N4833);
and and2836(N4831,N4834,N4835);
and and2843(N4842,N4844,N4845);
and and2844(N4843,N4846,N4847);
and and2851(N4854,N4856,N4857);
and and2852(N4855,N4858,N4859);
and and2859(N4866,N4868,N4869);
and and2860(N4867,N4870,N4871);
and and2867(N4878,N4880,N4881);
and and2868(N4879,N4882,N4883);
and and2875(N4890,N4892,N4893);
and and2876(N4891,N4894,N4895);
and and2883(N4902,N4904,N4905);
and and2884(N4903,N4906,N4907);
and and2891(N4914,N4916,N4917);
and and2892(N4915,N4918,N4919);
and and2899(N4926,N4928,N4929);
and and2900(N4927,N4930,N4931);
and and2907(N4938,N4940,N4941);
and and2908(N4939,N4942,N4943);
and and2915(N4950,N4952,N4953);
and and2916(N4951,N4954,N4955);
and and2923(N4962,N4964,N4965);
and and2924(N4963,N4966,N4967);
and and2931(N4974,N4976,N4977);
and and2932(N4975,N4978,N4979);
and and2939(N4985,N4987,N4988);
and and2940(N4986,N4989,N4990);
and and2947(N4996,N4998,N4999);
and and2948(N4997,N5000,N5001);
and and2955(N5007,N5009,N5010);
and and2956(N5008,N5011,N5012);
and and2963(N5018,N5020,N5021);
and and2964(N5019,N5022,N5023);
and and2971(N5029,N5031,N5032);
and and2972(N5030,N5033,N5034);
and and2979(N5040,N5042,N5043);
and and2980(N5041,N5044,N5045);
and and2987(N5051,N5053,N5054);
and and2988(N5052,N5055,N5056);
and and2995(N5062,N5064,N5065);
and and2996(N5063,N5066,N5067);
and and3003(N5073,N5075,N5076);
and and3004(N5074,N5077,N5078);
and and3011(N5084,N5086,N5087);
and and3012(N5085,N5088,N5089);
and and3019(N5095,N5097,N5098);
and and3020(N5096,N5099,N5100);
and and3027(N5106,N5108,N5109);
and and3028(N5107,N5110,N5111);
and and3035(N5117,N5119,N5120);
and and3036(N5118,N5121,N5122);
and and3043(N5128,N5130,N5131);
and and3044(N5129,N5132,N5133);
and and3051(N5139,N5141,N5142);
and and3052(N5140,N5143,N5144);
and and3059(N5150,N5152,N5153);
and and3060(N5151,N5154,N5155);
and and3067(N5161,N5163,N5164);
and and3068(N5162,N5165,N5166);
and and3075(N5172,N5174,N5175);
and and3076(N5173,N5176,N5177);
and and3083(N5183,N5185,N5186);
and and3084(N5184,N5187,N5188);
and and3091(N5193,N5195,N5196);
and and3092(N5194,N5197,N5198);
and and3099(N5203,N5205,N5206);
and and3100(N5204,N5207,N5208);
and and3107(N5213,N5215,N5216);
and and3108(N5214,N5217,N5218);
and and3115(N5223,N5225,N5226);
and and3116(N5224,N5227,N5228);
and and3123(N5233,N5235,N5236);
and and3124(N5234,N5237,N5238);
and and3131(N5243,N5245,N5246);
and and3132(N5244,N5247,N5248);
and and3139(N5253,N5255,N5256);
and and3140(N5254,N5257,N5258);
and and3147(N5262,N5264,N5265);
and and3148(N5263,N5266,N5267);
and and3155(N5271,N5273,N5274);
and and3156(N5272,N5275,N5276);
and and3163(N5280,N5282,N5283);
and and3164(N5281,N5284,N5285);
and and3170(N5294,N5296,N5297);
and and3171(N5295,N5298,N5299);
and and3177(N5307,N5309,N5310);
and and3178(N5308,N5311,N5312);
and and3184(N5320,N5322,N5323);
and and3185(N5321,N5324,N5325);
and and3191(N5332,N5334,N5335);
and and3192(N5333,N5336,N5337);
and and3198(N5344,N5346,N5347);
and and3199(N5345,N5348,N5349);
and and3205(N5356,N5358,N5359);
and and3206(N5357,N5360,N5361);
and and3212(N5368,N5370,N5371);
and and3213(N5369,N5372,N5373);
and and3219(N5379,N5381,N5382);
and and3220(N5380,N5383,N5384);
and and3226(N5390,N5392,N5393);
and and3227(N5391,N5394,N5395);
and and3233(N5401,N5403,N5404);
and and3234(N5402,N5405,N5406);
and and3240(N5412,N5414,N5415);
and and3241(N5413,N5416,N5417);
and and3247(N5423,N5425,N5426);
and and3248(N5424,N5427,N5428);
and and3254(N5433,N5435,N5436);
and and3255(N5434,N5437,N5438);
and and3261(N5443,N5445,N5446);
and and3262(N5444,N5447,N5448);
and and3268(N5453,N5455,N5456);
and and3269(N5454,N5457,N5458);
and and3275(N5463,N5465,N5466);
and and3276(N5464,N5467,N5468);
and and3282(N5472,N5474,N5475);
and and3283(N5473,N5476,N5477);
and and3289(N5481,N5483,N5484);
and and3290(N5482,N5485,N5486);
and and3296(N5490,N5492,N5493);
and and3297(N5491,N5494,N5495);
and and3(N391,N395,N396);
and and4(N392,N397,N398);
and and5(N393,N399,N400);
and and6(N394,R2,R3);
and and12(N408,N412,N413);
and and13(N409,in1,N414);
and and14(N410,N415,N416);
and and15(N411,N417,N418);
and and21(N425,N429,N430);
and and22(N426,N431,N432);
and and23(N427,N433,N434);
and and24(N428,N435,N436);
and and30(N442,N446,N447);
and and31(N443,N448,N449);
and and32(N444,N450,N451);
and and33(N445,R1,N452);
and and39(N459,N463,N464);
and and40(N460,N465,N466);
and and41(N461,R0,N467);
and and42(N462,N468,N469);
and and48(N476,N480,N481);
and and49(N477,in1,N482);
and and50(N478,N483,N484);
and and51(N479,N485,N486);
and and57(N492,N496,N497);
and and58(N493,N498,in1);
and and59(N494,N499,N500);
and and60(N495,N501,N502);
and and66(N508,N512,N513);
and and67(N509,N514,in1);
and and68(N510,R0,N515);
and and69(N511,N516,N517);
and and75(N524,N528,N529);
and and76(N525,in0,in1);
and and77(N526,N530,N531);
and and78(N527,N532,N533);
and and84(N540,N544,N545);
and and85(N541,N546,in2);
and and86(N542,N547,N548);
and and87(N543,N549,R3);
and and93(N556,N560,N561);
and and94(N557,N562,in2);
and and95(N558,N563,R1);
and and96(N559,R2,N564);
and and102(N572,N576,N577);
and and103(N573,in1,N578);
and and104(N574,N579,N580);
and and105(N575,R2,N581);
and and111(N588,N592,N593);
and and112(N589,N594,N595);
and and113(N590,R0,R1);
and and114(N591,N596,N597);
and and120(N604,N608,N609);
and and121(N605,N610,N611);
and and122(N606,N612,N613);
and and123(N607,R2,R3);
and and129(N620,N624,N625);
and and130(N621,N626,N627);
and and131(N622,in2,R0);
and and132(N623,N628,R3);
and and138(N636,N640,N641);
and and139(N637,N642,N643);
and and140(N638,N644,N645);
and and141(N639,N646,R3);
and and147(N652,N656,N657);
and and148(N653,N658,in1);
and and149(N654,N659,N660);
and and150(N655,N661,N662);
and and156(N668,N672,N673);
and and157(N669,N674,N675);
and and158(N670,N676,R0);
and and159(N671,N677,N678);
and and165(N684,N688,N689);
and and166(N685,N690,in1);
and and167(N686,N691,R0);
and and168(N687,R2,N692);
and and174(N700,N704,N705);
and and175(N701,N706,N707);
and and176(N702,R0,N708);
and and177(N703,N709,N710);
and and183(N716,N720,N721);
and and184(N717,in0,N722);
and and185(N718,N723,N724);
and and186(N719,N725,R3);
and and192(N732,N736,N737);
and and193(N733,N738,N739);
and and194(N734,N740,N741);
and and195(N735,R1,N742);
and and201(N748,N752,N753);
and and202(N749,N754,in1);
and and203(N750,in2,N755);
and and204(N751,N756,R2);
and and210(N764,N768,N769);
and and211(N765,N770,N771);
and and212(N766,N772,R1);
and and213(N767,N773,N774);
and and219(N780,N784,N785);
and and220(N781,in0,in1);
and and221(N782,N786,N787);
and and222(N783,N788,R3);
and and228(N796,N800,N801);
and and229(N797,N802,N803);
and and230(N798,N804,N805);
and and231(N799,R2,R3);
and and237(N812,N816,N817);
and and238(N813,N818,N819);
and and239(N814,N820,R1);
and and240(N815,R2,R3);
and and246(N827,N831,N832);
and and247(N828,in0,N833);
and and248(N829,N834,R1);
and and249(N830,N835,R3);
and and255(N842,N846,N847);
and and256(N843,N848,N849);
and and257(N844,R0,N850);
and and258(N845,N851,R3);
and and264(N857,N861,N862);
and and265(N858,N863,N864);
and and266(N859,N865,N866);
and and267(N860,R1,R3);
and and273(N872,N876,N877);
and and274(N873,N878,N879);
and and275(N874,N880,N881);
and and276(N875,R1,R2);
and and282(N887,N891,N892);
and and283(N888,N893,N894);
and and284(N889,R0,N895);
and and285(N890,R2,N896);
and and291(N902,N906,N907);
and and292(N903,N908,N909);
and and293(N904,R0,N910);
and and294(N905,R2,R3);
and and300(N917,N921,N922);
and and301(N918,in0,N923);
and and302(N919,N924,R0);
and and303(N920,N925,N926);
and and309(N932,N936,N937);
and and310(N933,N938,N939);
and and311(N934,in2,N940);
and and312(N935,N941,R3);
and and318(N947,N951,N952);
and and319(N948,N953,in1);
and and320(N949,N954,N955);
and and321(N950,R1,N956);
and and327(N962,N966,N967);
and and328(N963,N968,N969);
and and329(N964,N970,R1);
and and330(N965,R2,N971);
and and336(N977,N981,N982);
and and337(N978,in0,in1);
and and338(N979,N983,N984);
and and339(N980,N985,R3);
and and345(N992,N996,N997);
and and346(N993,N998,in2);
and and347(N994,N999,N1000);
and and348(N995,R2,N1001);
and and354(N1007,N1011,N1012);
and and355(N1008,N1013,N1014);
and and356(N1009,in2,N1015);
and and357(N1010,R2,R3);
and and363(N1022,N1026,N1027);
and and364(N1023,in0,N1028);
and and365(N1024,R0,N1029);
and and366(N1025,N1030,R3);
and and372(N1037,N1041,N1042);
and and373(N1038,in1,N1043);
and and374(N1039,R0,N1044);
and and375(N1040,N1045,R3);
and and381(N1052,N1056,N1057);
and and382(N1053,N1058,N1059);
and and383(N1054,in2,R0);
and and384(N1055,N1060,N1061);
and and390(N1067,N1071,N1072);
and and391(N1068,N1073,N1074);
and and392(N1069,N1075,N1076);
and and393(N1070,R2,R3);
and and399(N1082,N1086,N1087);
and and400(N1083,in1,N1088);
and and401(N1084,N1089,R1);
and and402(N1085,N1090,N1091);
and and408(N1097,N1101,N1102);
and and409(N1098,in0,in1);
and and410(N1099,N1103,R1);
and and411(N1100,N1104,N1105);
and and417(N1112,N1116,N1117);
and and418(N1113,N1118,N1119);
and and419(N1114,N1120,R1);
and and420(N1115,R2,N1121);
and and426(N1127,N1131,N1132);
and and427(N1128,N1133,N1134);
and and428(N1129,N1135,R0);
and and429(N1130,R2,N1136);
and and435(N1142,N1146,N1147);
and and436(N1143,in0,in2);
and and437(N1144,N1148,N1149);
and and438(N1145,R2,N1150);
and and444(N1157,N1161,N1162);
and and445(N1158,N1163,in1);
and and446(N1159,in2,R0);
and and447(N1160,N1164,R2);
and and453(N1172,N1176,N1177);
and and454(N1173,N1178,in2);
and and455(N1174,N1179,R1);
and and456(N1175,N1180,N1181);
and and462(N1187,N1191,N1192);
and and463(N1188,N1193,in1);
and and464(N1189,N1194,N1195);
and and465(N1190,R1,N1196);
and and471(N1202,N1206,N1207);
and and472(N1203,in0,N1208);
and and473(N1204,in2,N1209);
and and474(N1205,N1210,R3);
and and480(N1217,N1221,N1222);
and and481(N1218,in0,in1);
and and482(N1219,N1223,N1224);
and and483(N1220,N1225,R3);
and and489(N1232,N1236,N1237);
and and490(N1233,N1238,in1);
and and491(N1234,N1239,R0);
and and492(N1235,N1240,N1241);
and and498(N1247,N1251,N1252);
and and499(N1248,N1253,in1);
and and500(N1249,in2,R0);
and and501(N1250,N1254,N1255);
and and507(N1262,N1266,N1267);
and and508(N1263,N1268,N1269);
and and509(N1264,N1270,R1);
and and510(N1265,N1271,N1272);
and and516(N1277,N1281,N1282);
and and517(N1278,N1283,in1);
and and518(N1279,in2,R0);
and and519(N1280,N1284,N1285);
and and525(N1292,N1296,N1297);
and and526(N1293,N1298,in1);
and and527(N1294,N1299,N1300);
and and528(N1295,R1,R2);
and and534(N1307,N1311,N1312);
and and535(N1308,N1313,N1314);
and and536(N1309,in2,R0);
and and537(N1310,N1315,R2);
and and543(N1322,N1326,N1327);
and and544(N1323,in1,N1328);
and and545(N1324,R0,N1329);
and and546(N1325,R2,N1330);
and and552(N1337,N1341,N1342);
and and553(N1338,N1343,N1344);
and and554(N1339,N1345,R1);
and and555(N1340,R2,N1346);
and and561(N1352,N1356,N1357);
and and562(N1353,N1358,N1359);
and and563(N1354,N1360,N1361);
and and564(N1355,R2,R3);
and and570(N1367,N1371,N1372);
and and571(N1368,N1373,N1374);
and and572(N1369,N1375,R0);
and and573(N1370,R1,R2);
and and579(N1382,N1386,N1387);
and and580(N1383,N1388,N1389);
and and581(N1384,in2,N1390);
and and582(N1385,N1391,R2);
and and588(N1397,N1401,N1402);
and and589(N1398,N1403,in2);
and and590(N1399,N1404,R1);
and and591(N1400,R2,N1405);
and and597(N1412,N1416,N1417);
and and598(N1413,N1418,N1419);
and and599(N1414,N1420,N1421);
and and600(N1415,R2,R3);
and and606(N1427,N1431,N1432);
and and607(N1428,in0,N1433);
and and608(N1429,N1434,R1);
and and609(N1430,N1435,R3);
and and615(N1441,N1445,N1446);
and and616(N1442,N1447,N1448);
and and617(N1443,in2,N1449);
and and618(N1444,R1,N1450);
and and624(N1455,N1459,N1460);
and and625(N1456,N1461,in1);
and and626(N1457,in2,N1462);
and and627(N1458,R2,R3);
and and633(N1469,N1473,N1474);
and and634(N1470,in0,N1475);
and and635(N1471,in2,N1476);
and and636(N1472,R1,R2);
and and642(N1483,N1487,N1488);
and and643(N1484,in1,in2);
and and644(N1485,N1489,R1);
and and645(N1486,R2,R3);
and and651(N1497,N1501,N1502);
and and652(N1498,N1503,N1504);
and and653(N1499,N1505,R1);
and and654(N1500,N1506,R3);
and and660(N1511,N1515,N1516);
and and661(N1512,in1,N1517);
and and662(N1513,N1518,R1);
and and663(N1514,N1519,R3);
and and669(N1525,N1529,N1530);
and and670(N1526,in0,in1);
and and671(N1527,R0,N1531);
and and672(N1528,R2,N1532);
and and678(N1539,N1543,N1544);
and and679(N1540,in0,in2);
and and680(N1541,R0,N1545);
and and681(N1542,N1546,R3);
and and687(N1553,N1557,N1558);
and and688(N1554,in0,in1);
and and689(N1555,N1559,R0);
and and690(N1556,R1,R2);
and and696(N1567,N1571,N1572);
and and697(N1568,in0,in1);
and and698(N1569,in2,R1);
and and699(N1570,R2,N1573);
and and705(N1581,N1585,N1586);
and and706(N1582,in0,in1);
and and707(N1583,N1587,R0);
and and708(N1584,R1,N1588);
and and714(N1595,N1599,N1600);
and and715(N1596,N1601,in1);
and and716(N1597,in2,N1602);
and and717(N1598,R2,R3);
and and723(N1609,N1613,N1614);
and and724(N1610,N1615,N1616);
and and725(N1611,R0,N1617);
and and726(N1612,N1618,R3);
and and732(N1623,N1627,N1628);
and and733(N1624,N1629,in2);
and and734(N1625,N1630,N1631);
and and735(N1626,R2,R3);
and and741(N1637,N1641,N1642);
and and742(N1638,in1,N1643);
and and743(N1639,N1644,R1);
and and744(N1640,R2,R3);
and and750(N1651,N1655,N1656);
and and751(N1652,in0,N1657);
and and752(N1653,N1658,N1659);
and and753(N1654,R1,R2);
and and759(N1665,N1669,N1670);
and and760(N1666,N1671,in2);
and and761(N1667,R0,R1);
and and762(N1668,R2,N1672);
and and768(N1679,N1683,N1684);
and and769(N1680,N1685,in1);
and and770(N1681,N1686,N1687);
and and771(N1682,R2,R3);
and and777(N1693,N1697,N1698);
and and778(N1694,in1,N1699);
and and779(N1695,N1700,R1);
and and780(N1696,R2,N1701);
and and786(N1707,N1711,N1712);
and and787(N1708,in0,in2);
and and788(N1709,N1713,N1714);
and and789(N1710,N1715,R3);
and and795(N1721,N1725,N1726);
and and796(N1722,in0,in1);
and and797(N1723,N1727,N1728);
and and798(N1724,N1729,R3);
and and804(N1735,N1739,N1740);
and and805(N1736,in1,N1741);
and and806(N1737,R0,N1742);
and and807(N1738,R2,N1743);
and and813(N1749,N1753,N1754);
and and814(N1750,N1755,in1);
and and815(N1751,N1756,R0);
and and816(N1752,N1757,N1758);
and and822(N1763,N1767,N1768);
and and823(N1764,in1,N1769);
and and824(N1765,N1770,N1771);
and and825(N1766,R2,R3);
and and831(N1777,N1781,N1782);
and and832(N1778,N1783,in1);
and and833(N1779,N1784,R1);
and and834(N1780,N1785,R3);
and and840(N1791,N1795,N1796);
and and841(N1792,N1797,in1);
and and842(N1793,in2,N1798);
and and843(N1794,N1799,R2);
and and849(N1805,N1809,N1810);
and and850(N1806,N1811,N1812);
and and851(N1807,N1813,R0);
and and852(N1808,R1,N1814);
and and858(N1819,N1823,N1824);
and and859(N1820,in0,in1);
and and860(N1821,N1825,N1826);
and and861(N1822,N1827,R3);
and and867(N1833,N1837,N1838);
and and868(N1834,N1839,in1);
and and869(N1835,in2,N1840);
and and870(N1836,N1841,N1842);
and and876(N1847,N1851,N1852);
and and877(N1848,in0,in1);
and and878(N1849,in2,R0);
and and879(N1850,N1853,R2);
and and885(N1861,N1865,N1866);
and and886(N1862,N1867,in1);
and and887(N1863,N1868,N1869);
and and888(N1864,N1870,R3);
and and894(N1875,N1879,N1880);
and and895(N1876,in1,N1881);
and and896(N1877,N1882,R1);
and and897(N1878,R2,R3);
and and903(N1889,N1893,N1894);
and and904(N1890,N1895,in1);
and and905(N1891,N1896,R0);
and and906(N1892,R1,N1897);
and and912(N1903,N1907,N1908);
and and913(N1904,N1909,N1910);
and and914(N1905,R0,R1);
and and915(N1906,N1911,R3);
and and921(N1917,N1921,N1922);
and and922(N1918,N1923,N1924);
and and923(N1919,R0,N1925);
and and924(N1920,R2,N1926);
and and930(N1931,N1935,N1936);
and and931(N1932,N1937,N1938);
and and932(N1933,R0,N1939);
and and933(N1934,R2,N1940);
and and939(N1945,N1949,N1950);
and and940(N1946,N1951,in1);
and and941(N1947,N1952,R1);
and and942(N1948,N1953,N1954);
and and948(N1959,N1963,N1964);
and and949(N1960,N1965,N1966);
and and950(N1961,in2,N1967);
and and951(N1962,R2,N1968);
and and957(N1973,N1977,N1978);
and and958(N1974,N1979,N1980);
and and959(N1975,N1981,N1982);
and and960(N1976,R1,N1983);
and and966(N1987,N1991,N1992);
and and967(N1988,in0,in1);
and and968(N1989,N1993,R1);
and and969(N1990,R2,N1994);
and and975(N2001,N2005,N2006);
and and976(N2002,N2007,in1);
and and977(N2003,in2,N2008);
and and978(N2004,R2,R3);
and and984(N2015,N2019,N2020);
and and985(N2016,in0,in1);
and and986(N2017,N2021,N2022);
and and987(N2018,R2,R3);
and and993(N2029,N2033,N2034);
and and994(N2030,N2035,N2036);
and and995(N2031,in2,R0);
and and996(N2032,R1,N2037);
and and1002(N2043,N2047,N2048);
and and1003(N2044,N2049,N2050);
and and1004(N2045,in2,R0);
and and1005(N2046,N2051,R2);
and and1011(N2057,N2061,N2062);
and and1012(N2058,in1,N2063);
and and1013(N2059,R0,R1);
and and1014(N2060,R2,N2064);
and and1020(N2071,N2075,N2076);
and and1021(N2072,N2077,N2078);
and and1022(N2073,in2,N2079);
and and1023(N2074,N2080,R2);
and and1029(N2085,N2089,N2090);
and and1030(N2086,N2091,in1);
and and1031(N2087,R0,R1);
and and1032(N2088,R2,N2092);
and and1038(N2099,N2103,N2104);
and and1039(N2100,N2105,N2106);
and and1040(N2101,in2,R0);
and and1041(N2102,R1,N2107);
and and1047(N2113,N2117,N2118);
and and1048(N2114,in0,in2);
and and1049(N2115,R0,R1);
and and1050(N2116,R2,R3);
and and1056(N2126,N2130,N2131);
and and1057(N2127,in0,in1);
and and1058(N2128,in2,R0);
and and1059(N2129,R1,N2132);
and and1065(N2139,N2143,N2144);
and and1066(N2140,in1,in2);
and and1067(N2141,R0,N2145);
and and1068(N2142,R2,R3);
and and1074(N2152,N2156,N2157);
and and1075(N2153,N2158,in2);
and and1076(N2154,N2159,R1);
and and1077(N2155,R2,R3);
and and1083(N2165,N2169,N2170);
and and1084(N2166,N2171,N2172);
and and1085(N2167,N2173,R1);
and and1086(N2168,R2,R3);
and and1092(N2178,N2182,N2183);
and and1093(N2179,in0,in2);
and and1094(N2180,R0,N2184);
and and1095(N2181,R2,N2185);
and and1101(N2191,N2195,N2196);
and and1102(N2192,N2197,in1);
and and1103(N2193,in2,R0);
and and1104(N2194,N2198,R2);
and and1110(N2204,N2208,N2209);
and and1111(N2205,N2210,in1);
and and1112(N2206,in2,R0);
and and1113(N2207,R1,N2211);
and and1119(N2217,N2221,N2222);
and and1120(N2218,N2223,in2);
and and1121(N2219,R0,N2224);
and and1122(N2220,R2,R3);
and and1128(N2230,N2234,N2235);
and and1129(N2231,in0,in1);
and and1130(N2232,in2,N2236);
and and1131(N2233,R2,N2237);
and and1137(N2243,N2247,N2248);
and and1138(N2244,in0,in1);
and and1139(N2245,in2,N2249);
and and1140(N2246,R2,R3);
and and1146(N2256,N2260,N2261);
and and1147(N2257,N2262,N2263);
and and1148(N2258,in2,R0);
and and1149(N2259,N2264,R3);
and and1155(N2269,N2273,N2274);
and and1156(N2270,N2275,N2276);
and and1157(N2271,in2,R0);
and and1158(N2272,R1,N2277);
and and1164(N2282,N2286,N2287);
and and1165(N2283,in0,in1);
and and1166(N2284,in2,R0);
and and1167(N2285,N2288,N2289);
and and1173(N2295,N2299,N2300);
and and1174(N2296,N2301,in2);
and and1175(N2297,R0,R1);
and and1176(N2298,R2,R3);
and and1182(N2308,N2312,N2313);
and and1183(N2309,N2314,in2);
and and1184(N2310,N2315,R1);
and and1185(N2311,R2,R3);
and and1191(N2321,N2325,N2326);
and and1192(N2322,N2327,in1);
and and1193(N2323,N2328,R0);
and and1194(N2324,R1,R2);
and and1200(N2334,N2338,N2339);
and and1201(N2335,N2340,in1);
and and1202(N2336,in2,R1);
and and1203(N2337,N2341,N2342);
and and1209(N2347,N2351,N2352);
and and1210(N2348,in0,N2353);
and and1211(N2349,in2,N2354);
and and1212(N2350,N2355,R2);
and and1218(N2360,N2364,N2365);
and and1219(N2361,in0,N2366);
and and1220(N2362,in2,R1);
and and1221(N2363,N2367,R3);
and and1227(N2373,N2377,N2378);
and and1228(N2374,in0,in1);
and and1229(N2375,N2379,N2380);
and and1230(N2376,N2381,R2);
and and1236(N2386,N2390,N2391);
and and1237(N2387,in0,N2392);
and and1238(N2388,in2,R0);
and and1239(N2389,N2393,R2);
and and1245(N2399,N2403,N2404);
and and1246(N2400,in0,in1);
and and1247(N2401,in2,R0);
and and1248(N2402,N2405,N2406);
and and1254(N2412,N2416,N2417);
and and1255(N2413,in0,N2418);
and and1256(N2414,N2419,R0);
and and1257(N2415,R2,R3);
and and1263(N2425,N2429,N2430);
and and1264(N2426,N2431,in1);
and and1265(N2427,N2432,R0);
and and1266(N2428,R2,R3);
and and1272(N2438,N2442,N2443);
and and1273(N2439,N2444,in2);
and and1274(N2440,N2445,R1);
and and1275(N2441,R2,R3);
and and1281(N2451,N2455,N2456);
and and1282(N2452,in0,in1);
and and1283(N2453,in2,N2457);
and and1284(N2454,R1,N2458);
and and1290(N2464,N2468,N2469);
and and1291(N2465,in0,N2470);
and and1292(N2466,N2471,R1);
and and1293(N2467,N2472,R3);
and and1299(N2477,N2481,N2482);
and and1300(N2478,in1,N2483);
and and1301(N2479,N2484,R1);
and and1302(N2480,N2485,R3);
and and1308(N2490,N2494,N2495);
and and1309(N2491,N2496,in1);
and and1310(N2492,in2,R0);
and and1311(N2493,N2497,R2);
and and1317(N2503,N2507,N2508);
and and1318(N2504,N2509,in1);
and and1319(N2505,N2510,N2511);
and and1320(N2506,R1,R2);
and and1326(N2516,N2520,N2521);
and and1327(N2517,in0,N2522);
and and1328(N2518,in2,R0);
and and1329(N2519,R1,N2523);
and and1335(N2529,N2533,N2534);
and and1336(N2530,in0,in2);
and and1337(N2531,R0,R1);
and and1338(N2532,R2,N2535);
and and1344(N2542,N2546,N2547);
and and1345(N2543,N2548,in1);
and and1346(N2544,in2,R0);
and and1347(N2545,N2549,N2550);
and and1353(N2555,N2559,N2560);
and and1354(N2556,N2561,N2562);
and and1355(N2557,in2,R0);
and and1356(N2558,N2563,R2);
and and1362(N2568,N2572,N2573);
and and1363(N2569,N2574,N2575);
and and1364(N2570,N2576,R0);
and and1365(N2571,R1,R2);
and and1371(N2581,N2585,N2586);
and and1372(N2582,N2587,in1);
and and1373(N2583,in2,R0);
and and1374(N2584,N2588,R3);
and and1380(N2594,N2598,N2599);
and and1381(N2595,N2600,in1);
and and1382(N2596,N2601,N2602);
and and1383(N2597,R1,R3);
and and1389(N2607,N2611,N2612);
and and1390(N2608,in1,in2);
and and1391(N2609,R0,R1);
and and1392(N2610,R2,N2613);
and and1398(N2619,N2623,N2624);
and and1399(N2620,in0,in1);
and and1400(N2621,in2,N2625);
and and1401(N2622,R1,N2626);
and and1407(N2631,N2635,N2636);
and and1408(N2632,N2637,in1);
and and1409(N2633,in2,R1);
and and1410(N2634,R2,R3);
and and1416(N2643,N2647,N2648);
and and1417(N2644,in1,in2);
and and1418(N2645,R0,R1);
and and1419(N2646,R2,N2649);
and and1425(N2655,N2659,N2660);
and and1426(N2656,in0,in1);
and and1427(N2657,R0,R1);
and and1428(N2658,R2,N2661);
and and1434(N2667,N2671,N2672);
and and1435(N2668,in0,in1);
and and1436(N2669,R0,N2673);
and and1437(N2670,R2,R3);
and and1443(N2679,N2683,N2684);
and and1444(N2680,N2685,in1);
and and1445(N2681,in2,N2686);
and and1446(N2682,R2,R3);
and and1452(N2691,N2695,N2696);
and and1453(N2692,in1,in2);
and and1454(N2693,R0,R1);
and and1455(N2694,N2697,N2698);
and and1461(N2703,N2707,N2708);
and and1462(N2704,in0,in1);
and and1463(N2705,in2,N2709);
and and1464(N2706,R1,R2);
and and1470(N2715,N2719,N2720);
and and1471(N2716,N2721,in1);
and and1472(N2717,R0,R1);
and and1473(N2718,R2,N2722);
and and1479(N2727,N2731,N2732);
and and1480(N2728,in0,in1);
and and1481(N2729,N2733,R0);
and and1482(N2730,R2,N2734);
and and1488(N2739,N2743,N2744);
and and1489(N2740,in0,in2);
and and1490(N2741,R0,N2745);
and and1491(N2742,N2746,R3);
and and1497(N2751,N2755,N2756);
and and1498(N2752,in0,in1);
and and1499(N2753,R0,N2757);
and and1500(N2754,N2758,R3);
and and1506(N2763,N2767,N2768);
and and1507(N2764,in0,in1);
and and1508(N2765,in2,N2769);
and and1509(N2766,N2770,R2);
and and1515(N2775,N2779,N2780);
and and1516(N2776,N2781,in1);
and and1517(N2777,N2782,R0);
and and1518(N2778,R1,R2);
and and1524(N2787,N2791,N2792);
and and1525(N2788,in0,in1);
and and1526(N2789,N2793,R0);
and and1527(N2790,R1,R2);
and and1533(N2799,N2803,N2804);
and and1534(N2800,in0,in1);
and and1535(N2801,in2,R0);
and and1536(N2802,R1,N2805);
and and1542(N2811,N2815,N2816);
and and1543(N2812,in0,in1);
and and1544(N2813,in2,R0);
and and1545(N2814,N2817,R2);
and and1551(N2823,N2827,N2828);
and and1552(N2824,in0,in1);
and and1553(N2825,in2,N2829);
and and1554(N2826,N2830,R2);
and and1560(N2835,N2839,N2840);
and and1561(N2836,in0,in1);
and and1562(N2837,in2,N2841);
and and1563(N2838,R1,N2842);
and and1569(N2847,N2851,N2852);
and and1570(N2848,N2853,in1);
and and1571(N2849,in2,N2854);
and and1572(N2850,R1,N2855);
and and1578(N2859,N2863,N2864);
and and1579(N2860,in0,in1);
and and1580(N2861,N2865,N2866);
and and1581(N2862,R1,R2);
and and1587(N2871,N2875,N2876);
and and1588(N2872,N2877,in1);
and and1589(N2873,in2,R0);
and and1590(N2874,R1,R2);
and and1596(N2883,N2887,N2888);
and and1597(N2884,N2889,N2890);
and and1598(N2885,N2891,R0);
and and1599(N2886,R1,R2);
and and1605(N2895,N2899,N2900);
and and1606(N2896,N2901,N2902);
and and1607(N2897,N2903,R0);
and and1608(N2898,R1,R2);
and and1614(N2907,N2911,N2912);
and and1615(N2908,in0,in1);
and and1616(N2909,in2,N2913);
and and1617(N2910,R1,R2);
and and1623(N2919,N2923,N2924);
and and1624(N2920,N2925,N2926);
and and1625(N2921,in2,R0);
and and1626(N2922,R1,N2927);
and and1632(N2931,N2935,N2936);
and and1633(N2932,N2937,in1);
and and1634(N2933,in2,R0);
and and1635(N2934,N2938,R2);
and and1641(N2943,N2947,N2948);
and and1642(N2944,N2949,in1);
and and1643(N2945,N2950,R1);
and and1644(N2946,R2,R3);
and and1650(N2955,N2959,N2960);
and and1651(N2956,N2961,in1);
and and1652(N2957,N2962,R0);
and and1653(N2958,R1,R2);
and and1659(N2967,N2971,N2972);
and and1660(N2968,N2973,N2974);
and and1661(N2969,in2,R0);
and and1662(N2970,R1,R2);
and and1668(N2979,N2983,N2984);
and and1669(N2980,N2985,in1);
and and1670(N2981,in2,R0);
and and1671(N2982,R2,N2986);
and and1677(N2991,N2995,N2996);
and and1678(N2992,N2997,N2998);
and and1679(N2993,in2,N2999);
and and1680(N2994,R1,R3);
and and1686(N3003,N3007,N3008);
and and1687(N3004,in0,in1);
and and1688(N3005,in2,N3009);
and and1689(N3006,N3010,R2);
and and1695(N3015,N3019,N3020);
and and1696(N3016,in0,in1);
and and1697(N3017,in2,R0);
and and1698(N3018,R2,R3);
and and1704(N3027,N3031,N3032);
and and1705(N3028,N3033,in1);
and and1706(N3029,in2,N3034);
and and1707(N3030,R1,R2);
and and1713(N3039,N3043,N3044);
and and1714(N3040,in0,in1);
and and1715(N3041,R0,R1);
and and1716(N3042,R2,N3045);
and and1722(N3051,N3055,N3056);
and and1723(N3052,in0,in1);
and and1724(N3053,in2,R0);
and and1725(N3054,R1,N3057);
and and1731(N3063,N3067,N3068);
and and1732(N3064,N3069,in1);
and and1733(N3065,N3070,R0);
and and1734(N3066,R1,R2);
and and1740(N3075,N3079,N3080);
and and1741(N3076,N3081,in1);
and and1742(N3077,in2,R0);
and and1743(N3078,R1,R2);
and and1749(N3087,N3091,N3092);
and and1750(N3088,in0,in2);
and and1751(N3089,R0,R1);
and and1752(N3090,N3093,R3);
and and1758(N3098,N3102,N3103);
and and1759(N3099,in0,in2);
and and1760(N3100,R0,R1);
and and1761(N3101,R2,R3);
and and1767(N3109,N3113,N3114);
and and1768(N3110,N3115,in1);
and and1769(N3111,in2,R0);
and and1770(N3112,R1,R2);
and and1776(N3120,N3124,N3125);
and and1777(N3121,in0,in2);
and and1778(N3122,R0,N3126);
and and1779(N3123,R2,R3);
and and1785(N3131,N3135,N3136);
and and1786(N3132,in0,in2);
and and1787(N3133,R0,R1);
and and1788(N3134,R2,R3);
and and1794(N3142,N3146,N3147);
and and1795(N3143,in1,in2);
and and1796(N3144,R0,R1);
and and1797(N3145,R2,R3);
and and1803(N3153,N3157,N3158);
and and1804(N3154,in0,in1);
and and1805(N3155,in2,R0);
and and1806(N3156,R1,R2);
and and1812(N3164,N3168,N3169);
and and1813(N3165,N3170,in1);
and and1814(N3166,in2,R0);
and and1815(N3167,N3171,R2);
and and1821(N3175,N3179,N3180);
and and1822(N3176,in0,in1);
and and1823(N3177,in2,R0);
and and1824(N3178,N3181,R2);
and and1830(N3186,N3190,N3191);
and and1831(N3187,in1,in2);
and and1832(N3188,N3192,R1);
and and1833(N3189,R2,R3);
and and1839(N3197,N3201,N3202);
and and1840(N3198,in0,N3203);
and and1841(N3199,in2,N3204);
and and1842(N3200,R1,R2);
and and1848(N3208,N3212,N3213);
and and1849(N3209,N3214,in1);
and and1850(N3210,in2,N3215);
and and1851(N3211,R1,R2);
and and1857(N3219,N3223,N3224);
and and1858(N3220,in0,in1);
and and1859(N3221,in2,R0);
and and1860(N3222,R1,R2);
and and1866(N3230,N3234,N3235);
and and1867(N3231,in1,N3236);
and and1868(N3232,R0,R1);
and and1869(N3233,R2,R3);
and and1875(N3240,N3244,N3245);
and and1876(N3241,in0,in1);
and and1877(N3242,N3246,R1);
and and1878(N3243,R2,R3);
and and1884(N3250,N3254,N3255);
and and1885(N3251,in0,in1);
and and1886(N3252,in2,R0);
and and1887(N3253,R1,R3);
and and1893(N3259,N3263,N3264);
and and1894(N3260,N3265,in2);
and and1895(N3261,N3266,N3267);
and and1896(N3262,N3268,N3269);
and and1901(N3275,N3279,N3280);
and and1902(N3276,N3281,N3282);
and and1903(N3277,N3283,N3284);
and and1904(N3278,N3285,N3286);
and and1909(N3291,N3295,N3296);
and and1910(N3292,N3297,N3298);
and and1911(N3293,N3299,N3300);
and and1912(N3294,N3301,R4);
and and1917(N3307,N3311,N3312);
and and1918(N3308,N3313,N3314);
and and1919(N3309,N3315,R2);
and and1920(N3310,N3316,N3317);
and and1925(N3323,N3327,N3328);
and and1926(N3324,N3329,N3330);
and and1927(N3325,N3331,N3332);
and and1928(N3326,R3,N3333);
and and1933(N3339,N3343,N3344);
and and1934(N3340,N3345,R0);
and and1935(N3341,N3346,N3347);
and and1936(N3342,N3348,N3349);
and and1941(N3355,N3359,N3360);
and and1942(N3356,N3361,N3362);
and and1943(N3357,N3363,N3364);
and and1944(N3358,N3365,N3366);
and and1949(N3371,N3375,N3376);
and and1950(N3372,in2,N3377);
and and1951(N3373,N3378,N3379);
and and1952(N3374,N3380,N3381);
and and1957(N3386,N3390,N3391);
and and1958(N3387,N3392,N3393);
and and1959(N3388,N3394,R2);
and and1960(N3389,R4,N3395);
and and1965(N3401,N3405,N3406);
and and1966(N3402,N3407,N3408);
and and1967(N3403,R1,R2);
and and1968(N3404,N3409,N3410);
and and1973(N3416,N3420,N3421);
and and1974(N3417,in1,in2);
and and1975(N3418,N3422,N3423);
and and1976(N3419,N3424,N3425);
and and1981(N3431,N3435,N3436);
and and1982(N3432,N3437,N3438);
and and1983(N3433,R1,N3439);
and and1984(N3434,N3440,N3441);
and and1989(N3446,N3450,N3451);
and and1990(N3447,N3452,R0);
and and1991(N3448,N3453,N3454);
and and1992(N3449,R4,N3455);
and and1997(N3461,N3465,N3466);
and and1998(N3462,in1,N3467);
and and1999(N3463,N3468,N3469);
and and2000(N3464,R3,N3470);
and and2005(N3476,N3480,in0);
and and2006(N3477,N3481,N3482);
and and2007(N3478,N3483,N3484);
and and2008(N3479,R3,N3485);
and and2013(N3491,N3495,N3496);
and and2014(N3492,N3497,N3498);
and and2015(N3493,R1,N3499);
and and2016(N3494,N3500,N3501);
and and2021(N3506,N3510,N3511);
and and2022(N3507,N3512,in2);
and and2023(N3508,N3513,N3514);
and and2024(N3509,N3515,R4);
and and2029(N3521,N3525,N3526);
and and2030(N3522,in1,N3527);
and and2031(N3523,N3528,R2);
and and2032(N3524,N3529,N3530);
and and2037(N3535,N3539,N3540);
and and2038(N3536,N3541,R0);
and and2039(N3537,N3542,R3);
and and2040(N3538,N3543,R5);
and and2045(N3549,N3553,N3554);
and and2046(N3550,in2,N3555);
and and2047(N3551,R2,N3556);
and and2048(N3552,R4,N3557);
and and2053(N3563,N3567,in1);
and and2054(N3564,N3568,N3569);
and and2055(N3565,R1,R2);
and and2056(N3566,N3570,N3571);
and and2061(N3577,N3581,in0);
and and2062(N3578,N3582,N3583);
and and2063(N3579,N3584,R1);
and and2064(N3580,R2,N3585);
and and2069(N3591,N3595,in0);
and and2070(N3592,N3596,N3597);
and and2071(N3593,R2,N3598);
and and2072(N3594,N3599,N3600);
and and2077(N3605,N3609,in0);
and and2078(N3606,N3610,N3611);
and and2079(N3607,R2,R3);
and and2080(N3608,N3612,N3613);
and and2085(N3619,N3623,in0);
and and2086(N3620,in2,N3624);
and and2087(N3621,N3625,N3626);
and and2088(N3622,N3627,N3628);
and and2093(N3633,N3637,N3638);
and and2094(N3634,in1,N3639);
and and2095(N3635,R0,R3);
and and2096(N3636,N3640,N3641);
and and2101(N3647,N3651,N3652);
and and2102(N3648,in1,N3653);
and and2103(N3649,R0,N3654);
and and2104(N3650,N3655,N3656);
and and2109(N3661,N3665,N3666);
and and2110(N3662,in2,R0);
and and2111(N3663,R1,N3667);
and and2112(N3664,N3668,N3669);
and and2117(N3675,N3679,in0);
and and2118(N3676,N3680,R0);
and and2119(N3677,R1,N3681);
and and2120(N3678,N3682,N3683);
and and2125(N3689,N3693,in1);
and and2126(N3690,N3694,N3695);
and and2127(N3691,N3696,R2);
and and2128(N3692,N3697,N3698);
and and2133(N3703,N3707,in0);
and and2134(N3704,N3708,N3709);
and and2135(N3705,N3710,R2);
and and2136(N3706,N3711,N3712);
and and2141(N3717,N3721,in0);
and and2142(N3718,N3722,R0);
and and2143(N3719,R2,N3723);
and and2144(N3720,N3724,N3725);
and and2149(N3731,N3735,N3736);
and and2150(N3732,N3737,N3738);
and and2151(N3733,N3739,R3);
and and2152(N3734,N3740,R5);
and and2157(N3745,N3749,N3750);
and and2158(N3746,N3751,in2);
and and2159(N3747,N3752,R1);
and and2160(N3748,N3753,N3754);
and and2165(N3759,N3763,in0);
and and2166(N3760,in2,R0);
and and2167(N3761,N3764,N3765);
and and2168(N3762,N3766,N3767);
and and2173(N3773,N3777,in0);
and and2174(N3774,in1,N3778);
and and2175(N3775,R0,N3779);
and and2176(N3776,N3780,N3781);
and and2181(N3787,N3791,in0);
and and2182(N3788,in2,N3792);
and and2183(N3789,N3793,N3794);
and and2184(N3790,N3795,N3796);
and and2189(N3801,N3805,N3806);
and and2190(N3802,in2,N3807);
and and2191(N3803,R1,N3808);
and and2192(N3804,N3809,N3810);
and and2197(N3815,N3819,N3820);
and and2198(N3816,in1,N3821);
and and2199(N3817,R0,N3822);
and and2200(N3818,N3823,R4);
and and2205(N3829,N3833,N3834);
and and2206(N3830,in2,N3835);
and and2207(N3831,R2,N3836);
and and2208(N3832,R4,N3837);
and and2213(N3843,N3847,in0);
and and2214(N3844,N3848,N3849);
and and2215(N3845,R1,N3850);
and and2216(N3846,N3851,N3852);
and and2221(N3857,N3861,N3862);
and and2222(N3858,in1,N3863);
and and2223(N3859,R1,N3864);
and and2224(N3860,N3865,N3866);
and and2229(N3871,N3875,N3876);
and and2230(N3872,N3877,in2);
and and2231(N3873,R1,N3878);
and and2232(N3874,N3879,N3880);
and and2237(N3885,N3889,in1);
and and2238(N3886,N3890,N3891);
and and2239(N3887,R1,R3);
and and2240(N3888,R4,N3892);
and and2245(N3898,N3902,in0);
and and2246(N3899,N3903,N3904);
and and2247(N3900,R2,R3);
and and2248(N3901,R4,N3905);
and and2253(N3911,N3915,in0);
and and2254(N3912,N3916,R0);
and and2255(N3913,R1,R3);
and and2256(N3914,N3917,N3918);
and and2261(N3924,N3928,N3929);
and and2262(N3925,in2,R0);
and and2263(N3926,R1,N3930);
and and2264(N3927,R3,N3931);
and and2269(N3937,N3941,N3942);
and and2270(N3938,N3943,N3944);
and and2271(N3939,R0,R1);
and and2272(N3940,R2,R4);
and and2277(N3950,N3954,N3955);
and and2278(N3951,R0,R1);
and and2279(N3952,N3956,R3);
and and2280(N3953,R4,N3957);
and and2285(N3963,N3967,N3968);
and and2286(N3964,N3969,N3970);
and and2287(N3965,R0,R1);
and and2288(N3966,N3971,R3);
and and2293(N3976,N3980,in0);
and and2294(N3977,N3981,N3982);
and and2295(N3978,R2,N3983);
and and2296(N3979,R4,R5);
and and2301(N3989,N3993,in1);
and and2302(N3990,N3994,N3995);
and and2303(N3991,N3996,R2);
and and2304(N3992,R3,N3997);
and and2309(N4002,N4006,in0);
and and2310(N4003,N4007,N4008);
and and2311(N4004,R2,R3);
and and2312(N4005,N4009,N4010);
and and2317(N4015,N4019,in0);
and and2318(N4016,N4020,R0);
and and2319(N4017,R1,N4021);
and and2320(N4018,R4,N4022);
and and2325(N4028,N4032,N4033);
and and2326(N4029,in2,R0);
and and2327(N4030,R1,N4034);
and and2328(N4031,N4035,N4036);
and and2333(N4041,N4045,in0);
and and2334(N4042,N4046,R1);
and and2335(N4043,R2,N4047);
and and2336(N4044,R4,N4048);
and and2341(N4054,N4058,in0);
and and2342(N4055,in1,N4059);
and and2343(N4056,R0,N4060);
and and2344(N4057,N4061,N4062);
and and2349(N4067,N4071,in0);
and and2350(N4068,N4072,N4073);
and and2351(N4069,N4074,R3);
and and2352(N4070,N4075,R5);
and and2357(N4080,N4084,N4085);
and and2358(N4081,in2,N4086);
and and2359(N4082,N4087,R3);
and and2360(N4083,N4088,R5);
and and2365(N4093,N4097,N4098);
and and2366(N4094,N4099,N4100);
and and2367(N4095,N4101,R2);
and and2368(N4096,R3,R4);
and and2373(N4106,N4110,N4111);
and and2374(N4107,N4112,N4113);
and and2375(N4108,R1,N4114);
and and2376(N4109,R3,N4115);
and and2381(N4119,N4123,N4124);
and and2382(N4120,N4125,N4126);
and and2383(N4121,R2,N4127);
and and2384(N4122,R4,R5);
and and2389(N4132,N4136,in0);
and and2390(N4133,N4137,N4138);
and and2391(N4134,R2,N4139);
and and2392(N4135,N4140,R5);
and and2397(N4145,N4149,N4150);
and and2398(N4146,in2,N4151);
and and2399(N4147,R2,N4152);
and and2400(N4148,N4153,R5);
and and2405(N4158,N4162,in0);
and and2406(N4159,R0,N4163);
and and2407(N4160,N4164,N4165);
and and2408(N4161,R4,N4166);
and and2413(N4171,N4175,in0);
and and2414(N4172,N4176,R0);
and and2415(N4173,N4177,N4178);
and and2416(N4174,R4,N4179);
and and2421(N4184,N4188,in0);
and and2422(N4185,N4189,N4190);
and and2423(N4186,N4191,R3);
and and2424(N4187,R4,N4192);
and and2429(N4197,N4201,in1);
and and2430(N4198,N4202,N4203);
and and2431(N4199,N4204,R3);
and and2432(N4200,R4,N4205);
and and2437(N4210,N4214,in0);
and and2438(N4211,N4215,N4216);
and and2439(N4212,N4217,R3);
and and2440(N4213,R4,N4218);
and and2445(N4223,N4227,N4228);
and and2446(N4224,N4229,N4230);
and and2447(N4225,R0,R2);
and and2448(N4226,R3,R5);
and and2453(N4236,N4240,N4241);
and and2454(N4237,in1,in2);
and and2455(N4238,N4242,R1);
and and2456(N4239,N4243,R4);
and and2461(N4249,N4253,in0);
and and2462(N4250,N4254,R0);
and and2463(N4251,N4255,R3);
and and2464(N4252,R4,N4256);
and and2469(N4262,N4266,N4267);
and and2470(N4263,in1,N4268);
and and2471(N4264,N4269,R3);
and and2472(N4265,N4270,R5);
and and2477(N4275,N4279,N4280);
and and2478(N4276,N4281,R0);
and and2479(N4277,R1,N4282);
and and2480(N4278,N4283,N4284);
and and2485(N4288,N4292,in0);
and and2486(N4289,in1,in2);
and and2487(N4290,N4293,N4294);
and and2488(N4291,N4295,R3);
and and2493(N4301,N4305,in0);
and and2494(N4302,N4306,N4307);
and and2495(N4303,N4308,R2);
and and2496(N4304,R3,N4309);
and and2501(N4314,N4318,in0);
and and2502(N4315,N4319,N4320);
and and2503(N4316,R0,N4321);
and and2504(N4317,R2,N4322);
and and2509(N4327,N4331,N4332);
and and2510(N4328,in1,N4333);
and and2511(N4329,N4334,R2);
and and2512(N4330,N4335,R4);
and and2517(N4340,N4344,N4345);
and and2518(N4341,N4346,R0);
and and2519(N4342,N4347,R3);
and and2520(N4343,R4,N4348);
and and2525(N4353,N4357,N4358);
and and2526(N4354,in1,R0);
and and2527(N4355,R1,R3);
and and2528(N4356,N4359,N4360);
and and2533(N4366,N4370,in0);
and and2534(N4367,in2,N4371);
and and2535(N4368,R2,R3);
and and2536(N4369,N4372,N4373);
and and2541(N4379,N4383,in0);
and and2542(N4380,N4384,N4385);
and and2543(N4381,R2,N4386);
and and2544(N4382,N4387,R5);
and and2549(N4392,N4396,in0);
and and2550(N4393,N4397,R0);
and and2551(N4394,N4398,R3);
and and2552(N4395,R4,N4399);
and and2557(N4405,N4409,N4410);
and and2558(N4406,in1,N4411);
and and2559(N4407,N4412,R3);
and and2560(N4408,R4,N4413);
and and2565(N4418,N4422,in0);
and and2566(N4419,N4423,N4424);
and and2567(N4420,R1,N4425);
and and2568(N4421,N4426,R4);
and and2573(N4431,N4435,in0);
and and2574(N4432,N4436,N4437);
and and2575(N4433,R1,R2);
and and2576(N4434,N4438,N4439);
and and2581(N4444,N4448,N4449);
and and2582(N4445,in1,N4450);
and and2583(N4446,R0,R1);
and and2584(N4447,R3,N4451);
and and2589(N4457,N4461,in0);
and and2590(N4458,N4462,R0);
and and2591(N4459,N4463,R2);
and and2592(N4460,N4464,N4465);
and and2597(N4470,N4474,N4475);
and and2598(N4471,in1,in2);
and and2599(N4472,R0,R1);
and and2600(N4473,N4476,N4477);
and and2605(N4483,N4487,in0);
and and2606(N4484,N4488,N4489);
and and2607(N4485,R1,R2);
and and2608(N4486,N4490,N4491);
and and2613(N4496,N4500,in1);
and and2614(N4497,in2,R0);
and and2615(N4498,N4501,R3);
and and2616(N4499,N4502,R5);
and and2621(N4508,N4512,N4513);
and and2622(N4509,in2,R0);
and and2623(N4510,N4514,R3);
and and2624(N4511,R4,N4515);
and and2629(N4520,N4524,in0);
and and2630(N4521,in2,N4525);
and and2631(N4522,R1,R3);
and and2632(N4523,N4526,R5);
and and2637(N4532,N4536,in0);
and and2638(N4533,in1,N4537);
and and2639(N4534,R1,N4538);
and and2640(N4535,R3,N4539);
and and2645(N4544,N4548,N4549);
and and2646(N4545,in2,R0);
and and2647(N4546,R1,N4550);
and and2648(N4547,R4,N4551);
and and2653(N4556,N4560,in0);
and and2654(N4557,N4561,R1);
and and2655(N4558,N4562,R3);
and and2656(N4559,N4563,R5);
and and2661(N4568,N4572,in0);
and and2662(N4569,in1,in2);
and and2663(N4570,N4573,N4574);
and and2664(N4571,R2,N4575);
and and2669(N4580,N4584,N4585);
and and2670(N4581,in1,N4586);
and and2671(N4582,R1,R2);
and and2672(N4583,R3,N4587);
and and2677(N4592,N4596,N4597);
and and2678(N4593,R0,N4598);
and and2679(N4594,N4599,R3);
and and2680(N4595,R4,R5);
and and2685(N4604,N4608,in0);
and and2686(N4605,in2,N4609);
and and2687(N4606,R2,R3);
and and2688(N4607,N4610,R5);
and and2693(N4616,N4620,in0);
and and2694(N4617,in1,N4621);
and and2695(N4618,N4622,R2);
and and2696(N4619,R3,N4623);
and and2701(N4628,N4632,in0);
and and2702(N4629,N4633,N4634);
and and2703(N4630,N4635,R2);
and and2704(N4631,R3,R5);
and and2709(N4640,N4644,in0);
and and2710(N4641,N4645,R0);
and and2711(N4642,R1,N4646);
and and2712(N4643,N4647,R5);
and and2717(N4652,N4656,in1);
and and2718(N4653,N4657,R0);
and and2719(N4654,R1,N4658);
and and2720(N4655,N4659,R5);
and and2725(N4664,N4668,N4669);
and and2726(N4665,R0,R1);
and and2727(N4666,R2,R3);
and and2728(N4667,N4670,N4671);
and and2733(N4676,N4680,in0);
and and2734(N4677,N4681,R1);
and and2735(N4678,N4682,N4683);
and and2736(N4679,R4,R5);
and and2741(N4688,N4692,in0);
and and2742(N4689,in1,N4693);
and and2743(N4690,N4694,R3);
and and2744(N4691,N4695,R5);
and and2749(N4700,N4704,in0);
and and2750(N4701,N4705,R0);
and and2751(N4702,R2,N4706);
and and2752(N4703,N4707,N4708);
and and2757(N4712,N4716,in0);
and and2758(N4713,in1,N4717);
and and2759(N4714,R0,N4718);
and and2760(N4715,R4,N4719);
and and2765(N4724,N4728,N4729);
and and2766(N4725,N4730,in2);
and and2767(N4726,R0,R1);
and and2768(N4727,N4731,R4);
and and2773(N4736,N4740,in1);
and and2774(N4737,in2,N4741);
and and2775(N4738,R1,R2);
and and2776(N4739,N4742,N4743);
and and2781(N4748,N4752,in0);
and and2782(N4749,in1,in2);
and and2783(N4750,N4753,R1);
and and2784(N4751,N4754,N4755);
and and2789(N4760,N4764,in0);
and and2790(N4761,N4765,R0);
and and2791(N4762,N4766,R2);
and and2792(N4763,R3,N4767);
and and2797(N4772,N4776,N4777);
and and2798(N4773,in1,R0);
and and2799(N4774,N4778,R2);
and and2800(N4775,N4779,R4);
and and2805(N4784,N4788,N4789);
and and2806(N4785,in1,N4790);
and and2807(N4786,R0,R2);
and and2808(N4787,R4,R5);
and and2813(N4796,N4800,in0);
and and2814(N4797,N4801,R0);
and and2815(N4798,N4802,R3);
and and2816(N4799,R4,R5);
and and2821(N4808,N4812,in0);
and and2822(N4809,in2,R0);
and and2823(N4810,R1,N4813);
and and2824(N4811,R4,N4814);
and and2829(N4820,N4824,N4825);
and and2830(N4821,N4826,in2);
and and2831(N4822,R0,N4827);
and and2832(N4823,R3,R4);
and and2837(N4832,N4836,N4837);
and and2838(N4833,N4838,R0);
and and2839(N4834,R1,R2);
and and2840(N4835,R3,N4839);
and and2845(N4844,N4848,in0);
and and2846(N4845,in1,R0);
and and2847(N4846,N4849,N4850);
and and2848(N4847,R4,N4851);
and and2853(N4856,N4860,N4861);
and and2854(N4857,N4862,R1);
and and2855(N4858,N4863,R3);
and and2856(N4859,N4864,R5);
and and2861(N4868,N4872,N4873);
and and2862(N4869,N4874,R1);
and and2863(N4870,N4875,R3);
and and2864(N4871,N4876,R5);
and and2869(N4880,N4884,in0);
and and2870(N4881,R0,R1);
and and2871(N4882,N4885,N4886);
and and2872(N4883,R4,N4887);
and and2877(N4892,N4896,N4897);
and and2878(N4893,N4898,N4899);
and and2879(N4894,R0,R1);
and and2880(N4895,R3,N4900);
and and2885(N4904,N4908,in1);
and and2886(N4905,in2,R0);
and and2887(N4906,N4909,R3);
and and2888(N4907,N4910,R5);
and and2893(N4916,N4920,N4921);
and and2894(N4917,in1,in2);
and and2895(N4918,N4922,R1);
and and2896(N4919,R2,N4923);
and and2901(N4928,N4932,in0);
and and2902(N4929,N4933,R0);
and and2903(N4930,N4934,R3);
and and2904(N4931,R4,R5);
and and2909(N4940,N4944,in0);
and and2910(N4941,N4945,R0);
and and2911(N4942,R1,N4946);
and and2912(N4943,N4947,R4);
and and2917(N4952,N4956,in0);
and and2918(N4953,N4957,N4958);
and and2919(N4954,N4959,R2);
and and2920(N4955,R3,R5);
and and2925(N4964,N4968,N4969);
and and2926(N4965,in1,in2);
and and2927(N4966,N4970,N4971);
and and2928(N4967,R2,R4);
and and2933(N4976,N4980,in1);
and and2934(N4977,R0,R1);
and and2935(N4978,R2,R3);
and and2936(N4979,R4,N4981);
and and2941(N4987,N4991,in0);
and and2942(N4988,N4992,R0);
and and2943(N4989,R1,R2);
and and2944(N4990,R3,R4);
and and2949(N4998,N5002,in0);
and and2950(N4999,in1,in2);
and and2951(N5000,N5003,R1);
and and2952(N5001,R3,R4);
and and2957(N5009,N5013,N5014);
and and2958(N5010,in1,in2);
and and2959(N5011,R0,R1);
and and2960(N5012,N5015,R3);
and and2965(N5020,N5024,in0);
and and2966(N5021,N5025,R0);
and and2967(N5022,R1,N5026);
and and2968(N5023,R3,R5);
and and2973(N5031,N5035,in0);
and and2974(N5032,N5036,N5037);
and and2975(N5033,R2,R3);
and and2976(N5034,R4,N5038);
and and2981(N5042,N5046,N5047);
and and2982(N5043,R0,R1);
and and2983(N5044,R2,R3);
and and2984(N5045,N5048,R5);
and and2989(N5053,N5057,in0);
and and2990(N5054,R0,R1);
and and2991(N5055,N5058,R3);
and and2992(N5056,R4,N5059);
and and2997(N5064,N5068,N5069);
and and2998(N5065,in2,N5070);
and and2999(N5066,N5071,R2);
and and3000(N5067,R3,R4);
and and3005(N5075,N5079,in0);
and and3006(N5076,R0,N5080);
and and3007(N5077,N5081,R3);
and and3008(N5078,R4,R5);
and and3013(N5086,N5090,in0);
and and3014(N5087,in1,N5091);
and and3015(N5088,R1,R2);
and and3016(N5089,R3,N5092);
and and3021(N5097,N5101,in0);
and and3022(N5098,N5102,R1);
and and3023(N5099,R2,R3);
and and3024(N5100,R4,R5);
and and3029(N5108,N5112,in0);
and and3030(N5109,in1,R0);
and and3031(N5110,N5113,R2);
and and3032(N5111,N5114,R5);
and and3037(N5119,N5123,in0);
and and3038(N5120,in1,N5124);
and and3039(N5121,R0,R3);
and and3040(N5122,N5125,N5126);
and and3045(N5130,N5134,in0);
and and3046(N5131,in2,N5135);
and and3047(N5132,R2,N5136);
and and3048(N5133,R4,R5);
and and3053(N5141,N5145,N5146);
and and3054(N5142,in2,R1);
and and3055(N5143,R2,N5147);
and and3056(N5144,R4,R5);
and and3061(N5152,N5156,in1);
and and3062(N5153,N5157,R0);
and and3063(N5154,R1,R3);
and and3064(N5155,N5158,N5159);
and and3069(N5163,N5167,in0);
and and3070(N5164,R0,N5168);
and and3071(N5165,N5169,R3);
and and3072(N5166,R4,R5);
and and3077(N5174,N5178,N5179);
and and3078(N5175,N5180,in2);
and and3079(N5176,R0,R1);
and and3080(N5177,R4,N5181);
and and3085(N5185,N5189,in0);
and and3086(N5186,in1,R0);
and and3087(N5187,R1,R2);
and and3088(N5188,N5190,R5);
and and3093(N5195,N5199,in0);
and and3094(N5196,in1,N5200);
and and3095(N5197,N5201,R2);
and and3096(N5198,R3,R4);
and and3101(N5205,N5209,in0);
and and3102(N5206,in1,in2);
and and3103(N5207,R1,R2);
and and3104(N5208,N5210,R5);
and and3109(N5215,N5219,in0);
and and3110(N5216,N5220,N5221);
and and3111(N5217,R2,R3);
and and3112(N5218,R4,R5);
and and3117(N5225,N5229,in0);
and and3118(N5226,N5230,R0);
and and3119(N5227,R2,R3);
and and3120(N5228,N5231,R5);
and and3125(N5235,N5239,in0);
and and3126(N5236,in1,R0);
and and3127(N5237,R1,R2);
and and3128(N5238,R3,R4);
and and3133(N5245,N5249,in0);
and and3134(N5246,in2,R0);
and and3135(N5247,R1,R3);
and and3136(N5248,N5250,N5251);
and and3141(N5255,N5259,in0);
and and3142(N5256,in1,in2);
and and3143(N5257,R0,R2);
and and3144(N5258,R3,N5260);
and and3149(N5264,N5268,in0);
and and3150(N5265,N5269,in2);
and and3151(N5266,R0,R2);
and and3152(N5267,R3,R5);
and and3157(N5273,N5277,in0);
and and3158(N5274,in1,N5278);
and and3159(N5275,R2,R3);
and and3160(N5276,R4,R5);
and and3165(N5282,in0,N5286);
and and3166(N5283,N5287,N5288);
and and3167(N5284,N5289,N5290);
and and3168(N5285,N5291,N5292);
and and3172(N5296,in0,N5300);
and and3173(N5297,N5301,N5302);
and and3174(N5298,N5303,N5304);
and and3175(N5299,N5305,R7);
and and3179(N5309,N5313,N5314);
and and3180(N5310,R0,N5315);
and and3181(N5311,N5316,N5317);
and and3182(N5312,R6,N5318);
and and3186(N5322,in0,N5326);
and and3187(N5323,N5327,R1);
and and3188(N5324,N5328,N5329);
and and3189(N5325,N5330,R6);
and and3193(N5334,in1,R0);
and and3194(N5335,R1,N5338);
and and3195(N5336,N5339,N5340);
and and3196(N5337,N5341,N5342);
and and3200(N5346,in0,N5350);
and and3201(N5347,R1,N5351);
and and3202(N5348,N5352,R5);
and and3203(N5349,N5353,N5354);
and and3207(N5358,in0,N5362);
and and3208(N5359,N5363,R1);
and and3209(N5360,N5364,N5365);
and and3210(N5361,N5366,R6);
and and3214(N5370,in0,R0);
and and3215(N5371,R1,N5374);
and and3216(N5372,N5375,N5376);
and and3217(N5373,R5,N5377);
and and3221(N5381,in0,in2);
and and3222(N5382,R0,N5385);
and and3223(N5383,N5386,N5387);
and and3224(N5384,R6,N5388);
and and3228(N5392,N5396,R0);
and and3229(N5393,N5397,R3);
and and3230(N5394,N5398,N5399);
and and3231(N5395,R6,R7);
and and3235(N5403,N5407,N5408);
and and3236(N5404,R1,R3);
and and3237(N5405,R4,N5409);
and and3238(N5406,N5410,R7);
and and3242(N5414,in0,N5418);
and and3243(N5415,R1,R2);
and and3244(N5416,N5419,N5420);
and and3245(N5417,N5421,R6);
and and3249(N5425,in0,N5429);
and and3250(N5426,R1,R2);
and and3251(N5427,N5430,R5);
and and3252(N5428,R6,N5431);
and and3256(N5435,in0,N5439);
and and3257(N5436,R0,R1);
and and3258(N5437,N5440,R4);
and and3259(N5438,R5,N5441);
and and3263(N5445,in0,N5449);
and and3264(N5446,R1,R3);
and and3265(N5447,R4,N5450);
and and3266(N5448,N5451,R7);
and and3270(N5455,in0,N5459);
and and3271(N5456,R0,R3);
and and3272(N5457,N5460,N5461);
and and3273(N5458,R6,R7);
and and3277(N5465,in0,N5469);
and and3278(N5466,R1,R2);
and and3279(N5467,N5470,R4);
and and3280(N5468,R6,R7);
and and3284(N5474,in1,in2);
and and3285(N5475,R1,R3);
and and3286(N5476,N5478,R5);
and and3287(N5477,R6,N5479);
and and3291(N5483,in2,R1);
and and3292(N5484,R2,R3);
and and3293(N5485,N5487,R5);
and and3294(N5486,R6,N5488);
and and3298(N5492,in0,R0);
and and3299(N5493,R1,N5496);
and and3300(N5494,R3,R4);
and and3301(N5495,R5,R6);
and and7(N395,N401,N402);
and and8(N396,N403,N404);
and and16(N412,N419,N420);
and and17(N413,R6,N421);
and and25(N429,R4,N437);
and and26(N430,R6,N438);
and and34(N446,N453,R5);
and and35(N447,N454,N455);
and and43(N463,N470,N471);
and and44(N464,N472,R7);
and and52(N480,R4,N487);
and and53(N481,N488,R7);
and and61(N496,R4,R5);
and and62(N497,N503,N504);
and and70(N512,N518,R5);
and and71(N513,N519,N520);
and and79(N528,N534,N535);
and and80(N529,N536,R7);
and and88(N544,R4,N550);
and and89(N545,N551,N552);
and and97(N560,N565,N566);
and and98(N561,N567,N568);
and and106(N576,N582,N583);
and and107(N577,N584,R7);
and and115(N592,N598,R5);
and and116(N593,N599,N600);
and and124(N608,N614,R5);
and and125(N609,N615,N616);
and and133(N624,N629,N630);
and and134(N625,N631,N632);
and and142(N640,N647,N648);
and and143(N641,R6,R7);
and and151(N656,R4,N663);
and and152(N657,R6,N664);
and and160(N672,R4,N679);
and and161(N673,R6,N680);
and and169(N688,N693,N694);
and and170(N689,N695,N696);
and and178(N704,R4,R5);
and and179(N705,N711,N712);
and and187(N720,N726,R5);
and and188(N721,N727,N728);
and and196(N736,N743,R4);
and and197(N737,N744,R7);
and and205(N752,N757,N758);
and and206(N753,N759,N760);
and and214(N768,R4,N775);
and and215(N769,R6,N776);
and and223(N784,N789,N790);
and and224(N785,N791,N792);
and and232(N800,N806,N807);
and and233(N801,N808,R7);
and and241(N816,R4,N821);
and and242(N817,N822,N823);
and and250(N831,R4,N836);
and and251(N832,N837,N838);
and and259(N846,N852,R5);
and and260(N847,N853,R7);
and and268(N861,R4,R5);
and and269(N862,N867,N868);
and and277(N876,N882,R4);
and and278(N877,R5,N883);
and and286(N891,R4,N897);
and and287(N892,R6,N898);
and and295(N906,N911,N912);
and and296(N907,R6,N913);
and and304(N921,R3,N927);
and and305(N922,R6,N928);
and and313(N936,R4,R5);
and and314(N937,N942,N943);
and and322(N951,R3,N957);
and and323(N952,N958,R6);
and and331(N966,N972,N973);
and and332(N967,R6,R7);
and and340(N981,N986,N987);
and and341(N982,R6,N988);
and and349(N996,R4,N1002);
and and350(N997,R6,N1003);
and and358(N1011,N1016,N1017);
and and359(N1012,R6,N1018);
and and367(N1026,N1031,N1032);
and and368(N1027,N1033,R7);
and and376(N1041,N1046,N1047);
and and377(N1042,N1048,R7);
and and385(N1056,R3,N1062);
and and386(N1057,N1063,R7);
and and394(N1071,N1077,R5);
and and395(N1072,R6,N1078);
and and403(N1086,N1092,N1093);
and and404(N1087,R6,R7);
and and412(N1101,N1106,N1107);
and and413(N1102,R6,N1108);
and and421(N1116,N1122,R5);
and and422(N1117,R6,N1123);
and and430(N1131,N1137,R5);
and and431(N1132,N1138,R7);
and and439(N1146,N1151,N1152);
and and440(N1147,R6,N1153);
and and448(N1161,N1165,N1166);
and and449(N1162,N1167,N1168);
and and457(N1176,N1182,R5);
and and458(N1177,R6,N1183);
and and466(N1191,N1197,R5);
and and467(N1192,R6,N1198);
and and475(N1206,N1211,R5);
and and476(N1207,N1212,N1213);
and and484(N1221,N1226,R5);
and and485(N1222,N1227,N1228);
and and493(N1236,R3,R4);
and and494(N1237,N1242,N1243);
and and502(N1251,N1256,N1257);
and and503(N1252,N1258,R7);
and and511(N1266,R4,R5);
and and512(N1267,N1273,R7);
and and520(N1281,N1286,R4);
and and521(N1282,N1287,N1288);
and and529(N1296,N1301,N1302);
and and530(N1297,N1303,R7);
and and538(N1311,N1316,R5);
and and539(N1312,N1317,N1318);
and and547(N1326,N1331,R5);
and and548(N1327,N1332,N1333);
and and556(N1341,R4,N1347);
and and557(N1342,R6,N1348);
and and565(N1356,R4,N1362);
and and566(N1357,R6,N1363);
and and574(N1371,N1376,R5);
and and575(N1372,N1377,N1378);
and and583(N1386,N1392,R4);
and and584(N1387,N1393,R7);
and and592(N1401,N1406,R5);
and and593(N1402,N1407,N1408);
and and601(N1416,R4,N1422);
and and602(N1417,N1423,R7);
and and610(N1431,N1436,N1437);
and and611(N1432,R6,R7);
and and619(N1445,R3,N1451);
and and620(N1446,R6,R7);
and and628(N1459,R4,N1463);
and and629(N1460,N1464,N1465);
and and637(N1473,R3,N1477);
and and638(N1474,N1478,N1479);
and and646(N1487,N1490,N1491);
and and647(N1488,N1492,N1493);
and and655(N1501,R4,N1507);
and and656(N1502,R6,R7);
and and664(N1515,R4,N1520);
and and665(N1516,R6,N1521);
and and673(N1529,N1533,N1534);
and and674(N1530,N1535,R7);
and and682(N1543,N1547,N1548);
and and683(N1544,R6,N1549);
and and691(N1557,N1560,N1561);
and and692(N1558,N1562,N1563);
and and700(N1571,N1574,N1575);
and and701(N1572,N1576,N1577);
and and709(N1585,R4,N1589);
and and710(N1586,N1590,N1591);
and and718(N1599,N1603,R5);
and and719(N1600,N1604,N1605);
and and727(N1613,R4,N1619);
and and728(N1614,R6,R7);
and and736(N1627,N1632,R5);
and and737(N1628,R6,N1633);
and and745(N1641,N1645,R5);
and and746(N1642,N1646,N1647);
and and754(N1655,R3,N1660);
and and755(N1656,R5,N1661);
and and763(N1669,N1673,N1674);
and and764(N1670,R6,N1675);
and and772(N1683,N1688,R5);
and and773(N1684,N1689,R7);
and and781(N1697,N1702,R5);
and and782(N1698,R6,N1703);
and and790(N1711,N1716,N1717);
and and791(N1712,R6,R7);
and and799(N1725,N1730,N1731);
and and800(N1726,R6,R7);
and and808(N1739,N1744,N1745);
and and809(N1740,R6,R7);
and and817(N1753,R3,N1759);
and and818(N1754,R6,R7);
and and826(N1767,R4,R5);
and and827(N1768,N1772,N1773);
and and835(N1781,N1786,R5);
and and836(N1782,N1787,R7);
and and844(N1795,N1800,R5);
and and845(N1796,N1801,R7);
and and853(N1809,R4,R5);
and and854(N1810,R6,N1815);
and and862(N1823,R4,N1828);
and and863(N1824,R6,N1829);
and and871(N1837,R3,R4);
and and872(N1838,N1843,R6);
and and880(N1851,N1854,N1855);
and and881(N1852,N1856,N1857);
and and889(N1865,R4,N1871);
and and890(N1866,R6,R7);
and and898(N1879,N1883,N1884);
and and899(N1880,N1885,R7);
and and907(N1893,N1898,R4);
and and908(N1894,R6,N1899);
and and916(N1907,R4,N1912);
and and917(N1908,R6,N1913);
and and925(N1921,R4,N1927);
and and926(N1922,R6,R7);
and and934(N1935,R4,R5);
and and935(N1936,R6,N1941);
and and943(N1949,R4,R5);
and and944(N1950,N1955,R7);
and and952(N1963,R4,N1969);
and and953(N1964,R6,R7);
and and961(N1977,R3,R4);
and and962(N1978,R5,R6);
and and970(N1991,N1995,N1996);
and and971(N1992,N1997,R7);
and and979(N2005,N2009,N2010);
and and980(N2006,N2011,R7);
and and988(N2019,N2023,N2024);
and and989(N2020,N2025,R7);
and and997(N2033,R3,N2038);
and and998(N2034,R5,N2039);
and and1006(N2047,R4,N2052);
and and1007(N2048,N2053,R7);
and and1015(N2061,N2065,N2066);
and and1016(N2062,N2067,R7);
and and1024(N2075,R3,R4);
and and1025(N2076,N2081,R6);
and and1033(N2089,N2093,R5);
and and1034(N2090,N2094,N2095);
and and1042(N2103,R4,R5);
and and1043(N2104,N2108,N2109);
and and1051(N2117,N2119,N2120);
and and1052(N2118,N2121,N2122);
and and1060(N2130,R3,N2133);
and and1061(N2131,N2134,N2135);
and and1069(N2143,R4,N2146);
and and1070(N2144,N2147,N2148);
and and1078(N2156,N2160,R5);
and and1079(N2157,N2161,R7);
and and1087(N2169,R4,R5);
and and1088(N2170,N2174,R7);
and and1096(N2182,R4,N2186);
and and1097(N2183,R6,N2187);
and and1105(N2195,R3,N2199);
and and1106(N2196,N2200,R6);
and and1114(N2208,R3,N2212);
and and1115(N2209,N2213,R7);
and and1123(N2221,N2225,R5);
and and1124(N2222,N2226,R7);
and and1132(N2234,R4,N2238);
and and1133(N2235,R6,N2239);
and and1141(N2247,N2250,N2251);
and and1142(N2248,R6,N2252);
and and1150(N2260,R4,R5);
and and1151(N2261,R6,N2265);
and and1159(N2273,R4,R5);
and and1160(N2274,N2278,R7);
and and1168(N2286,R3,N2290);
and and1169(N2287,N2291,R7);
and and1177(N2299,N2302,N2303);
and and1178(N2300,N2304,R7);
and and1186(N2312,R4,R5);
and and1187(N2313,N2316,N2317);
and and1195(N2325,R3,N2329);
and and1196(N2326,R6,N2330);
and and1204(N2338,R4,R5);
and and1205(N2339,R6,N2343);
and and1213(N2351,R3,R4);
and and1214(N2352,R5,N2356);
and and1222(N2364,N2368,R5);
and and1223(N2365,N2369,R7);
and and1231(N2377,R4,R5);
and and1232(N2378,N2382,R7);
and and1240(N2390,R3,N2394);
and and1241(N2391,R5,N2395);
and and1249(N2403,R3,R4);
and and1250(N2404,N2407,N2408);
and and1258(N2416,R4,N2420);
and and1259(N2417,R6,N2421);
and and1267(N2429,R4,N2433);
and and1268(N2430,R6,N2434);
and and1276(N2442,R4,N2446);
and and1277(N2443,R6,N2447);
and and1285(N2455,R4,N2459);
and and1286(N2456,R6,N2460);
and and1294(N2468,R4,R5);
and and1295(N2469,N2473,R7);
and and1303(N2481,R4,R5);
and and1304(N2482,N2486,R7);
and and1312(N2494,R3,N2498);
and and1313(N2495,N2499,R7);
and and1321(N2507,N2512,R4);
and and1322(N2508,R5,R7);
and and1330(N2520,R3,R5);
and and1331(N2521,N2524,N2525);
and and1339(N2533,N2536,N2537);
and and1340(N2534,N2538,R7);
and and1348(N2546,R3,R4);
and and1349(N2547,R5,N2551);
and and1357(N2559,R3,R4);
and and1358(N2560,R5,N2564);
and and1366(N2572,N2577,R4);
and and1367(N2573,R6,R7);
and and1375(N2585,R4,N2589);
and and1376(N2586,N2590,R7);
and and1384(N2598,N2603,R5);
and and1385(N2599,R6,R7);
and and1393(N2611,N2614,R5);
and and1394(N2612,N2615,R7);
and and1402(N2623,R3,N2627);
and and1403(N2624,R6,R7);
and and1411(N2635,N2638,N2639);
and and1412(N2636,R6,R7);
and and1420(N2647,N2650,R5);
and and1421(N2648,R6,N2651);
and and1429(N2659,N2662,N2663);
and and1430(N2660,R6,R7);
and and1438(N2671,R4,N2674);
and and1439(N2672,N2675,R7);
and and1447(N2683,R4,R5);
and and1448(N2684,N2687,R7);
and and1456(N2695,R4,R5);
and and1457(N2696,N2699,R7);
and and1465(N2707,N2710,R5);
and and1466(N2708,N2711,R7);
and and1474(N2719,R4,R5);
and and1475(N2720,R6,N2723);
and and1483(N2731,R4,R5);
and and1484(N2732,N2735,R7);
and and1492(N2743,R4,N2747);
and and1493(N2744,R6,R7);
and and1501(N2755,R4,N2759);
and and1502(N2756,R6,R7);
and and1510(N2767,R3,R5);
and and1511(N2768,R6,N2771);
and and1519(N2779,R3,R4);
and and1520(N2780,N2783,R7);
and and1528(N2791,R3,N2794);
and and1529(N2792,N2795,R7);
and and1537(N2803,N2806,R5);
and and1538(N2804,N2807,R7);
and and1546(N2815,N2818,N2819);
and and1547(N2816,R6,R7);
and and1555(N2827,R3,R4);
and and1556(N2828,R5,N2831);
and and1564(N2839,R3,R5);
and and1565(N2840,N2843,R7);
and and1573(N2851,R3,R5);
and and1574(N2852,R6,R7);
and and1582(N2863,R4,R5);
and and1583(N2864,R6,N2867);
and and1591(N2875,N2878,R4);
and and1592(N2876,R6,N2879);
and and1600(N2887,R3,R4);
and and1601(N2888,R5,R6);
and and1609(N2899,R3,R4);
and and1610(N2900,R5,R7);
and and1618(N2911,R3,N2914);
and and1619(N2912,N2915,R7);
and and1627(N2923,R3,R5);
and and1628(N2924,R6,R7);
and and1636(N2935,R4,N2939);
and and1637(N2936,R6,R7);
and and1645(N2947,R4,R5);
and and1646(N2948,R6,N2951);
and and1654(N2959,N2963,R5);
and and1655(N2960,R6,R7);
and and1663(N2971,N2975,R5);
and and1664(N2972,R6,R7);
and and1672(N2983,R4,R5);
and and1673(N2984,R6,N2987);
and and1681(N2995,R4,R5);
and and1682(N2996,R6,R7);
and and1690(N3007,R3,N3011);
and and1691(N3008,R6,R7);
and and1699(N3019,N3021,N3022);
and and1700(N3020,N3023,R7);
and and1708(N3031,R4,R5);
and and1709(N3032,N3035,R7);
and and1717(N3043,R4,R5);
and and1718(N3044,N3046,N3047);
and and1726(N3055,R4,R5);
and and1727(N3056,N3058,N3059);
and and1735(N3067,R4,N3071);
and and1736(N3068,R6,R7);
and and1744(N3079,N3082,N3083);
and and1745(N3080,R5,R7);
and and1753(N3091,R4,R5);
and and1754(N3092,N3094,R7);
and and1762(N3102,N3104,R5);
and and1763(N3103,N3105,R7);
and and1771(N3113,R3,R5);
and and1772(N3114,N3116,R7);
and and1780(N3124,R4,R5);
and and1781(N3125,R6,N3127);
and and1789(N3135,R4,N3137);
and and1790(N3136,R6,N3138);
and and1798(N3146,R4,N3148);
and and1799(N3147,N3149,R7);
and and1807(N3157,R3,N3159);
and and1808(N3158,N3160,R6);
and and1816(N3168,R3,R5);
and and1817(N3169,R6,R7);
and and1825(N3179,R3,R4);
and and1826(N3180,R6,N3182);
and and1834(N3190,R4,R5);
and and1835(N3191,R6,N3193);
and and1843(N3201,R3,R4);
and and1844(N3202,R5,R6);
and and1852(N3212,R3,R4);
and and1853(N3213,R6,R7);
and and1861(N3223,N3225,R5);
and and1862(N3224,N3226,R7);
and and1870(N3234,R4,R5);
and and1871(N3235,R6,R7);
and and1879(N3244,R4,R5);
and and1880(N3245,R6,R7);
and and1888(N3254,R4,R5);
and and1889(N3255,R6,R7);
and and1897(N3263,N3270,N3271);
and and1905(N3279,R6,N3287);
and and1913(N3295,N3302,N3303);
and and1921(N3311,N3318,N3319);
and and1929(N3327,N3334,N3335);
and and1937(N3343,N3350,N3351);
and and1945(N3359,R6,N3367);
and and1953(N3375,N3382,R7);
and and1961(N3390,N3396,N3397);
and and1969(N3405,N3411,N3412);
and and1977(N3420,N3426,N3427);
and and1985(N3435,R6,N3442);
and and1993(N3450,N3456,N3457);
and and2001(N3465,N3471,N3472);
and and2009(N3480,N3486,N3487);
and and2017(N3495,N3502,R7);
and and2025(N3510,N3516,N3517);
and and2033(N3525,R5,N3531);
and and2041(N3539,N3544,N3545);
and and2049(N3553,N3558,N3559);
and and2057(N3567,N3572,N3573);
and and2065(N3581,N3586,N3587);
and and2073(N3595,N3601,R7);
and and2081(N3609,N3614,N3615);
and and2089(N3623,R6,N3629);
and and2097(N3637,N3642,N3643);
and and2105(N3651,R6,N3657);
and and2113(N3665,N3670,N3671);
and and2121(N3679,N3684,N3685);
and and2129(N3693,R6,N3699);
and and2137(N3707,R6,N3713);
and and2145(N3721,N3726,N3727);
and and2153(N3735,R6,N3741);
and and2161(N3749,N3755,R7);
and and2169(N3763,N3768,N3769);
and and2177(N3777,N3782,N3783);
and and2185(N3791,N3797,R7);
and and2193(N3805,R6,N3811);
and and2201(N3819,N3824,N3825);
and and2209(N3833,N3838,N3839);
and and2217(N3847,N3853,R7);
and and2225(N3861,N3867,R7);
and and2233(N3875,R6,N3881);
and and2241(N3889,N3893,N3894);
and and2249(N3902,N3906,N3907);
and and2257(N3915,N3919,N3920);
and and2265(N3928,N3932,N3933);
and and2273(N3941,N3945,N3946);
and and2281(N3954,N3958,N3959);
and and2289(N3967,N3972,R7);
and and2297(N3980,N3984,N3985);
and and2305(N3993,N3998,R6);
and and2313(N4006,R6,N4011);
and and2321(N4019,N4023,N4024);
and and2329(N4032,R5,N4037);
and and2337(N4045,N4049,N4050);
and and2345(N4058,R6,N4063);
and and2353(N4071,N4076,R7);
and and2361(N4084,N4089,R7);
and and2369(N4097,R5,N4102);
and and2377(N4110,R5,R7);
and and2385(N4123,N4128,R7);
and and2393(N4136,N4141,R7);
and and2401(N4149,N4154,R7);
and and2409(N4162,N4167,R7);
and and2417(N4175,R6,N4180);
and and2425(N4188,R6,N4193);
and and2433(N4201,N4206,R7);
and and2441(N4214,N4219,R7);
and and2449(N4227,N4231,N4232);
and and2457(N4240,N4244,N4245);
and and2465(N4253,N4257,N4258);
and and2473(N4266,R6,N4271);
and and2481(N4279,R6,R7);
and and2489(N4292,N4296,N4297);
and and2497(N4305,N4310,R7);
and and2505(N4318,R5,N4323);
and and2513(N4331,N4336,R7);
and and2521(N4344,N4349,R7);
and and2529(N4357,N4361,N4362);
and and2537(N4370,N4374,N4375);
and and2545(N4383,N4388,R7);
and and2553(N4396,N4400,N4401);
and and2561(N4409,N4414,R7);
and and2569(N4422,N4427,R6);
and and2577(N4435,N4440,R7);
and and2585(N4448,N4452,N4453);
and and2593(N4461,R5,N4466);
and and2601(N4474,N4478,N4479);
and and2609(N4487,N4492,R7);
and and2617(N4500,N4503,N4504);
and and2625(N4512,R6,N4516);
and and2633(N4524,N4527,N4528);
and and2641(N4536,R5,N4540);
and and2649(N4548,N4552,R7);
and and2657(N4560,R6,N4564);
and and2665(N4572,N4576,R7);
and and2673(N4584,R6,N4588);
and and2681(N4596,N4600,R7);
and and2689(N4608,N4611,N4612);
and and2697(N4620,R5,N4624);
and and2705(N4632,R6,N4636);
and and2713(N4644,N4648,R7);
and and2721(N4656,N4660,R7);
and and2729(N4668,R6,N4672);
and and2737(N4680,R6,N4684);
and and2745(N4692,N4696,R7);
and and2753(N4704,R6,R7);
and and2761(N4716,R6,N4720);
and and2769(N4728,N4732,R6);
and and2777(N4740,N4744,R6);
and and2785(N4752,N4756,R7);
and and2793(N4764,N4768,R7);
and and2801(N4776,N4780,R7);
and and2809(N4788,N4791,N4792);
and and2817(N4800,N4803,N4804);
and and2825(N4812,N4815,N4816);
and and2833(N4824,N4828,R7);
and and2841(N4836,R6,N4840);
and and2849(N4848,R6,N4852);
and and2857(N4860,R6,R7);
and and2865(N4872,R6,R7);
and and2873(N4884,R6,N4888);
and and2881(N4896,R6,R7);
and and2889(N4908,N4911,N4912);
and and2897(N4920,N4924,R6);
and and2905(N4932,N4935,N4936);
and and2913(N4944,R5,N4948);
and and2921(N4956,R6,N4960);
and and2929(N4968,N4972,R7);
and and2937(N4980,N4982,N4983);
and and2945(N4991,N4993,N4994);
and and2953(N5002,N5004,N5005);
and and2961(N5013,R4,N5016);
and and2969(N5024,N5027,R7);
and and2977(N5035,R6,R7);
and and2985(N5046,N5049,R7);
and and2993(N5057,N5060,R7);
and and3001(N5068,R5,R7);
and and3009(N5079,R6,N5082);
and and3017(N5090,R6,N5093);
and and3025(N5101,N5103,N5104);
and and3033(N5112,N5115,R7);
and and3041(N5123,R6,R7);
and and3049(N5134,N5137,R7);
and and3057(N5145,R6,N5148);
and and3065(N5156,R6,R7);
and and3073(N5167,N5170,R7);
and and3081(N5178,R6,R7);
and and3089(N5189,R6,N5191);
and and3097(N5199,R5,R6);
and and3105(N5209,R6,N5211);
and and3113(N5219,R6,R7);
and and3121(N5229,R6,R7);
and and3129(N5239,N5240,N5241);
and and3137(N5249,R6,R7);
and and3145(N5259,R5,R6);
and and3153(N5268,R6,R7);
and and3161(N5277,R6,R7);
and and3302(N5931,N5932,N5933);
and and3311(N5949,N5950,N5951);
and and3320(N5967,N5968,N5969);
and and3329(N5985,N5986,N5987);
and and3338(N6002,N6003,N6004);
and and3347(N6019,N6020,N6021);
and and3356(N6036,N6037,N6038);
and and3365(N6053,N6054,N6055);
and and3374(N6069,N6070,N6071);
and and3383(N6085,N6086,N6087);
and and3392(N6101,N6102,N6103);
and and3401(N6117,N6118,N6119);
and and3410(N6133,N6134,N6135);
and and3419(N6149,N6150,N6151);
and and3428(N6165,N6166,N6167);
and and3437(N6181,N6182,N6183);
and and3446(N6197,N6198,N6199);
and and3455(N6213,N6214,N6215);
and and3464(N6229,N6230,N6231);
and and3473(N6245,N6246,N6247);
and and3482(N6261,N6262,N6263);
and and3491(N6277,N6278,N6279);
and and3500(N6293,N6294,N6295);
and and3509(N6308,N6309,N6310);
and and3518(N6323,N6324,N6325);
and and3527(N6338,N6339,N6340);
and and3536(N6353,N6354,N6355);
and and3545(N6368,N6369,N6370);
and and3554(N6383,N6384,N6385);
and and3563(N6398,N6399,N6400);
and and3572(N6413,N6414,N6415);
and and3581(N6428,N6429,N6430);
and and3590(N6443,N6444,N6445);
and and3599(N6458,N6459,N6460);
and and3608(N6473,N6474,N6475);
and and3617(N6488,N6489,N6490);
and and3626(N6503,N6504,N6505);
and and3635(N6518,N6519,N6520);
and and3644(N6533,N6534,N6535);
and and3653(N6548,N6549,N6550);
and and3662(N6563,N6564,N6565);
and and3671(N6578,N6579,N6580);
and and3680(N6593,N6594,N6595);
and and3689(N6608,N6609,N6610);
and and3698(N6623,N6624,N6625);
and and3707(N6638,N6639,N6640);
and and3716(N6653,N6654,N6655);
and and3725(N6668,N6669,N6670);
and and3734(N6683,N6684,N6685);
and and3743(N6698,N6699,N6700);
and and3752(N6712,N6713,N6714);
and and3761(N6726,N6727,N6728);
and and3770(N6740,N6741,N6742);
and and3779(N6754,N6755,N6756);
and and3788(N6768,N6769,N6770);
and and3797(N6782,N6783,N6784);
and and3806(N6796,N6797,N6798);
and and3815(N6810,N6811,N6812);
and and3824(N6824,N6825,N6826);
and and3833(N6838,N6839,N6840);
and and3842(N6852,N6853,N6854);
and and3851(N6866,N6867,N6868);
and and3860(N6880,N6881,N6882);
and and3869(N6894,N6895,N6896);
and and3878(N6908,N6909,N6910);
and and3887(N6922,N6923,N6924);
and and3896(N6936,N6937,N6938);
and and3905(N6950,N6951,N6952);
and and3914(N6964,N6965,N6966);
and and3923(N6978,N6979,N6980);
and and3932(N6992,N6993,N6994);
and and3941(N7006,N7007,N7008);
and and3950(N7020,N7021,N7022);
and and3959(N7034,N7035,N7036);
and and3968(N7048,N7049,N7050);
and and3977(N7062,N7063,N7064);
and and3986(N7076,N7077,N7078);
and and3995(N7090,N7091,N7092);
and and4004(N7104,N7105,N7106);
and and4013(N7118,N7119,N7120);
and and4022(N7131,N7132,N7133);
and and4031(N7144,N7145,N7146);
and and4040(N7157,N7158,N7159);
and and4049(N7170,N7171,N7172);
and and4058(N7183,N7184,N7185);
and and4067(N7196,N7197,N7198);
and and4076(N7209,N7210,N7211);
and and4085(N7222,N7223,N7224);
and and4094(N7235,N7236,N7237);
and and4103(N7248,N7249,N7250);
and and4112(N7261,N7262,N7263);
and and4121(N7274,N7275,N7276);
and and4130(N7287,N7288,N7289);
and and4139(N7300,N7301,N7302);
and and4148(N7313,N7314,N7315);
and and4157(N7326,N7327,N7328);
and and4166(N7339,N7340,N7341);
and and4175(N7352,N7353,N7354);
and and4184(N7365,N7366,N7367);
and and4193(N7378,N7379,N7380);
and and4202(N7391,N7392,N7393);
and and4211(N7404,N7405,N7406);
and and4220(N7417,N7418,N7419);
and and4229(N7430,N7431,N7432);
and and4238(N7443,N7444,N7445);
and and4247(N7456,N7457,N7458);
and and4256(N7469,N7470,N7471);
and and4265(N7482,N7483,N7484);
and and4274(N7495,N7496,N7497);
and and4283(N7508,N7509,N7510);
and and4292(N7521,N7522,N7523);
and and4301(N7534,N7535,N7536);
and and4310(N7547,N7548,N7549);
and and4319(N7560,N7561,N7562);
and and4328(N7573,N7574,N7575);
and and4337(N7586,N7587,N7588);
and and4346(N7599,N7600,N7601);
and and4355(N7612,N7613,N7614);
and and4364(N7624,N7625,N7626);
and and4373(N7636,N7637,N7638);
and and4382(N7648,N7649,N7650);
and and4391(N7660,N7661,N7662);
and and4400(N7672,N7673,N7674);
and and4409(N7684,N7685,N7686);
and and4418(N7696,N7697,N7698);
and and4427(N7708,N7709,N7710);
and and4436(N7720,N7721,N7722);
and and4445(N7732,N7733,N7734);
and and4454(N7744,N7745,N7746);
and and4463(N7756,N7757,N7758);
and and4472(N7768,N7769,N7770);
and and4481(N7780,N7781,N7782);
and and4490(N7792,N7793,N7794);
and and4499(N7804,N7805,N7806);
and and4508(N7816,N7817,N7818);
and and4517(N7828,N7829,N7830);
and and4526(N7840,N7841,N7842);
and and4535(N7852,N7853,N7854);
and and4544(N7864,N7865,N7866);
and and4553(N7876,N7877,N7878);
and and4562(N7888,N7889,N7890);
and and4571(N7900,N7901,N7902);
and and4580(N7911,N7912,N7913);
and and4589(N7922,N7923,N7924);
and and4598(N7933,N7934,N7935);
and and4607(N7944,N7945,N7946);
and and4616(N7955,N7956,N7957);
and and4625(N7966,N7967,N7968);
and and4634(N7977,N7978,N7979);
and and4643(N7988,N7989,N7990);
and and4652(N7999,N8000,N8001);
and and4661(N8010,N8011,N8012);
and and4670(N8021,N8022,N8023);
and and4679(N8032,N8033,N8034);
and and4688(N8042,N8043,N8044);
and and4697(N8052,N8053,N8054);
and and4706(N8062,N8063,N8064);
and and4715(N8072,N8073,N8074);
and and4724(N8082,N8083,N8084);
and and4733(N8092,N8093,N8094);
and and4742(N8102,N8103,N8104);
and and4751(N8112,N8113,N8114);
and and4760(N8121,N8122,N8123);
and and4768(N8137,N8138,N8139);
and and4776(N8153,N8154,N8155);
and and4784(N8168,N8169,N8170);
and and4792(N8183,N8184,N8185);
and and4800(N8198,N8199,N8200);
and and4808(N8213,N8214,N8215);
and and4816(N8228,N8229,N8230);
and and4824(N8243,N8244,N8245);
and and4832(N8258,N8259,N8260);
and and4840(N8273,N8274,N8275);
and and4848(N8288,N8289,N8290);
and and4856(N8303,N8304,N8305);
and and4864(N8318,N8319,N8320);
and and4872(N8333,N8334,N8335);
and and4880(N8348,N8349,N8350);
and and4888(N8363,N8364,N8365);
and and4896(N8377,N8378,N8379);
and and4904(N8391,N8392,N8393);
and and4912(N8405,N8406,N8407);
and and4920(N8419,N8420,N8421);
and and4928(N8433,N8434,N8435);
and and4936(N8447,N8448,N8449);
and and4944(N8461,N8462,N8463);
and and4952(N8475,N8476,N8477);
and and4960(N8489,N8490,N8491);
and and4968(N8503,N8504,N8505);
and and4976(N8517,N8518,N8519);
and and4984(N8531,N8532,N8533);
and and4992(N8545,N8546,N8547);
and and5000(N8559,N8560,N8561);
and and5008(N8573,N8574,N8575);
and and5016(N8587,N8588,N8589);
and and5024(N8601,N8602,N8603);
and and5032(N8615,N8616,N8617);
and and5040(N8629,N8630,N8631);
and and5048(N8643,N8644,N8645);
and and5056(N8657,N8658,N8659);
and and5064(N8671,N8672,N8673);
and and5072(N8685,N8686,N8687);
and and5080(N8699,N8700,N8701);
and and5088(N8713,N8714,N8715);
and and5096(N8727,N8728,N8729);
and and5104(N8741,N8742,N8743);
and and5112(N8755,N8756,N8757);
and and5120(N8769,N8770,N8771);
and and5128(N8783,N8784,N8785);
and and5136(N8797,N8798,N8799);
and and5144(N8811,N8812,N8813);
and and5152(N8825,N8826,N8827);
and and5160(N8839,N8840,N8841);
and and5168(N8853,N8854,N8855);
and and5176(N8867,N8868,N8869);
and and5184(N8881,N8882,N8883);
and and5192(N8895,N8896,N8897);
and and5200(N8908,N8909,N8910);
and and5208(N8921,N8922,N8923);
and and5216(N8934,N8935,N8936);
and and5224(N8947,N8948,N8949);
and and5232(N8960,N8961,N8962);
and and5240(N8973,N8974,N8975);
and and5248(N8986,N8987,N8988);
and and5256(N8999,N9000,N9001);
and and5264(N9012,N9013,N9014);
and and5272(N9025,N9026,N9027);
and and5280(N9038,N9039,N9040);
and and5288(N9051,N9052,N9053);
and and5296(N9064,N9065,N9066);
and and5304(N9077,N9078,N9079);
and and5312(N9090,N9091,N9092);
and and5320(N9103,N9104,N9105);
and and5328(N9116,N9117,N9118);
and and5336(N9129,N9130,N9131);
and and5344(N9142,N9143,N9144);
and and5352(N9155,N9156,N9157);
and and5360(N9168,N9169,N9170);
and and5368(N9181,N9182,N9183);
and and5376(N9194,N9195,N9196);
and and5384(N9207,N9208,N9209);
and and5392(N9220,N9221,N9222);
and and5400(N9233,N9234,N9235);
and and5408(N9246,N9247,N9248);
and and5416(N9259,N9260,N9261);
and and5424(N9272,N9273,N9274);
and and5432(N9285,N9286,N9287);
and and5440(N9298,N9299,N9300);
and and5448(N9311,N9312,N9313);
and and5456(N9324,N9325,N9326);
and and5464(N9337,N9338,N9339);
and and5472(N9350,N9351,N9352);
and and5480(N9363,N9364,N9365);
and and5488(N9376,N9377,N9378);
and and5496(N9389,N9390,N9391);
and and5504(N9402,N9403,N9404);
and and5512(N9415,N9416,N9417);
and and5520(N9428,N9429,N9430);
and and5528(N9441,N9442,N9443);
and and5536(N9454,N9455,N9456);
and and5544(N9467,N9468,N9469);
and and5552(N9480,N9481,N9482);
and and5560(N9493,N9494,N9495);
and and5568(N9506,N9507,N9508);
and and5576(N9519,N9520,N9521);
and and5584(N9532,N9533,N9534);
and and5592(N9545,N9546,N9547);
and and5600(N9558,N9559,N9560);
and and5608(N9571,N9572,N9573);
and and5616(N9584,N9585,N9586);
and and5624(N9597,N9598,N9599);
and and5632(N9610,N9611,N9612);
and and5640(N9623,N9624,N9625);
and and5648(N9636,N9637,N9638);
and and5656(N9648,N9649,N9650);
and and5664(N9660,N9661,N9662);
and and5672(N9672,N9673,N9674);
and and5680(N9684,N9685,N9686);
and and5688(N9696,N9697,N9698);
and and5696(N9708,N9709,N9710);
and and5704(N9720,N9721,N9722);
and and5712(N9732,N9733,N9734);
and and5720(N9744,N9745,N9746);
and and5728(N9756,N9757,N9758);
and and5736(N9768,N9769,N9770);
and and5744(N9780,N9781,N9782);
and and5752(N9792,N9793,N9794);
and and5760(N9804,N9805,N9806);
and and5768(N9816,N9817,N9818);
and and5776(N9828,N9829,N9830);
and and5784(N9840,N9841,N9842);
and and5792(N9852,N9853,N9854);
and and5800(N9864,N9865,N9866);
and and5808(N9876,N9877,N9878);
and and5816(N9888,N9889,N9890);
and and5824(N9900,N9901,N9902);
and and5832(N9912,N9913,N9914);
and and5840(N9924,N9925,N9926);
and and5848(N9936,N9937,N9938);
and and5856(N9948,N9949,N9950);
and and5864(N9960,N9961,N9962);
and and5872(N9972,N9973,N9974);
and and5880(N9984,N9985,N9986);
and and5888(N9996,N9997,N9998);
and and5896(N10008,N10009,N10010);
and and5904(N10020,N10021,N10022);
and and5912(N10032,N10033,N10034);
and and5920(N10044,N10045,N10046);
and and5928(N10056,N10057,N10058);
and and5936(N10068,N10069,N10070);
and and5944(N10080,N10081,N10082);
and and5952(N10092,N10093,N10094);
and and5960(N10104,N10105,N10106);
and and5968(N10116,N10117,N10118);
and and5976(N10128,N10129,N10130);
and and5984(N10140,N10141,N10142);
and and5992(N10152,N10153,N10154);
and and6000(N10164,N10165,N10166);
and and6008(N10176,N10177,N10178);
and and6016(N10188,N10189,N10190);
and and6024(N10200,N10201,N10202);
and and6032(N10211,N10212,N10213);
and and6040(N10222,N10223,N10224);
and and6048(N10233,N10234,N10235);
and and6056(N10244,N10245,N10246);
and and6064(N10255,N10256,N10257);
and and6072(N10266,N10267,N10268);
and and6080(N10277,N10278,N10279);
and and6088(N10288,N10289,N10290);
and and6096(N10299,N10300,N10301);
and and6104(N10310,N10311,N10312);
and and6112(N10321,N10322,N10323);
and and6120(N10332,N10333,N10334);
and and6128(N10343,N10344,N10345);
and and6136(N10354,N10355,N10356);
and and6144(N10365,N10366,N10367);
and and6152(N10376,N10377,N10378);
and and6160(N10387,N10388,N10389);
and and6168(N10398,N10399,N10400);
and and6176(N10409,N10410,N10411);
and and6184(N10420,N10421,N10422);
and and6192(N10431,N10432,N10433);
and and6200(N10442,N10443,N10444);
and and6208(N10453,N10454,N10455);
and and6216(N10464,N10465,N10466);
and and6224(N10475,N10476,N10477);
and and6232(N10486,N10487,N10488);
and and6240(N10497,N10498,N10499);
and and6248(N10508,N10509,N10510);
and and6256(N10519,N10520,N10521);
and and6264(N10530,N10531,N10532);
and and6272(N10541,N10542,N10543);
and and6280(N10552,N10553,N10554);
and and6288(N10563,N10564,N10565);
and and6296(N10574,N10575,N10576);
and and6304(N10585,N10586,N10587);
and and6312(N10596,N10597,N10598);
and and6320(N10607,N10608,N10609);
and and6328(N10618,N10619,N10620);
and and6336(N10629,N10630,N10631);
and and6344(N10640,N10641,N10642);
and and6352(N10651,N10652,N10653);
and and6360(N10662,N10663,N10664);
and and6368(N10673,N10674,N10675);
and and6376(N10683,N10684,N10685);
and and6384(N10693,N10694,N10695);
and and6392(N10703,N10704,N10705);
and and6400(N10713,N10714,N10715);
and and6408(N10723,N10724,N10725);
and and6416(N10733,N10734,N10735);
and and6424(N10743,N10744,N10745);
and and6432(N10753,N10754,N10755);
and and6440(N10763,N10764,N10765);
and and6448(N10773,N10774,N10775);
and and6456(N10783,N10784,N10785);
and and6464(N10793,N10794,N10795);
and and6472(N10803,N10804,N10805);
and and6480(N10813,N10814,N10815);
and and6488(N10823,N10824,N10825);
and and6496(N10833,N10834,N10835);
and and6504(N10843,N10844,N10845);
and and6512(N10853,N10854,N10855);
and and6520(N10863,N10864,N10865);
and and6528(N10873,N10874,N10875);
and and6536(N10883,N10884,N10885);
and and6544(N10893,N10894,N10895);
and and6552(N10903,N10904,N10905);
and and6560(N10913,N10914,N10915);
and and6568(N10923,N10924,N10925);
and and6576(N10932,N10933,N10934);
and and6584(N10941,N10942,N10943);
and and6592(N10950,N10951,N10952);
and and6600(N10959,N10960,N10961);
and and6608(N10968,N10969,N10970);
and and6615(N10981,N10982,N10983);
and and6622(N10994,N10995,N10996);
and and6629(N11007,N11008,N11009);
and and6636(N11019,N11020,N11021);
and and6643(N11031,N11032,N11033);
and and6650(N11043,N11044,N11045);
and and6657(N11055,N11056,N11057);
and and6664(N11067,N11068,N11069);
and and6671(N11079,N11080,N11081);
and and6678(N11091,N11092,N11093);
and and6685(N11103,N11104,N11105);
and and6692(N11115,N11116,N11117);
and and6699(N11126,N11127,N11128);
and and6706(N11137,N11138,N11139);
and and6713(N11148,N11149,N11150);
and and6720(N11159,N11160,N11161);
and and6727(N11170,N11171,N11172);
and and6734(N11181,N11182,N11183);
and and6741(N11192,N11193,N11194);
and and6748(N11203,N11204,N11205);
and and6755(N11214,N11215,N11216);
and and6762(N11225,N11226,N11227);
and and6769(N11236,N11237,N11238);
and and6776(N11247,N11248,N11249);
and and6783(N11258,N11259,N11260);
and and6790(N11269,N11270,N11271);
and and6797(N11279,N11280,N11281);
and and6804(N11289,N11290,N11291);
and and6811(N11299,N11300,N11301);
and and6818(N11309,N11310,N11311);
and and6825(N11319,N11320,N11321);
and and6832(N11329,N11330,N11331);
and and6839(N11339,N11340,N11341);
and and6846(N11349,N11350,N11351);
and and6853(N11359,N11360,N11361);
and and6860(N11369,N11370,N11371);
and and6867(N11379,N11380,N11381);
and and6874(N11389,N11390,N11391);
and and6881(N11399,N11400,N11401);
and and6888(N11408,N11409,N11410);
and and6894(N11420,N11421,N11422);
and and3303(N5932,N5934,N5935);
and and3304(N5933,N5936,N5937);
and and3312(N5950,N5952,N5953);
and and3313(N5951,N5954,N5955);
and and3321(N5968,N5970,N5971);
and and3322(N5969,N5972,N5973);
and and3330(N5986,N5988,N5989);
and and3331(N5987,N5990,N5991);
and and3339(N6003,N6005,N6006);
and and3340(N6004,N6007,N6008);
and and3348(N6020,N6022,N6023);
and and3349(N6021,N6024,N6025);
and and3357(N6037,N6039,N6040);
and and3358(N6038,N6041,N6042);
and and3366(N6054,N6056,N6057);
and and3367(N6055,N6058,N6059);
and and3375(N6070,N6072,N6073);
and and3376(N6071,N6074,N6075);
and and3384(N6086,N6088,N6089);
and and3385(N6087,N6090,N6091);
and and3393(N6102,N6104,N6105);
and and3394(N6103,N6106,N6107);
and and3402(N6118,N6120,N6121);
and and3403(N6119,N6122,N6123);
and and3411(N6134,N6136,N6137);
and and3412(N6135,N6138,N6139);
and and3420(N6150,N6152,N6153);
and and3421(N6151,N6154,N6155);
and and3429(N6166,N6168,N6169);
and and3430(N6167,N6170,N6171);
and and3438(N6182,N6184,N6185);
and and3439(N6183,N6186,N6187);
and and3447(N6198,N6200,N6201);
and and3448(N6199,N6202,N6203);
and and3456(N6214,N6216,N6217);
and and3457(N6215,N6218,N6219);
and and3465(N6230,N6232,N6233);
and and3466(N6231,N6234,N6235);
and and3474(N6246,N6248,N6249);
and and3475(N6247,N6250,N6251);
and and3483(N6262,N6264,N6265);
and and3484(N6263,N6266,N6267);
and and3492(N6278,N6280,N6281);
and and3493(N6279,N6282,N6283);
and and3501(N6294,N6296,N6297);
and and3502(N6295,N6298,N6299);
and and3510(N6309,N6311,N6312);
and and3511(N6310,N6313,N6314);
and and3519(N6324,N6326,N6327);
and and3520(N6325,N6328,N6329);
and and3528(N6339,N6341,N6342);
and and3529(N6340,N6343,N6344);
and and3537(N6354,N6356,N6357);
and and3538(N6355,N6358,N6359);
and and3546(N6369,N6371,N6372);
and and3547(N6370,N6373,N6374);
and and3555(N6384,N6386,N6387);
and and3556(N6385,N6388,N6389);
and and3564(N6399,N6401,N6402);
and and3565(N6400,N6403,N6404);
and and3573(N6414,N6416,N6417);
and and3574(N6415,N6418,N6419);
and and3582(N6429,N6431,N6432);
and and3583(N6430,N6433,N6434);
and and3591(N6444,N6446,N6447);
and and3592(N6445,N6448,N6449);
and and3600(N6459,N6461,N6462);
and and3601(N6460,N6463,N6464);
and and3609(N6474,N6476,N6477);
and and3610(N6475,N6478,N6479);
and and3618(N6489,N6491,N6492);
and and3619(N6490,N6493,N6494);
and and3627(N6504,N6506,N6507);
and and3628(N6505,N6508,N6509);
and and3636(N6519,N6521,N6522);
and and3637(N6520,N6523,N6524);
and and3645(N6534,N6536,N6537);
and and3646(N6535,N6538,N6539);
and and3654(N6549,N6551,N6552);
and and3655(N6550,N6553,N6554);
and and3663(N6564,N6566,N6567);
and and3664(N6565,N6568,N6569);
and and3672(N6579,N6581,N6582);
and and3673(N6580,N6583,N6584);
and and3681(N6594,N6596,N6597);
and and3682(N6595,N6598,N6599);
and and3690(N6609,N6611,N6612);
and and3691(N6610,N6613,N6614);
and and3699(N6624,N6626,N6627);
and and3700(N6625,N6628,N6629);
and and3708(N6639,N6641,N6642);
and and3709(N6640,N6643,N6644);
and and3717(N6654,N6656,N6657);
and and3718(N6655,N6658,N6659);
and and3726(N6669,N6671,N6672);
and and3727(N6670,N6673,N6674);
and and3735(N6684,N6686,N6687);
and and3736(N6685,N6688,N6689);
and and3744(N6699,N6701,N6702);
and and3745(N6700,N6703,N6704);
and and3753(N6713,N6715,N6716);
and and3754(N6714,N6717,N6718);
and and3762(N6727,N6729,N6730);
and and3763(N6728,N6731,N6732);
and and3771(N6741,N6743,N6744);
and and3772(N6742,N6745,N6746);
and and3780(N6755,N6757,N6758);
and and3781(N6756,N6759,N6760);
and and3789(N6769,N6771,N6772);
and and3790(N6770,N6773,N6774);
and and3798(N6783,N6785,N6786);
and and3799(N6784,N6787,N6788);
and and3807(N6797,N6799,N6800);
and and3808(N6798,N6801,N6802);
and and3816(N6811,N6813,N6814);
and and3817(N6812,N6815,N6816);
and and3825(N6825,N6827,N6828);
and and3826(N6826,N6829,N6830);
and and3834(N6839,N6841,N6842);
and and3835(N6840,N6843,N6844);
and and3843(N6853,N6855,N6856);
and and3844(N6854,N6857,N6858);
and and3852(N6867,N6869,N6870);
and and3853(N6868,N6871,N6872);
and and3861(N6881,N6883,N6884);
and and3862(N6882,N6885,N6886);
and and3870(N6895,N6897,N6898);
and and3871(N6896,N6899,N6900);
and and3879(N6909,N6911,N6912);
and and3880(N6910,N6913,N6914);
and and3888(N6923,N6925,N6926);
and and3889(N6924,N6927,N6928);
and and3897(N6937,N6939,N6940);
and and3898(N6938,N6941,N6942);
and and3906(N6951,N6953,N6954);
and and3907(N6952,N6955,N6956);
and and3915(N6965,N6967,N6968);
and and3916(N6966,N6969,N6970);
and and3924(N6979,N6981,N6982);
and and3925(N6980,N6983,N6984);
and and3933(N6993,N6995,N6996);
and and3934(N6994,N6997,N6998);
and and3942(N7007,N7009,N7010);
and and3943(N7008,N7011,N7012);
and and3951(N7021,N7023,N7024);
and and3952(N7022,N7025,N7026);
and and3960(N7035,N7037,N7038);
and and3961(N7036,N7039,N7040);
and and3969(N7049,N7051,N7052);
and and3970(N7050,N7053,N7054);
and and3978(N7063,N7065,N7066);
and and3979(N7064,N7067,N7068);
and and3987(N7077,N7079,N7080);
and and3988(N7078,N7081,N7082);
and and3996(N7091,N7093,N7094);
and and3997(N7092,N7095,N7096);
and and4005(N7105,N7107,N7108);
and and4006(N7106,N7109,N7110);
and and4014(N7119,N7121,N7122);
and and4015(N7120,N7123,N7124);
and and4023(N7132,N7134,N7135);
and and4024(N7133,N7136,N7137);
and and4032(N7145,N7147,N7148);
and and4033(N7146,N7149,N7150);
and and4041(N7158,N7160,N7161);
and and4042(N7159,N7162,N7163);
and and4050(N7171,N7173,N7174);
and and4051(N7172,N7175,N7176);
and and4059(N7184,N7186,N7187);
and and4060(N7185,N7188,N7189);
and and4068(N7197,N7199,N7200);
and and4069(N7198,N7201,N7202);
and and4077(N7210,N7212,N7213);
and and4078(N7211,N7214,N7215);
and and4086(N7223,N7225,N7226);
and and4087(N7224,N7227,N7228);
and and4095(N7236,N7238,N7239);
and and4096(N7237,N7240,N7241);
and and4104(N7249,N7251,N7252);
and and4105(N7250,N7253,N7254);
and and4113(N7262,N7264,N7265);
and and4114(N7263,N7266,N7267);
and and4122(N7275,N7277,N7278);
and and4123(N7276,N7279,N7280);
and and4131(N7288,N7290,N7291);
and and4132(N7289,N7292,N7293);
and and4140(N7301,N7303,N7304);
and and4141(N7302,N7305,N7306);
and and4149(N7314,N7316,N7317);
and and4150(N7315,N7318,N7319);
and and4158(N7327,N7329,N7330);
and and4159(N7328,N7331,N7332);
and and4167(N7340,N7342,N7343);
and and4168(N7341,N7344,N7345);
and and4176(N7353,N7355,N7356);
and and4177(N7354,N7357,N7358);
and and4185(N7366,N7368,N7369);
and and4186(N7367,N7370,N7371);
and and4194(N7379,N7381,N7382);
and and4195(N7380,N7383,N7384);
and and4203(N7392,N7394,N7395);
and and4204(N7393,N7396,N7397);
and and4212(N7405,N7407,N7408);
and and4213(N7406,N7409,N7410);
and and4221(N7418,N7420,N7421);
and and4222(N7419,N7422,N7423);
and and4230(N7431,N7433,N7434);
and and4231(N7432,N7435,N7436);
and and4239(N7444,N7446,N7447);
and and4240(N7445,N7448,N7449);
and and4248(N7457,N7459,N7460);
and and4249(N7458,N7461,N7462);
and and4257(N7470,N7472,N7473);
and and4258(N7471,N7474,N7475);
and and4266(N7483,N7485,N7486);
and and4267(N7484,N7487,N7488);
and and4275(N7496,N7498,N7499);
and and4276(N7497,N7500,N7501);
and and4284(N7509,N7511,N7512);
and and4285(N7510,N7513,N7514);
and and4293(N7522,N7524,N7525);
and and4294(N7523,N7526,N7527);
and and4302(N7535,N7537,N7538);
and and4303(N7536,N7539,N7540);
and and4311(N7548,N7550,N7551);
and and4312(N7549,N7552,N7553);
and and4320(N7561,N7563,N7564);
and and4321(N7562,N7565,N7566);
and and4329(N7574,N7576,N7577);
and and4330(N7575,N7578,N7579);
and and4338(N7587,N7589,N7590);
and and4339(N7588,N7591,N7592);
and and4347(N7600,N7602,N7603);
and and4348(N7601,N7604,N7605);
and and4356(N7613,N7615,N7616);
and and4357(N7614,N7617,N7618);
and and4365(N7625,N7627,N7628);
and and4366(N7626,N7629,N7630);
and and4374(N7637,N7639,N7640);
and and4375(N7638,N7641,N7642);
and and4383(N7649,N7651,N7652);
and and4384(N7650,N7653,N7654);
and and4392(N7661,N7663,N7664);
and and4393(N7662,N7665,N7666);
and and4401(N7673,N7675,N7676);
and and4402(N7674,N7677,N7678);
and and4410(N7685,N7687,N7688);
and and4411(N7686,N7689,N7690);
and and4419(N7697,N7699,N7700);
and and4420(N7698,N7701,N7702);
and and4428(N7709,N7711,N7712);
and and4429(N7710,N7713,N7714);
and and4437(N7721,N7723,N7724);
and and4438(N7722,N7725,N7726);
and and4446(N7733,N7735,N7736);
and and4447(N7734,N7737,N7738);
and and4455(N7745,N7747,N7748);
and and4456(N7746,N7749,N7750);
and and4464(N7757,N7759,N7760);
and and4465(N7758,N7761,N7762);
and and4473(N7769,N7771,N7772);
and and4474(N7770,N7773,N7774);
and and4482(N7781,N7783,N7784);
and and4483(N7782,N7785,N7786);
and and4491(N7793,N7795,N7796);
and and4492(N7794,N7797,N7798);
and and4500(N7805,N7807,N7808);
and and4501(N7806,N7809,N7810);
and and4509(N7817,N7819,N7820);
and and4510(N7818,N7821,N7822);
and and4518(N7829,N7831,N7832);
and and4519(N7830,N7833,N7834);
and and4527(N7841,N7843,N7844);
and and4528(N7842,N7845,N7846);
and and4536(N7853,N7855,N7856);
and and4537(N7854,N7857,N7858);
and and4545(N7865,N7867,N7868);
and and4546(N7866,N7869,N7870);
and and4554(N7877,N7879,N7880);
and and4555(N7878,N7881,N7882);
and and4563(N7889,N7891,N7892);
and and4564(N7890,N7893,N7894);
and and4572(N7901,N7903,N7904);
and and4573(N7902,N7905,N7906);
and and4581(N7912,N7914,N7915);
and and4582(N7913,N7916,N7917);
and and4590(N7923,N7925,N7926);
and and4591(N7924,N7927,N7928);
and and4599(N7934,N7936,N7937);
and and4600(N7935,N7938,N7939);
and and4608(N7945,N7947,N7948);
and and4609(N7946,N7949,N7950);
and and4617(N7956,N7958,N7959);
and and4618(N7957,N7960,N7961);
and and4626(N7967,N7969,N7970);
and and4627(N7968,N7971,N7972);
and and4635(N7978,N7980,N7981);
and and4636(N7979,N7982,N7983);
and and4644(N7989,N7991,N7992);
and and4645(N7990,N7993,N7994);
and and4653(N8000,N8002,N8003);
and and4654(N8001,N8004,N8005);
and and4662(N8011,N8013,N8014);
and and4663(N8012,N8015,N8016);
and and4671(N8022,N8024,N8025);
and and4672(N8023,N8026,N8027);
and and4680(N8033,N8035,N8036);
and and4681(N8034,N8037,N8038);
and and4689(N8043,N8045,N8046);
and and4690(N8044,N8047,N8048);
and and4698(N8053,N8055,N8056);
and and4699(N8054,N8057,N8058);
and and4707(N8063,N8065,N8066);
and and4708(N8064,N8067,N8068);
and and4716(N8073,N8075,N8076);
and and4717(N8074,N8077,N8078);
and and4725(N8083,N8085,N8086);
and and4726(N8084,N8087,N8088);
and and4734(N8093,N8095,N8096);
and and4735(N8094,N8097,N8098);
and and4743(N8103,N8105,N8106);
and and4744(N8104,N8107,N8108);
and and4752(N8113,N8115,N8116);
and and4753(N8114,N8117,N8118);
and and4761(N8122,N8124,N8125);
and and4762(N8123,N8126,N8127);
and and4769(N8138,N8140,N8141);
and and4770(N8139,N8142,N8143);
and and4777(N8154,N8156,N8157);
and and4778(N8155,N8158,N8159);
and and4785(N8169,N8171,N8172);
and and4786(N8170,N8173,N8174);
and and4793(N8184,N8186,N8187);
and and4794(N8185,N8188,N8189);
and and4801(N8199,N8201,N8202);
and and4802(N8200,N8203,N8204);
and and4809(N8214,N8216,N8217);
and and4810(N8215,N8218,N8219);
and and4817(N8229,N8231,N8232);
and and4818(N8230,N8233,N8234);
and and4825(N8244,N8246,N8247);
and and4826(N8245,N8248,N8249);
and and4833(N8259,N8261,N8262);
and and4834(N8260,N8263,N8264);
and and4841(N8274,N8276,N8277);
and and4842(N8275,N8278,N8279);
and and4849(N8289,N8291,N8292);
and and4850(N8290,N8293,N8294);
and and4857(N8304,N8306,N8307);
and and4858(N8305,N8308,N8309);
and and4865(N8319,N8321,N8322);
and and4866(N8320,N8323,N8324);
and and4873(N8334,N8336,N8337);
and and4874(N8335,N8338,N8339);
and and4881(N8349,N8351,N8352);
and and4882(N8350,N8353,N8354);
and and4889(N8364,N8366,N8367);
and and4890(N8365,N8368,N8369);
and and4897(N8378,N8380,N8381);
and and4898(N8379,N8382,N8383);
and and4905(N8392,N8394,N8395);
and and4906(N8393,N8396,N8397);
and and4913(N8406,N8408,N8409);
and and4914(N8407,N8410,N8411);
and and4921(N8420,N8422,N8423);
and and4922(N8421,N8424,N8425);
and and4929(N8434,N8436,N8437);
and and4930(N8435,N8438,N8439);
and and4937(N8448,N8450,N8451);
and and4938(N8449,N8452,N8453);
and and4945(N8462,N8464,N8465);
and and4946(N8463,N8466,N8467);
and and4953(N8476,N8478,N8479);
and and4954(N8477,N8480,N8481);
and and4961(N8490,N8492,N8493);
and and4962(N8491,N8494,N8495);
and and4969(N8504,N8506,N8507);
and and4970(N8505,N8508,N8509);
and and4977(N8518,N8520,N8521);
and and4978(N8519,N8522,N8523);
and and4985(N8532,N8534,N8535);
and and4986(N8533,N8536,N8537);
and and4993(N8546,N8548,N8549);
and and4994(N8547,N8550,N8551);
and and5001(N8560,N8562,N8563);
and and5002(N8561,N8564,N8565);
and and5009(N8574,N8576,N8577);
and and5010(N8575,N8578,N8579);
and and5017(N8588,N8590,N8591);
and and5018(N8589,N8592,N8593);
and and5025(N8602,N8604,N8605);
and and5026(N8603,N8606,N8607);
and and5033(N8616,N8618,N8619);
and and5034(N8617,N8620,N8621);
and and5041(N8630,N8632,N8633);
and and5042(N8631,N8634,N8635);
and and5049(N8644,N8646,N8647);
and and5050(N8645,N8648,N8649);
and and5057(N8658,N8660,N8661);
and and5058(N8659,N8662,N8663);
and and5065(N8672,N8674,N8675);
and and5066(N8673,N8676,N8677);
and and5073(N8686,N8688,N8689);
and and5074(N8687,N8690,N8691);
and and5081(N8700,N8702,N8703);
and and5082(N8701,N8704,N8705);
and and5089(N8714,N8716,N8717);
and and5090(N8715,N8718,N8719);
and and5097(N8728,N8730,N8731);
and and5098(N8729,N8732,N8733);
and and5105(N8742,N8744,N8745);
and and5106(N8743,N8746,N8747);
and and5113(N8756,N8758,N8759);
and and5114(N8757,N8760,N8761);
and and5121(N8770,N8772,N8773);
and and5122(N8771,N8774,N8775);
and and5129(N8784,N8786,N8787);
and and5130(N8785,N8788,N8789);
and and5137(N8798,N8800,N8801);
and and5138(N8799,N8802,N8803);
and and5145(N8812,N8814,N8815);
and and5146(N8813,N8816,N8817);
and and5153(N8826,N8828,N8829);
and and5154(N8827,N8830,N8831);
and and5161(N8840,N8842,N8843);
and and5162(N8841,N8844,N8845);
and and5169(N8854,N8856,N8857);
and and5170(N8855,N8858,N8859);
and and5177(N8868,N8870,N8871);
and and5178(N8869,N8872,N8873);
and and5185(N8882,N8884,N8885);
and and5186(N8883,N8886,N8887);
and and5193(N8896,N8898,N8899);
and and5194(N8897,N8900,N8901);
and and5201(N8909,N8911,N8912);
and and5202(N8910,N8913,N8914);
and and5209(N8922,N8924,N8925);
and and5210(N8923,N8926,N8927);
and and5217(N8935,N8937,N8938);
and and5218(N8936,N8939,N8940);
and and5225(N8948,N8950,N8951);
and and5226(N8949,N8952,N8953);
and and5233(N8961,N8963,N8964);
and and5234(N8962,N8965,N8966);
and and5241(N8974,N8976,N8977);
and and5242(N8975,N8978,N8979);
and and5249(N8987,N8989,N8990);
and and5250(N8988,N8991,N8992);
and and5257(N9000,N9002,N9003);
and and5258(N9001,N9004,N9005);
and and5265(N9013,N9015,N9016);
and and5266(N9014,N9017,N9018);
and and5273(N9026,N9028,N9029);
and and5274(N9027,N9030,N9031);
and and5281(N9039,N9041,N9042);
and and5282(N9040,N9043,N9044);
and and5289(N9052,N9054,N9055);
and and5290(N9053,N9056,N9057);
and and5297(N9065,N9067,N9068);
and and5298(N9066,N9069,N9070);
and and5305(N9078,N9080,N9081);
and and5306(N9079,N9082,N9083);
and and5313(N9091,N9093,N9094);
and and5314(N9092,N9095,N9096);
and and5321(N9104,N9106,N9107);
and and5322(N9105,N9108,N9109);
and and5329(N9117,N9119,N9120);
and and5330(N9118,N9121,N9122);
and and5337(N9130,N9132,N9133);
and and5338(N9131,N9134,N9135);
and and5345(N9143,N9145,N9146);
and and5346(N9144,N9147,N9148);
and and5353(N9156,N9158,N9159);
and and5354(N9157,N9160,N9161);
and and5361(N9169,N9171,N9172);
and and5362(N9170,N9173,N9174);
and and5369(N9182,N9184,N9185);
and and5370(N9183,N9186,N9187);
and and5377(N9195,N9197,N9198);
and and5378(N9196,N9199,N9200);
and and5385(N9208,N9210,N9211);
and and5386(N9209,N9212,N9213);
and and5393(N9221,N9223,N9224);
and and5394(N9222,N9225,N9226);
and and5401(N9234,N9236,N9237);
and and5402(N9235,N9238,N9239);
and and5409(N9247,N9249,N9250);
and and5410(N9248,N9251,N9252);
and and5417(N9260,N9262,N9263);
and and5418(N9261,N9264,N9265);
and and5425(N9273,N9275,N9276);
and and5426(N9274,N9277,N9278);
and and5433(N9286,N9288,N9289);
and and5434(N9287,N9290,N9291);
and and5441(N9299,N9301,N9302);
and and5442(N9300,N9303,N9304);
and and5449(N9312,N9314,N9315);
and and5450(N9313,N9316,N9317);
and and5457(N9325,N9327,N9328);
and and5458(N9326,N9329,N9330);
and and5465(N9338,N9340,N9341);
and and5466(N9339,N9342,N9343);
and and5473(N9351,N9353,N9354);
and and5474(N9352,N9355,N9356);
and and5481(N9364,N9366,N9367);
and and5482(N9365,N9368,N9369);
and and5489(N9377,N9379,N9380);
and and5490(N9378,N9381,N9382);
and and5497(N9390,N9392,N9393);
and and5498(N9391,N9394,N9395);
and and5505(N9403,N9405,N9406);
and and5506(N9404,N9407,N9408);
and and5513(N9416,N9418,N9419);
and and5514(N9417,N9420,N9421);
and and5521(N9429,N9431,N9432);
and and5522(N9430,N9433,N9434);
and and5529(N9442,N9444,N9445);
and and5530(N9443,N9446,N9447);
and and5537(N9455,N9457,N9458);
and and5538(N9456,N9459,N9460);
and and5545(N9468,N9470,N9471);
and and5546(N9469,N9472,N9473);
and and5553(N9481,N9483,N9484);
and and5554(N9482,N9485,N9486);
and and5561(N9494,N9496,N9497);
and and5562(N9495,N9498,N9499);
and and5569(N9507,N9509,N9510);
and and5570(N9508,N9511,N9512);
and and5577(N9520,N9522,N9523);
and and5578(N9521,N9524,N9525);
and and5585(N9533,N9535,N9536);
and and5586(N9534,N9537,N9538);
and and5593(N9546,N9548,N9549);
and and5594(N9547,N9550,N9551);
and and5601(N9559,N9561,N9562);
and and5602(N9560,N9563,N9564);
and and5609(N9572,N9574,N9575);
and and5610(N9573,N9576,N9577);
and and5617(N9585,N9587,N9588);
and and5618(N9586,N9589,N9590);
and and5625(N9598,N9600,N9601);
and and5626(N9599,N9602,N9603);
and and5633(N9611,N9613,N9614);
and and5634(N9612,N9615,N9616);
and and5641(N9624,N9626,N9627);
and and5642(N9625,N9628,N9629);
and and5649(N9637,N9639,N9640);
and and5650(N9638,N9641,N9642);
and and5657(N9649,N9651,N9652);
and and5658(N9650,N9653,N9654);
and and5665(N9661,N9663,N9664);
and and5666(N9662,N9665,N9666);
and and5673(N9673,N9675,N9676);
and and5674(N9674,N9677,N9678);
and and5681(N9685,N9687,N9688);
and and5682(N9686,N9689,N9690);
and and5689(N9697,N9699,N9700);
and and5690(N9698,N9701,N9702);
and and5697(N9709,N9711,N9712);
and and5698(N9710,N9713,N9714);
and and5705(N9721,N9723,N9724);
and and5706(N9722,N9725,N9726);
and and5713(N9733,N9735,N9736);
and and5714(N9734,N9737,N9738);
and and5721(N9745,N9747,N9748);
and and5722(N9746,N9749,N9750);
and and5729(N9757,N9759,N9760);
and and5730(N9758,N9761,N9762);
and and5737(N9769,N9771,N9772);
and and5738(N9770,N9773,N9774);
and and5745(N9781,N9783,N9784);
and and5746(N9782,N9785,N9786);
and and5753(N9793,N9795,N9796);
and and5754(N9794,N9797,N9798);
and and5761(N9805,N9807,N9808);
and and5762(N9806,N9809,N9810);
and and5769(N9817,N9819,N9820);
and and5770(N9818,N9821,N9822);
and and5777(N9829,N9831,N9832);
and and5778(N9830,N9833,N9834);
and and5785(N9841,N9843,N9844);
and and5786(N9842,N9845,N9846);
and and5793(N9853,N9855,N9856);
and and5794(N9854,N9857,N9858);
and and5801(N9865,N9867,N9868);
and and5802(N9866,N9869,N9870);
and and5809(N9877,N9879,N9880);
and and5810(N9878,N9881,N9882);
and and5817(N9889,N9891,N9892);
and and5818(N9890,N9893,N9894);
and and5825(N9901,N9903,N9904);
and and5826(N9902,N9905,N9906);
and and5833(N9913,N9915,N9916);
and and5834(N9914,N9917,N9918);
and and5841(N9925,N9927,N9928);
and and5842(N9926,N9929,N9930);
and and5849(N9937,N9939,N9940);
and and5850(N9938,N9941,N9942);
and and5857(N9949,N9951,N9952);
and and5858(N9950,N9953,N9954);
and and5865(N9961,N9963,N9964);
and and5866(N9962,N9965,N9966);
and and5873(N9973,N9975,N9976);
and and5874(N9974,N9977,N9978);
and and5881(N9985,N9987,N9988);
and and5882(N9986,N9989,N9990);
and and5889(N9997,N9999,N10000);
and and5890(N9998,N10001,N10002);
and and5897(N10009,N10011,N10012);
and and5898(N10010,N10013,N10014);
and and5905(N10021,N10023,N10024);
and and5906(N10022,N10025,N10026);
and and5913(N10033,N10035,N10036);
and and5914(N10034,N10037,N10038);
and and5921(N10045,N10047,N10048);
and and5922(N10046,N10049,N10050);
and and5929(N10057,N10059,N10060);
and and5930(N10058,N10061,N10062);
and and5937(N10069,N10071,N10072);
and and5938(N10070,N10073,N10074);
and and5945(N10081,N10083,N10084);
and and5946(N10082,N10085,N10086);
and and5953(N10093,N10095,N10096);
and and5954(N10094,N10097,N10098);
and and5961(N10105,N10107,N10108);
and and5962(N10106,N10109,N10110);
and and5969(N10117,N10119,N10120);
and and5970(N10118,N10121,N10122);
and and5977(N10129,N10131,N10132);
and and5978(N10130,N10133,N10134);
and and5985(N10141,N10143,N10144);
and and5986(N10142,N10145,N10146);
and and5993(N10153,N10155,N10156);
and and5994(N10154,N10157,N10158);
and and6001(N10165,N10167,N10168);
and and6002(N10166,N10169,N10170);
and and6009(N10177,N10179,N10180);
and and6010(N10178,N10181,N10182);
and and6017(N10189,N10191,N10192);
and and6018(N10190,N10193,N10194);
and and6025(N10201,N10203,N10204);
and and6026(N10202,N10205,N10206);
and and6033(N10212,N10214,N10215);
and and6034(N10213,N10216,N10217);
and and6041(N10223,N10225,N10226);
and and6042(N10224,N10227,N10228);
and and6049(N10234,N10236,N10237);
and and6050(N10235,N10238,N10239);
and and6057(N10245,N10247,N10248);
and and6058(N10246,N10249,N10250);
and and6065(N10256,N10258,N10259);
and and6066(N10257,N10260,N10261);
and and6073(N10267,N10269,N10270);
and and6074(N10268,N10271,N10272);
and and6081(N10278,N10280,N10281);
and and6082(N10279,N10282,N10283);
and and6089(N10289,N10291,N10292);
and and6090(N10290,N10293,N10294);
and and6097(N10300,N10302,N10303);
and and6098(N10301,N10304,N10305);
and and6105(N10311,N10313,N10314);
and and6106(N10312,N10315,N10316);
and and6113(N10322,N10324,N10325);
and and6114(N10323,N10326,N10327);
and and6121(N10333,N10335,N10336);
and and6122(N10334,N10337,N10338);
and and6129(N10344,N10346,N10347);
and and6130(N10345,N10348,N10349);
and and6137(N10355,N10357,N10358);
and and6138(N10356,N10359,N10360);
and and6145(N10366,N10368,N10369);
and and6146(N10367,N10370,N10371);
and and6153(N10377,N10379,N10380);
and and6154(N10378,N10381,N10382);
and and6161(N10388,N10390,N10391);
and and6162(N10389,N10392,N10393);
and and6169(N10399,N10401,N10402);
and and6170(N10400,N10403,N10404);
and and6177(N10410,N10412,N10413);
and and6178(N10411,N10414,N10415);
and and6185(N10421,N10423,N10424);
and and6186(N10422,N10425,N10426);
and and6193(N10432,N10434,N10435);
and and6194(N10433,N10436,N10437);
and and6201(N10443,N10445,N10446);
and and6202(N10444,N10447,N10448);
and and6209(N10454,N10456,N10457);
and and6210(N10455,N10458,N10459);
and and6217(N10465,N10467,N10468);
and and6218(N10466,N10469,N10470);
and and6225(N10476,N10478,N10479);
and and6226(N10477,N10480,N10481);
and and6233(N10487,N10489,N10490);
and and6234(N10488,N10491,N10492);
and and6241(N10498,N10500,N10501);
and and6242(N10499,N10502,N10503);
and and6249(N10509,N10511,N10512);
and and6250(N10510,N10513,N10514);
and and6257(N10520,N10522,N10523);
and and6258(N10521,N10524,N10525);
and and6265(N10531,N10533,N10534);
and and6266(N10532,N10535,N10536);
and and6273(N10542,N10544,N10545);
and and6274(N10543,N10546,N10547);
and and6281(N10553,N10555,N10556);
and and6282(N10554,N10557,N10558);
and and6289(N10564,N10566,N10567);
and and6290(N10565,N10568,N10569);
and and6297(N10575,N10577,N10578);
and and6298(N10576,N10579,N10580);
and and6305(N10586,N10588,N10589);
and and6306(N10587,N10590,N10591);
and and6313(N10597,N10599,N10600);
and and6314(N10598,N10601,N10602);
and and6321(N10608,N10610,N10611);
and and6322(N10609,N10612,N10613);
and and6329(N10619,N10621,N10622);
and and6330(N10620,N10623,N10624);
and and6337(N10630,N10632,N10633);
and and6338(N10631,N10634,N10635);
and and6345(N10641,N10643,N10644);
and and6346(N10642,N10645,N10646);
and and6353(N10652,N10654,N10655);
and and6354(N10653,N10656,N10657);
and and6361(N10663,N10665,N10666);
and and6362(N10664,N10667,N10668);
and and6369(N10674,N10676,N10677);
and and6370(N10675,N10678,N10679);
and and6377(N10684,N10686,N10687);
and and6378(N10685,N10688,N10689);
and and6385(N10694,N10696,N10697);
and and6386(N10695,N10698,N10699);
and and6393(N10704,N10706,N10707);
and and6394(N10705,N10708,N10709);
and and6401(N10714,N10716,N10717);
and and6402(N10715,N10718,N10719);
and and6409(N10724,N10726,N10727);
and and6410(N10725,N10728,N10729);
and and6417(N10734,N10736,N10737);
and and6418(N10735,N10738,N10739);
and and6425(N10744,N10746,N10747);
and and6426(N10745,N10748,N10749);
and and6433(N10754,N10756,N10757);
and and6434(N10755,N10758,N10759);
and and6441(N10764,N10766,N10767);
and and6442(N10765,N10768,N10769);
and and6449(N10774,N10776,N10777);
and and6450(N10775,N10778,N10779);
and and6457(N10784,N10786,N10787);
and and6458(N10785,N10788,N10789);
and and6465(N10794,N10796,N10797);
and and6466(N10795,N10798,N10799);
and and6473(N10804,N10806,N10807);
and and6474(N10805,N10808,N10809);
and and6481(N10814,N10816,N10817);
and and6482(N10815,N10818,N10819);
and and6489(N10824,N10826,N10827);
and and6490(N10825,N10828,N10829);
and and6497(N10834,N10836,N10837);
and and6498(N10835,N10838,N10839);
and and6505(N10844,N10846,N10847);
and and6506(N10845,N10848,N10849);
and and6513(N10854,N10856,N10857);
and and6514(N10855,N10858,N10859);
and and6521(N10864,N10866,N10867);
and and6522(N10865,N10868,N10869);
and and6529(N10874,N10876,N10877);
and and6530(N10875,N10878,N10879);
and and6537(N10884,N10886,N10887);
and and6538(N10885,N10888,N10889);
and and6545(N10894,N10896,N10897);
and and6546(N10895,N10898,N10899);
and and6553(N10904,N10906,N10907);
and and6554(N10905,N10908,N10909);
and and6561(N10914,N10916,N10917);
and and6562(N10915,N10918,N10919);
and and6569(N10924,N10926,N10927);
and and6570(N10925,N10928,N10929);
and and6577(N10933,N10935,N10936);
and and6578(N10934,N10937,N10938);
and and6585(N10942,N10944,N10945);
and and6586(N10943,N10946,N10947);
and and6593(N10951,N10953,N10954);
and and6594(N10952,N10955,N10956);
and and6601(N10960,N10962,N10963);
and and6602(N10961,N10964,N10965);
and and6609(N10969,N10971,N10972);
and and6610(N10970,N10973,N10974);
and and6616(N10982,N10984,N10985);
and and6617(N10983,N10986,N10987);
and and6623(N10995,N10997,N10998);
and and6624(N10996,N10999,N11000);
and and6630(N11008,N11010,N11011);
and and6631(N11009,N11012,N11013);
and and6637(N11020,N11022,N11023);
and and6638(N11021,N11024,N11025);
and and6644(N11032,N11034,N11035);
and and6645(N11033,N11036,N11037);
and and6651(N11044,N11046,N11047);
and and6652(N11045,N11048,N11049);
and and6658(N11056,N11058,N11059);
and and6659(N11057,N11060,N11061);
and and6665(N11068,N11070,N11071);
and and6666(N11069,N11072,N11073);
and and6672(N11080,N11082,N11083);
and and6673(N11081,N11084,N11085);
and and6679(N11092,N11094,N11095);
and and6680(N11093,N11096,N11097);
and and6686(N11104,N11106,N11107);
and and6687(N11105,N11108,N11109);
and and6693(N11116,N11118,N11119);
and and6694(N11117,N11120,N11121);
and and6700(N11127,N11129,N11130);
and and6701(N11128,N11131,N11132);
and and6707(N11138,N11140,N11141);
and and6708(N11139,N11142,N11143);
and and6714(N11149,N11151,N11152);
and and6715(N11150,N11153,N11154);
and and6721(N11160,N11162,N11163);
and and6722(N11161,N11164,N11165);
and and6728(N11171,N11173,N11174);
and and6729(N11172,N11175,N11176);
and and6735(N11182,N11184,N11185);
and and6736(N11183,N11186,N11187);
and and6742(N11193,N11195,N11196);
and and6743(N11194,N11197,N11198);
and and6749(N11204,N11206,N11207);
and and6750(N11205,N11208,N11209);
and and6756(N11215,N11217,N11218);
and and6757(N11216,N11219,N11220);
and and6763(N11226,N11228,N11229);
and and6764(N11227,N11230,N11231);
and and6770(N11237,N11239,N11240);
and and6771(N11238,N11241,N11242);
and and6777(N11248,N11250,N11251);
and and6778(N11249,N11252,N11253);
and and6784(N11259,N11261,N11262);
and and6785(N11260,N11263,N11264);
and and6791(N11270,N11272,N11273);
and and6792(N11271,N11274,N11275);
and and6798(N11280,N11282,N11283);
and and6799(N11281,N11284,N11285);
and and6805(N11290,N11292,N11293);
and and6806(N11291,N11294,N11295);
and and6812(N11300,N11302,N11303);
and and6813(N11301,N11304,N11305);
and and6819(N11310,N11312,N11313);
and and6820(N11311,N11314,N11315);
and and6826(N11320,N11322,N11323);
and and6827(N11321,N11324,N11325);
and and6833(N11330,N11332,N11333);
and and6834(N11331,N11334,N11335);
and and6840(N11340,N11342,N11343);
and and6841(N11341,N11344,N11345);
and and6847(N11350,N11352,N11353);
and and6848(N11351,N11354,N11355);
and and6854(N11360,N11362,N11363);
and and6855(N11361,N11364,N11365);
and and6861(N11370,N11372,N11373);
and and6862(N11371,N11374,N11375);
and and6868(N11380,N11382,N11383);
and and6869(N11381,N11384,N11385);
and and6875(N11390,N11392,N11393);
and and6876(N11391,N11394,N11395);
and and6882(N11400,N11402,N11403);
and and6883(N11401,N11404,N11405);
and and6889(N11409,N11411,N11412);
and and6890(N11410,N11413,in0);
and and6895(N11421,N11423,N11424);
and and6896(N11422,N11425,in0);
and and3305(N5934,N5938,N5939);
and and3306(N5935,N5940,N5941);
and and3307(N5936,N5942,R1);
and and3308(N5937,N5943,N5944);
and and3314(N5952,N5956,N5957);
and and3315(N5953,N5958,N5959);
and and3316(N5954,N5960,N5961);
and and3317(N5955,N5962,R2);
and and3323(N5970,N5974,N5975);
and and3324(N5971,N5976,N5977);
and and3325(N5972,N5978,N5979);
and and3326(N5973,N5980,N5981);
and and3332(N5988,N5992,N5993);
and and3333(N5989,N5994,N5995);
and and3334(N5990,R0,N5996);
and and3335(N5991,N5997,N5998);
and and3341(N6005,N6009,N6010);
and and3342(N6006,N6011,N6012);
and and3343(N6007,N6013,R0);
and and3344(N6008,N6014,R2);
and and3350(N6022,N6026,N6027);
and and3351(N6023,N6028,N6029);
and and3352(N6024,N6030,N6031);
and and3353(N6025,N6032,N6033);
and and3359(N6039,N6043,N6044);
and and3360(N6040,N6045,N6046);
and and3361(N6041,N6047,R1);
and and3362(N6042,N6048,N6049);
and and3368(N6056,N6060,N6061);
and and3369(N6057,N6062,in2);
and and3370(N6058,N6063,R1);
and and3371(N6059,N6064,R3);
and and3377(N6072,N6076,N6077);
and and3378(N6073,N6078,N6079);
and and3379(N6074,R0,N6080);
and and3380(N6075,R2,N6081);
and and3386(N6088,N6092,N6093);
and and3387(N6089,in1,N6094);
and and3388(N6090,N6095,N6096);
and and3389(N6091,N6097,R3);
and and3395(N6104,N6108,N6109);
and and3396(N6105,N6110,in1);
and and3397(N6106,N6111,N6112);
and and3398(N6107,N6113,R3);
and and3404(N6120,N6124,N6125);
and and3405(N6121,N6126,N6127);
and and3406(N6122,R0,N6128);
and and3407(N6123,R2,N6129);
and and3413(N6136,N6140,N6141);
and and3414(N6137,N6142,in2);
and and3415(N6138,N6143,R1);
and and3416(N6139,R2,N6144);
and and3422(N6152,N6156,N6157);
and and3423(N6153,in0,N6158);
and and3424(N6154,N6159,N6160);
and and3425(N6155,R2,N6161);
and and3431(N6168,N6172,N6173);
and and3432(N6169,N6174,N6175);
and and3433(N6170,R0,N6176);
and and3434(N6171,N6177,R3);
and and3440(N6184,N6188,N6189);
and and3441(N6185,N6190,in2);
and and3442(N6186,N6191,N6192);
and and3443(N6187,N6193,N6194);
and and3449(N6200,N6204,N6205);
and and3450(N6201,N6206,N6207);
and and3451(N6202,N6208,N6209);
and and3452(N6203,N6210,R3);
and and3458(N6216,N6220,N6221);
and and3459(N6217,N6222,N6223);
and and3460(N6218,N6224,N6225);
and and3461(N6219,N6226,R3);
and and3467(N6232,N6236,N6237);
and and3468(N6233,N6238,N6239);
and and3469(N6234,N6240,N6241);
and and3470(N6235,R1,N6242);
and and3476(N6248,N6252,N6253);
and and3477(N6249,N6254,in1);
and and3478(N6250,N6255,N6256);
and and3479(N6251,N6257,N6258);
and and3485(N6264,N6268,N6269);
and and3486(N6265,N6270,in1);
and and3487(N6266,in2,N6271);
and and3488(N6267,N6272,N6273);
and and3494(N6280,N6284,N6285);
and and3495(N6281,N6286,N6287);
and and3496(N6282,N6288,N6289);
and and3497(N6283,R2,R3);
and and3503(N6296,N6300,N6301);
and and3504(N6297,N6302,in2);
and and3505(N6298,N6303,N6304);
and and3506(N6299,R2,R3);
and and3512(N6311,N6315,N6316);
and and3513(N6312,in0,N6317);
and and3514(N6313,N6318,R0);
and and3515(N6314,R1,R3);
and and3521(N6326,N6330,N6331);
and and3522(N6327,N6332,N6333);
and and3523(N6328,R0,R1);
and and3524(N6329,R2,N6334);
and and3530(N6341,N6345,N6346);
and and3531(N6342,N6347,N6348);
and and3532(N6343,N6349,R1);
and and3533(N6344,N6350,R3);
and and3539(N6356,N6360,N6361);
and and3540(N6357,N6362,in1);
and and3541(N6358,N6363,R0);
and and3542(N6359,N6364,N6365);
and and3548(N6371,N6375,N6376);
and and3549(N6372,N6377,N6378);
and and3550(N6373,in2,N6379);
and and3551(N6374,N6380,R3);
and and3557(N6386,N6390,N6391);
and and3558(N6387,N6392,N6393);
and and3559(N6388,N6394,R1);
and and3560(N6389,N6395,N6396);
and and3566(N6401,N6405,N6406);
and and3567(N6402,N6407,N6408);
and and3568(N6403,N6409,N6410);
and and3569(N6404,R1,R2);
and and3575(N6416,N6420,N6421);
and and3576(N6417,N6422,in1);
and and3577(N6418,R0,R1);
and and3578(N6419,N6423,N6424);
and and3584(N6431,N6435,N6436);
and and3585(N6432,N6437,in2);
and and3586(N6433,R0,R1);
and and3587(N6434,N6438,N6439);
and and3593(N6446,N6450,N6451);
and and3594(N6447,N6452,in2);
and and3595(N6448,N6453,N6454);
and and3596(N6449,N6455,R3);
and and3602(N6461,N6465,N6466);
and and3603(N6462,in0,N6467);
and and3604(N6463,N6468,N6469);
and and3605(N6464,N6470,R3);
and and3611(N6476,N6480,N6481);
and and3612(N6477,N6482,N6483);
and and3613(N6478,N6484,N6485);
and and3614(N6479,N6486,R2);
and and3620(N6491,N6495,N6496);
and and3621(N6492,N6497,N6498);
and and3622(N6493,in2,N6499);
and and3623(N6494,N6500,R2);
and and3629(N6506,N6510,N6511);
and and3630(N6507,in1,N6512);
and and3631(N6508,R0,N6513);
and and3632(N6509,R2,N6514);
and and3638(N6521,N6525,N6526);
and and3639(N6522,N6527,N6528);
and and3640(N6523,N6529,N6530);
and and3641(N6524,N6531,R3);
and and3647(N6536,N6540,N6541);
and and3648(N6537,N6542,in1);
and and3649(N6538,in2,N6543);
and and3650(N6539,R1,N6544);
and and3656(N6551,N6555,N6556);
and and3657(N6552,N6557,in1);
and and3658(N6553,N6558,N6559);
and and3659(N6554,N6560,R3);
and and3665(N6566,N6570,N6571);
and and3666(N6567,N6572,N6573);
and and3667(N6568,N6574,N6575);
and and3668(N6569,R2,N6576);
and and3674(N6581,N6585,N6586);
and and3675(N6582,in1,N6587);
and and3676(N6583,N6588,R1);
and and3677(N6584,R2,N6589);
and and3683(N6596,N6600,N6601);
and and3684(N6597,in0,in1);
and and3685(N6598,in2,N6602);
and and3686(N6599,N6603,N6604);
and and3692(N6611,N6615,N6616);
and and3693(N6612,N6617,in1);
and and3694(N6613,in2,N6618);
and and3695(N6614,R1,N6619);
and and3701(N6626,N6630,N6631);
and and3702(N6627,N6632,N6633);
and and3703(N6628,in2,N6634);
and and3704(N6629,N6635,R2);
and and3710(N6641,N6645,N6646);
and and3711(N6642,N6647,N6648);
and and3712(N6643,in2,R0);
and and3713(N6644,N6649,R2);
and and3719(N6656,N6660,N6661);
and and3720(N6657,N6662,N6663);
and and3721(N6658,R0,R1);
and and3722(N6659,N6664,N6665);
and and3728(N6671,N6675,N6676);
and and3729(N6672,N6677,N6678);
and and3730(N6673,in2,N6679);
and and3731(N6674,N6680,R2);
and and3737(N6686,N6690,N6691);
and and3738(N6687,N6692,N6693);
and and3739(N6688,in2,N6694);
and and3740(N6689,R1,R2);
and and3746(N6701,N6705,N6706);
and and3747(N6702,N6707,in1);
and and3748(N6703,in2,N6708);
and and3749(N6704,R1,R2);
and and3755(N6715,N6719,N6720);
and and3756(N6716,in1,N6721);
and and3757(N6717,R0,N6722);
and and3758(N6718,N6723,R3);
and and3764(N6729,N6733,N6734);
and and3765(N6730,N6735,in2);
and and3766(N6731,R0,N6736);
and and3767(N6732,R2,R3);
and and3773(N6743,N6747,N6748);
and and3774(N6744,N6749,in2);
and and3775(N6745,R0,R1);
and and3776(N6746,N6750,N6751);
and and3782(N6757,N6761,N6762);
and and3783(N6758,N6763,N6764);
and and3784(N6759,R0,R1);
and and3785(N6760,R2,N6765);
and and3791(N6771,N6775,N6776);
and and3792(N6772,in0,N6777);
and and3793(N6773,in2,R0);
and and3794(N6774,N6778,N6779);
and and3800(N6785,N6789,N6790);
and and3801(N6786,N6791,in1);
and and3802(N6787,in2,N6792);
and and3803(N6788,N6793,R3);
and and3809(N6799,N6803,N6804);
and and3810(N6800,N6805,N6806);
and and3811(N6801,N6807,R0);
and and3812(N6802,R1,N6808);
and and3818(N6813,N6817,N6818);
and and3819(N6814,N6819,in1);
and and3820(N6815,in2,N6820);
and and3821(N6816,R1,N6821);
and and3827(N6827,N6831,N6832);
and and3828(N6828,N6833,in1);
and and3829(N6829,N6834,R0);
and and3830(N6830,R1,N6835);
and and3836(N6841,N6845,N6846);
and and3837(N6842,N6847,N6848);
and and3838(N6843,in2,R0);
and and3839(N6844,R1,N6849);
and and3845(N6855,N6859,N6860);
and and3846(N6856,N6861,in1);
and and3847(N6857,N6862,R0);
and and3848(N6858,R1,N6863);
and and3854(N6869,N6873,N6874);
and and3855(N6870,in0,N6875);
and and3856(N6871,in2,R0);
and and3857(N6872,R1,R2);
and and3863(N6883,N6887,N6888);
and and3864(N6884,in0,in1);
and and3865(N6885,N6889,N6890);
and and3866(N6886,R2,R3);
and and3872(N6897,N6901,N6902);
and and3873(N6898,in1,in2);
and and3874(N6899,N6903,R1);
and and3875(N6900,R2,N6904);
and and3881(N6911,N6915,N6916);
and and3882(N6912,in0,N6917);
and and3883(N6913,in2,N6918);
and and3884(N6914,R1,R2);
and and3890(N6925,N6929,N6930);
and and3891(N6926,in0,in2);
and and3892(N6927,R0,N6931);
and and3893(N6928,N6932,N6933);
and and3899(N6939,N6943,N6944);
and and3900(N6940,in1,in2);
and and3901(N6941,N6945,N6946);
and and3902(N6942,N6947,R3);
and and3908(N6953,N6957,N6958);
and and3909(N6954,in0,in2);
and and3910(N6955,R0,N6959);
and and3911(N6956,R2,N6960);
and and3917(N6967,N6971,N6972);
and and3918(N6968,in0,in1);
and and3919(N6969,N6973,R0);
and and3920(N6970,N6974,N6975);
and and3926(N6981,N6985,N6986);
and and3927(N6982,N6987,in1);
and and3928(N6983,N6988,R0);
and and3929(N6984,N6989,R2);
and and3935(N6995,N6999,N7000);
and and3936(N6996,N7001,N7002);
and and3937(N6997,R0,R1);
and and3938(N6998,N7003,R3);
and and3944(N7009,N7013,N7014);
and and3945(N7010,in0,N7015);
and and3946(N7011,in2,N7016);
and and3947(N7012,R1,N7017);
and and3953(N7023,N7027,N7028);
and and3954(N7024,N7029,in1);
and and3955(N7025,R0,R1);
and and3956(N7026,N7030,N7031);
and and3962(N7037,N7041,N7042);
and and3963(N7038,in0,in1);
and and3964(N7039,N7043,N7044);
and and3965(N7040,R1,R2);
and and3971(N7051,N7055,N7056);
and and3972(N7052,in0,in1);
and and3973(N7053,N7057,N7058);
and and3974(N7054,R2,R3);
and and3980(N7065,N7069,N7070);
and and3981(N7066,in1,N7071);
and and3982(N7067,R0,R1);
and and3983(N7068,N7072,R3);
and and3989(N7079,N7083,N7084);
and and3990(N7080,N7085,N7086);
and and3991(N7081,in2,R0);
and and3992(N7082,R1,R2);
and and3998(N7093,N7097,N7098);
and and3999(N7094,N7099,in1);
and and4000(N7095,N7100,R0);
and and4001(N7096,R1,N7101);
and and4007(N7107,N7111,N7112);
and and4008(N7108,in1,N7113);
and and4009(N7109,R0,N7114);
and and4010(N7110,N7115,R3);
and and4016(N7121,N7125,N7126);
and and4017(N7122,N7127,in1);
and and4018(N7123,R0,R1);
and and4019(N7124,R2,R3);
and and4025(N7134,N7138,N7139);
and and4026(N7135,in0,N7140);
and and4027(N7136,R0,R1);
and and4028(N7137,R2,R3);
and and4034(N7147,N7151,N7152);
and and4035(N7148,in1,in2);
and and4036(N7149,R0,R1);
and and4037(N7150,R2,R3);
and and4043(N7160,N7164,N7165);
and and4044(N7161,in0,in1);
and and4045(N7162,R0,R1);
and and4046(N7163,R2,N7166);
and and4052(N7173,N7177,N7178);
and and4053(N7174,in1,in2);
and and4054(N7175,R0,R1);
and and4055(N7176,N7179,R3);
and and4061(N7186,N7190,N7191);
and and4062(N7187,in0,in1);
and and4063(N7188,R0,N7192);
and and4064(N7189,R2,R3);
and and4070(N7199,N7203,N7204);
and and4071(N7200,N7205,N7206);
and and4072(N7201,R0,R1);
and and4073(N7202,R2,R3);
and and4079(N7212,N7216,N7217);
and and4080(N7213,N7218,in2);
and and4081(N7214,N7219,R1);
and and4082(N7215,R2,R3);
and and4088(N7225,N7229,N7230);
and and4089(N7226,N7231,in2);
and and4090(N7227,N7232,R1);
and and4091(N7228,N7233,R3);
and and4097(N7238,N7242,N7243);
and and4098(N7239,in0,N7244);
and and4099(N7240,N7245,R0);
and and4100(N7241,R1,N7246);
and and4106(N7251,N7255,N7256);
and and4107(N7252,N7257,in2);
and and4108(N7253,R0,N7258);
and and4109(N7254,N7259,R3);
and and4115(N7264,N7268,N7269);
and and4116(N7265,in0,N7270);
and and4117(N7266,R0,N7271);
and and4118(N7267,N7272,R3);
and and4124(N7277,N7281,N7282);
and and4125(N7278,N7283,N7284);
and and4126(N7279,R0,R1);
and and4127(N7280,R2,N7285);
and and4133(N7290,N7294,N7295);
and and4134(N7291,N7296,N7297);
and and4135(N7292,in2,R0);
and and4136(N7293,R2,N7298);
and and4142(N7303,N7307,N7308);
and and4143(N7304,in1,N7309);
and and4144(N7305,N7310,R1);
and and4145(N7306,R2,R3);
and and4151(N7316,N7320,N7321);
and and4152(N7317,N7322,N7323);
and and4153(N7318,N7324,R0);
and and4154(N7319,R1,N7325);
and and4160(N7329,N7333,N7334);
and and4161(N7330,N7335,N7336);
and and4162(N7331,in2,R0);
and and4163(N7332,R1,N7337);
and and4169(N7342,N7346,N7347);
and and4170(N7343,N7348,in2);
and and4171(N7344,R0,N7349);
and and4172(N7345,R2,N7350);
and and4178(N7355,N7359,N7360);
and and4179(N7356,in1,N7361);
and and4180(N7357,R0,N7362);
and and4181(N7358,R2,N7363);
and and4187(N7368,N7372,N7373);
and and4188(N7369,in0,N7374);
and and4189(N7370,N7375,R0);
and and4190(N7371,N7376,R2);
and and4196(N7381,N7385,N7386);
and and4197(N7382,N7387,N7388);
and and4198(N7383,R0,R1);
and and4199(N7384,R2,N7389);
and and4205(N7394,N7398,N7399);
and and4206(N7395,N7400,N7401);
and and4207(N7396,in2,R0);
and and4208(N7397,R2,N7402);
and and4214(N7407,N7411,N7412);
and and4215(N7408,N7413,in1);
and and4216(N7409,N7414,R0);
and and4217(N7410,R2,N7415);
and and4223(N7420,N7424,N7425);
and and4224(N7421,in0,N7426);
and and4225(N7422,in2,N7427);
and and4226(N7423,R2,N7428);
and and4232(N7433,N7437,N7438);
and and4233(N7434,in1,in2);
and and4234(N7435,N7439,N7440);
and and4235(N7436,R2,N7441);
and and4241(N7446,N7450,N7451);
and and4242(N7447,N7452,N7453);
and and4243(N7448,R0,N7454);
and and4244(N7449,R2,R3);
and and4250(N7459,N7463,N7464);
and and4251(N7460,N7465,in1);
and and4252(N7461,in2,N7466);
and and4253(N7462,R2,R3);
and and4259(N7472,N7476,N7477);
and and4260(N7473,in0,N7478);
and and4261(N7474,N7479,N7480);
and and4262(N7475,R1,N7481);
and and4268(N7485,N7489,N7490);
and and4269(N7486,N7491,in1);
and and4270(N7487,N7492,R1);
and and4271(N7488,N7493,R3);
and and4277(N7498,N7502,N7503);
and and4278(N7499,N7504,in1);
and and4279(N7500,N7505,R1);
and and4280(N7501,R2,N7506);
and and4286(N7511,N7515,N7516);
and and4287(N7512,in0,N7517);
and and4288(N7513,N7518,R1);
and and4289(N7514,R2,N7519);
and and4295(N7524,N7528,N7529);
and and4296(N7525,N7530,in1);
and and4297(N7526,in2,R0);
and and4298(N7527,R1,R2);
and and4304(N7537,N7541,N7542);
and and4305(N7538,in0,in1);
and and4306(N7539,N7543,N7544);
and and4307(N7540,R2,R3);
and and4313(N7550,N7554,N7555);
and and4314(N7551,in0,in2);
and and4315(N7552,R0,N7556);
and and4316(N7553,N7557,R3);
and and4322(N7563,N7567,N7568);
and and4323(N7564,N7569,in2);
and and4324(N7565,R0,R1);
and and4325(N7566,N7570,R3);
and and4331(N7576,N7580,N7581);
and and4332(N7577,in0,in1);
and and4333(N7578,in2,R1);
and and4334(N7579,R2,N7582);
and and4340(N7589,N7593,N7594);
and and4341(N7590,N7595,in1);
and and4342(N7591,N7596,R0);
and and4343(N7592,R2,R3);
and and4349(N7602,N7606,N7607);
and and4350(N7603,N7608,in1);
and and4351(N7604,in2,R0);
and and4352(N7605,N7609,R3);
and and4358(N7615,N7619,N7620);
and and4359(N7616,in0,in1);
and and4360(N7617,in2,R1);
and and4361(N7618,R2,R3);
and and4367(N7627,N7631,N7632);
and and4368(N7628,N7633,in1);
and and4369(N7629,R0,R1);
and and4370(N7630,N7634,R3);
and and4376(N7639,N7643,N7644);
and and4377(N7640,N7645,in2);
and and4378(N7641,R0,R1);
and and4379(N7642,N7646,R3);
and and4385(N7651,N7655,N7656);
and and4386(N7652,in1,in2);
and and4387(N7653,R0,R1);
and and4388(N7654,N7657,R3);
and and4394(N7663,N7667,N7668);
and and4395(N7664,in0,in1);
and and4396(N7665,N7669,R0);
and and4397(N7666,R1,N7670);
and and4403(N7675,N7679,N7680);
and and4404(N7676,N7681,in1);
and and4405(N7677,N7682,R0);
and and4406(N7678,R1,R3);
and and4412(N7687,N7691,N7692);
and and4413(N7688,in1,in2);
and and4414(N7689,R0,N7693);
and and4415(N7690,R2,R3);
and and4421(N7699,N7703,N7704);
and and4422(N7700,N7705,in1);
and and4423(N7701,in2,N7706);
and and4424(N7702,R1,R2);
and and4430(N7711,N7715,N7716);
and and4431(N7712,N7717,in2);
and and4432(N7713,N7718,N7719);
and and4433(N7714,R2,R3);
and and4439(N7723,N7727,N7728);
and and4440(N7724,in0,in1);
and and4441(N7725,N7729,R1);
and and4442(N7726,N7730,R3);
and and4448(N7735,N7739,N7740);
and and4449(N7736,N7741,in1);
and and4450(N7737,in2,R1);
and and4451(N7738,N7742,R3);
and and4457(N7747,N7751,N7752);
and and4458(N7748,in0,N7753);
and and4459(N7749,N7754,R0);
and and4460(N7750,R2,R3);
and and4466(N7759,N7763,N7764);
and and4467(N7760,N7765,in1);
and and4468(N7761,N7766,R0);
and and4469(N7762,R1,R3);
and and4475(N7771,N7775,N7776);
and and4476(N7772,N7777,in1);
and and4477(N7773,in2,R0);
and and4478(N7774,R1,N7778);
and and4484(N7783,N7787,N7788);
and and4485(N7784,in0,N7789);
and and4486(N7785,R0,R1);
and and4487(N7786,R2,R3);
and and4493(N7795,N7799,N7800);
and and4494(N7796,in0,N7801);
and and4495(N7797,in2,R0);
and and4496(N7798,R1,N7802);
and and4502(N7807,N7811,N7812);
and and4503(N7808,in0,in1);
and and4504(N7809,R0,R1);
and and4505(N7810,N7813,R3);
and and4511(N7819,N7823,N7824);
and and4512(N7820,in1,N7825);
and and4513(N7821,N7826,R1);
and and4514(N7822,N7827,R3);
and and4520(N7831,N7835,N7836);
and and4521(N7832,N7837,N7838);
and and4522(N7833,N7839,R1);
and and4523(N7834,R2,R3);
and and4529(N7843,N7847,N7848);
and and4530(N7844,in0,in1);
and and4531(N7845,N7849,N7850);
and and4532(N7846,R1,R3);
and and4538(N7855,N7859,N7860);
and and4539(N7856,in0,in1);
and and4540(N7857,N7861,N7862);
and and4541(N7858,R1,R2);
and and4547(N7867,N7871,N7872);
and and4548(N7868,N7873,in1);
and and4549(N7869,in2,R0);
and and4550(N7870,R1,R2);
and and4556(N7879,N7883,N7884);
and and4557(N7880,in0,in1);
and and4558(N7881,in2,R0);
and and4559(N7882,R1,N7885);
and and4565(N7891,N7895,N7896);
and and4566(N7892,N7897,in1);
and and4567(N7893,in2,R0);
and and4568(N7894,N7898,R2);
and and4574(N7903,N7907,N7908);
and and4575(N7904,in0,N7909);
and and4576(N7905,R0,R1);
and and4577(N7906,N7910,R3);
and and4583(N7914,N7918,N7919);
and and4584(N7915,in0,in2);
and and4585(N7916,N7920,R1);
and and4586(N7917,R2,N7921);
and and4592(N7925,N7929,N7930);
and and4593(N7926,in0,in2);
and and4594(N7927,R0,R1);
and and4595(N7928,R2,R3);
and and4601(N7936,N7940,N7941);
and and4602(N7937,in0,in1);
and and4603(N7938,N7942,R0);
and and4604(N7939,R1,R2);
and and4610(N7947,N7951,N7952);
and and4611(N7948,in0,in1);
and and4612(N7949,in2,R0);
and and4613(N7950,N7953,R3);
and and4619(N7958,N7962,N7963);
and and4620(N7959,in0,in1);
and and4621(N7960,in2,R0);
and and4622(N7961,R1,R2);
and and4628(N7969,N7973,N7974);
and and4629(N7970,in0,in1);
and and4630(N7971,R0,N7975);
and and4631(N7972,R2,R3);
and and4637(N7980,N7984,N7985);
and and4638(N7981,in1,N7986);
and and4639(N7982,R0,R1);
and and4640(N7983,R2,R3);
and and4646(N7991,N7995,N7996);
and and4647(N7992,in1,in2);
and and4648(N7993,N7997,R1);
and and4649(N7994,R2,R3);
and and4655(N8002,N8006,N8007);
and and4656(N8003,in0,N8008);
and and4657(N8004,in2,R0);
and and4658(N8005,R1,R2);
and and4664(N8013,N8017,N8018);
and and4665(N8014,N8019,in1);
and and4666(N8015,in2,R0);
and and4667(N8016,N8020,R2);
and and4673(N8024,N8028,N8029);
and and4674(N8025,in0,in1);
and and4675(N8026,R0,R1);
and and4676(N8027,R2,N8030);
and and4682(N8035,N8039,N8040);
and and4683(N8036,in0,in1);
and and4684(N8037,in2,R0);
and and4685(N8038,R1,N8041);
and and4691(N8045,N8049,N8050);
and and4692(N8046,in0,in1);
and and4693(N8047,N8051,R0);
and and4694(N8048,R1,R3);
and and4700(N8055,N8059,N8060);
and and4701(N8056,in0,in1);
and and4702(N8057,R0,R1);
and and4703(N8058,R2,R3);
and and4709(N8065,N8069,N8070);
and and4710(N8066,N8071,in1);
and and4711(N8067,in2,R0);
and and4712(N8068,R1,R2);
and and4718(N8075,N8079,N8080);
and and4719(N8076,in0,in1);
and and4720(N8077,in2,R0);
and and4721(N8078,R1,R3);
and and4727(N8085,N8089,N8090);
and and4728(N8086,in0,N8091);
and and4729(N8087,in2,R1);
and and4730(N8088,R2,R3);
and and4736(N8095,N8099,N8100);
and and4737(N8096,in0,in1);
and and4738(N8097,in2,R0);
and and4739(N8098,N8101,R2);
and and4745(N8105,N8109,N8110);
and and4746(N8106,in0,in1);
and and4747(N8107,in2,R1);
and and4748(N8108,R2,R3);
and and4754(N8115,N8119,N8120);
and and4755(N8116,in0,in1);
and and4756(N8117,in2,R0);
and and4757(N8118,R1,R2);
and and4763(N8124,N8128,N8129);
and and4764(N8125,N8130,N8131);
and and4765(N8126,N8132,N8133);
and and4766(N8127,N8134,N8135);
and and4771(N8140,N8144,N8145);
and and4772(N8141,in1,N8146);
and and4773(N8142,N8147,N8148);
and and4774(N8143,N8149,N8150);
and and4779(N8156,N8160,N8161);
and and4780(N8157,N8162,N8163);
and and4781(N8158,N8164,N8165);
and and4782(N8159,R4,R5);
and and4787(N8171,N8175,N8176);
and and4788(N8172,N8177,N8178);
and and4789(N8173,N8179,N8180);
and and4790(N8174,R3,N8181);
and and4795(N8186,N8190,in0);
and and4796(N8187,in1,N8191);
and and4797(N8188,N8192,N8193);
and and4798(N8189,N8194,N8195);
and and4803(N8201,N8205,in1);
and and4804(N8202,in2,N8206);
and and4805(N8203,N8207,N8208);
and and4806(N8204,N8209,N8210);
and and4811(N8216,N8220,in1);
and and4812(N8217,N8221,N8222);
and and4813(N8218,N8223,N8224);
and and4814(N8219,N8225,N8226);
and and4819(N8231,N8235,N8236);
and and4820(N8232,N8237,N8238);
and and4821(N8233,R1,N8239);
and and4822(N8234,N8240,N8241);
and and4827(N8246,N8250,N8251);
and and4828(N8247,N8252,N8253);
and and4829(N8248,R1,N8254);
and and4830(N8249,N8255,R5);
and and4835(N8261,N8265,N8266);
and and4836(N8262,in2,N8267);
and and4837(N8263,N8268,N8269);
and and4838(N8264,N8270,R4);
and and4843(N8276,N8280,in0);
and and4844(N8277,N8281,N8282);
and and4845(N8278,N8283,R2);
and and4846(N8279,N8284,N8285);
and and4851(N8291,N8295,N8296);
and and4852(N8292,N8297,R0);
and and4853(N8293,N8298,N8299);
and and4854(N8294,N8300,N8301);
and and4859(N8306,N8310,N8311);
and and4860(N8307,N8312,R0);
and and4861(N8308,N8313,N8314);
and and4862(N8309,N8315,R4);
and and4867(N8321,N8325,in1);
and and4868(N8322,N8326,N8327);
and and4869(N8323,N8328,R3);
and and4870(N8324,N8329,N8330);
and and4875(N8336,N8340,in0);
and and4876(N8337,N8341,N8342);
and and4877(N8338,R0,N8343);
and and4878(N8339,N8344,N8345);
and and4883(N8351,N8355,in0);
and and4884(N8352,N8356,N8357);
and and4885(N8353,N8358,N8359);
and and4886(N8354,N8360,N8361);
and and4891(N8366,N8370,N8371);
and and4892(N8367,in2,N8372);
and and4893(N8368,N8373,R2);
and and4894(N8369,N8374,R5);
and and4899(N8380,N8384,in0);
and and4900(N8381,N8385,N8386);
and and4901(N8382,N8387,N8388);
and and4902(N8383,R3,N8389);
and and4907(N8394,N8398,in0);
and and4908(N8395,in2,N8399);
and and4909(N8396,N8400,N8401);
and and4910(N8397,N8402,N8403);
and and4915(N8408,N8412,in0);
and and4916(N8409,in1,N8413);
and and4917(N8410,N8414,N8415);
and and4918(N8411,N8416,N8417);
and and4923(N8422,N8426,in0);
and and4924(N8423,N8427,N8428);
and and4925(N8424,N8429,R2);
and and4926(N8425,R4,N8430);
and and4931(N8436,N8440,in0);
and and4932(N8437,N8441,N8442);
and and4933(N8438,N8443,R1);
and and4934(N8439,R2,N8444);
and and4939(N8450,N8454,N8455);
and and4940(N8451,N8456,N8457);
and and4941(N8452,R2,R3);
and and4942(N8453,N8458,N8459);
and and4947(N8464,N8468,N8469);
and and4948(N8465,N8470,R0);
and and4949(N8466,R1,N8471);
and and4950(N8467,N8472,N8473);
and and4955(N8478,N8482,N8483);
and and4956(N8479,N8484,N8485);
and and4957(N8480,R2,R3);
and and4958(N8481,N8486,R5);
and and4963(N8492,N8496,N8497);
and and4964(N8493,N8498,in2);
and and4965(N8494,N8499,R1);
and and4966(N8495,N8500,N8501);
and and4971(N8506,N8510,N8511);
and and4972(N8507,in1,N8512);
and and4973(N8508,R0,R3);
and and4974(N8509,N8513,N8514);
and and4979(N8520,N8524,N8525);
and and4980(N8521,in2,R0);
and and4981(N8522,N8526,R3);
and and4982(N8523,N8527,N8528);
and and4987(N8534,N8538,N8539);
and and4988(N8535,N8540,in2);
and and4989(N8536,R0,N8541);
and and4990(N8537,N8542,N8543);
and and4995(N8548,N8552,in0);
and and4996(N8549,N8553,N8554);
and and4997(N8550,N8555,N8556);
and and4998(N8551,R4,N8557);
and and5003(N8562,N8566,N8567);
and and5004(N8563,in1,N8568);
and and5005(N8564,N8569,N8570);
and and5006(N8565,R4,N8571);
and and5011(N8576,N8580,N8581);
and and5012(N8577,N8582,R0);
and and5013(N8578,N8583,N8584);
and and5014(N8579,R4,N8585);
and and5019(N8590,N8594,N8595);
and and5020(N8591,in2,R0);
and and5021(N8592,N8596,R2);
and and5022(N8593,N8597,N8598);
and and5027(N8604,N8608,N8609);
and and5028(N8605,in1,R0);
and and5029(N8606,R2,N8610);
and and5030(N8607,N8611,N8612);
and and5035(N8618,N8622,in0);
and and5036(N8619,N8623,R0);
and and5037(N8620,R2,N8624);
and and5038(N8621,N8625,N8626);
and and5043(N8632,N8636,N8637);
and and5044(N8633,R0,N8638);
and and5045(N8634,N8639,N8640);
and and5046(N8635,R4,R5);
and and5051(N8646,N8650,N8651);
and and5052(N8647,in1,N8652);
and and5053(N8648,N8653,R1);
and and5054(N8649,N8654,N8655);
and and5059(N8660,N8664,N8665);
and and5060(N8661,N8666,in2);
and and5061(N8662,N8667,R1);
and and5062(N8663,N8668,N8669);
and and5067(N8674,N8678,in0);
and and5068(N8675,N8679,N8680);
and and5069(N8676,N8681,N8682);
and and5070(N8677,R3,N8683);
and and5075(N8688,N8692,N8693);
and and5076(N8689,in2,N8694);
and and5077(N8690,N8695,R3);
and and5078(N8691,N8696,R5);
and and5083(N8702,N8706,in0);
and and5084(N8703,N8707,in2);
and and5085(N8704,N8708,N8709);
and and5086(N8705,R2,N8710);
and and5091(N8716,N8720,N8721);
and and5092(N8717,in1,R0);
and and5093(N8718,N8722,N8723);
and and5094(N8719,N8724,N8725);
and and5099(N8730,N8734,in0);
and and5100(N8731,N8735,N8736);
and and5101(N8732,R0,N8737);
and and5102(N8733,R4,N8738);
and and5107(N8744,N8748,N8749);
and and5108(N8745,N8750,N8751);
and and5109(N8746,R1,R2);
and and5110(N8747,N8752,N8753);
and and5115(N8758,N8762,in1);
and and5116(N8759,N8763,N8764);
and and5117(N8760,R1,N8765);
and and5118(N8761,N8766,N8767);
and and5123(N8772,N8776,N8777);
and and5124(N8773,N8778,in2);
and and5125(N8774,N8779,R1);
and and5126(N8775,N8780,N8781);
and and5131(N8786,N8790,N8791);
and and5132(N8787,N8792,R0);
and and5133(N8788,R1,N8793);
and and5134(N8789,N8794,N8795);
and and5139(N8800,N8804,in0);
and and5140(N8801,in1,R0);
and and5141(N8802,N8805,N8806);
and and5142(N8803,N8807,N8808);
and and5147(N8814,N8818,N8819);
and and5148(N8815,N8820,N8821);
and and5149(N8816,N8822,R2);
and and5150(N8817,N8823,R4);
and and5155(N8828,N8832,N8833);
and and5156(N8829,N8834,R1);
and and5157(N8830,R2,N8835);
and and5158(N8831,N8836,R5);
and and5163(N8842,N8846,N8847);
and and5164(N8843,in1,R0);
and and5165(N8844,N8848,R3);
and and5166(N8845,N8849,N8850);
and and5171(N8856,N8860,in0);
and and5172(N8857,N8861,N8862);
and and5173(N8858,N8863,R2);
and and5174(N8859,R4,N8864);
and and5179(N8870,N8874,in0);
and and5180(N8871,in1,N8875);
and and5181(N8872,N8876,R2);
and and5182(N8873,N8877,N8878);
and and5187(N8884,N8888,in0);
and and5188(N8885,N8889,N8890);
and and5189(N8886,N8891,R1);
and and5190(N8887,N8892,N8893);
and and5195(N8898,N8902,in0);
and and5196(N8899,in1,in2);
and and5197(N8900,N8903,R1);
and and5198(N8901,N8904,N8905);
and and5203(N8911,N8915,N8916);
and and5204(N8912,N8917,R1);
and and5205(N8913,N8918,R3);
and and5206(N8914,N8919,N8920);
and and5211(N8924,N8928,in0);
and and5212(N8925,N8929,N8930);
and and5213(N8926,R1,N8931);
and and5214(N8927,R3,R5);
and and5219(N8937,N8941,N8942);
and and5220(N8938,R0,R1);
and and5221(N8939,N8943,N8944);
and and5222(N8940,R4,N8945);
and and5227(N8950,N8954,in0);
and and5228(N8951,N8955,in2);
and and5229(N8952,N8956,R3);
and and5230(N8953,R4,N8957);
and and5235(N8963,N8967,in0);
and and5236(N8964,in1,N8968);
and and5237(N8965,N8969,R3);
and and5238(N8966,R4,N8970);
and and5243(N8976,N8980,in0);
and and5244(N8977,N8981,N8982);
and and5245(N8978,N8983,R3);
and and5246(N8979,R4,R5);
and and5251(N8989,N8993,N8994);
and and5252(N8990,N8995,in2);
and and5253(N8991,R0,N8996);
and and5254(N8992,R3,N8997);
and and5259(N9002,N9006,in0);
and and5260(N9003,N9007,N9008);
and and5261(N9004,R1,N9009);
and and5262(N9005,N9010,N9011);
and and5267(N9015,N9019,in0);
and and5268(N9016,in1,R0);
and and5269(N9017,N9020,R3);
and and5270(N9018,N9021,N9022);
and and5275(N9028,N9032,N9033);
and and5276(N9029,N9034,R1);
and and5277(N9030,N9035,N9036);
and and5278(N9031,R4,R5);
and and5283(N9041,N9045,N9046);
and and5284(N9042,in1,in2);
and and5285(N9043,R0,N9047);
and and5286(N9044,N9048,N9049);
and and5291(N9054,N9058,in0);
and and5292(N9055,in2,R0);
and and5293(N9056,N9059,N9060);
and and5294(N9057,N9061,N9062);
and and5299(N9067,N9071,in0);
and and5300(N9068,in1,R0);
and and5301(N9069,N9072,N9073);
and and5302(N9070,N9074,N9075);
and and5307(N9080,N9084,N9085);
and and5308(N9081,N9086,R0);
and and5309(N9082,R2,N9087);
and and5310(N9083,N9088,N9089);
and and5315(N9093,N9097,N9098);
and and5316(N9094,N9099,N9100);
and and5317(N9095,R1,R3);
and and5318(N9096,N9101,R5);
and and5323(N9106,N9110,in0);
and and5324(N9107,N9111,N9112);
and and5325(N9108,R2,N9113);
and and5326(N9109,N9114,R5);
and and5331(N9119,N9123,in1);
and and5332(N9120,in2,N9124);
and and5333(N9121,N9125,R2);
and and5334(N9122,N9126,N9127);
and and5339(N9132,N9136,in0);
and and5340(N9133,N9137,R0);
and and5341(N9134,N9138,N9139);
and and5342(N9135,R4,N9140);
and and5347(N9145,N9149,in1);
and and5348(N9146,N9150,N9151);
and and5349(N9147,N9152,R3);
and and5350(N9148,R4,N9153);
and and5355(N9158,N9162,N9163);
and and5356(N9159,in2,N9164);
and and5357(N9160,N9165,R3);
and and5358(N9161,R4,N9166);
and and5363(N9171,N9175,in0);
and and5364(N9172,N9176,N9177);
and and5365(N9173,R1,N9178);
and and5366(N9174,N9179,R5);
and and5371(N9184,N9188,in1);
and and5372(N9185,in2,N9189);
and and5373(N9186,R1,N9190);
and and5374(N9187,N9191,R5);
and and5379(N9197,N9201,in0);
and and5380(N9198,N9202,in2);
and and5381(N9199,N9203,R1);
and and5382(N9200,N9204,R5);
and and5387(N9210,N9214,in0);
and and5388(N9211,in1,N9215);
and and5389(N9212,N9216,R1);
and and5390(N9213,N9217,R5);
and and5395(N9223,N9227,N9228);
and and5396(N9224,in1,in2);
and and5397(N9225,N9229,N9230);
and and5398(N9226,R3,N9231);
and and5403(N9236,N9240,N9241);
and and5404(N9237,N9242,R0);
and and5405(N9238,R1,N9243);
and and5406(N9239,N9244,R4);
and and5411(N9249,N9253,in0);
and and5412(N9250,in2,R1);
and and5413(N9251,N9254,N9255);
and and5414(N9252,R4,N9256);
and and5419(N9262,N9266,in0);
and and5420(N9263,in1,R1);
and and5421(N9264,N9267,N9268);
and and5422(N9265,R4,N9269);
and and5427(N9275,N9279,N9280);
and and5428(N9276,N9281,N9282);
and and5429(N9277,R1,R3);
and and5430(N9278,R4,N9283);
and and5435(N9288,N9292,N9293);
and and5436(N9289,in2,N9294);
and and5437(N9290,N9295,R3);
and and5438(N9291,N9296,R5);
and and5443(N9301,N9305,in0);
and and5444(N9302,in2,R0);
and and5445(N9303,N9306,N9307);
and and5446(N9304,N9308,N9309);
and and5451(N9314,N9318,in0);
and and5452(N9315,in1,R0);
and and5453(N9316,N9319,N9320);
and and5454(N9317,N9321,N9322);
and and5459(N9327,N9331,N9332);
and and5460(N9328,N9333,R0);
and and5461(N9329,R1,N9334);
and and5462(N9330,N9335,N9336);
and and5467(N9340,N9344,N9345);
and and5468(N9341,N9346,R1);
and and5469(N9342,N9347,N9348);
and and5470(N9343,R4,R5);
and and5475(N9353,N9357,N9358);
and and5476(N9354,in1,in2);
and and5477(N9355,R0,N9359);
and and5478(N9356,N9360,R4);
and and5483(N9366,N9370,in0);
and and5484(N9367,in2,R0);
and and5485(N9368,N9371,N9372);
and and5486(N9369,N9373,R4);
and and5491(N9379,N9383,in0);
and and5492(N9380,in1,R0);
and and5493(N9381,N9384,N9385);
and and5494(N9382,N9386,R4);
and and5499(N9392,N9396,N9397);
and and5500(N9393,in1,N9398);
and and5501(N9394,N9399,R1);
and and5502(N9395,R2,N9400);
and and5507(N9405,N9409,N9410);
and and5508(N9406,in1,N9411);
and and5509(N9407,N9412,R2);
and and5510(N9408,R3,N9413);
and and5515(N9418,N9422,in0);
and and5516(N9419,N9423,N9424);
and and5517(N9420,N9425,R2);
and and5518(N9421,R3,N9426);
and and5523(N9431,N9435,N9436);
and and5524(N9432,N9437,R0);
and and5525(N9433,R1,R3);
and and5526(N9434,N9438,R5);
and and5531(N9444,N9448,N9449);
and and5532(N9445,in1,R0);
and and5533(N9446,N9450,R2);
and and5534(N9447,N9451,N9452);
and and5539(N9457,N9461,N9462);
and and5540(N9458,N9463,in2);
and and5541(N9459,R0,R1);
and and5542(N9460,N9464,N9465);
and and5547(N9470,N9474,N9475);
and and5548(N9471,N9476,R1);
and and5549(N9472,R2,N9477);
and and5550(N9473,R4,N9478);
and and5555(N9483,N9487,N9488);
and and5556(N9484,R0,N9489);
and and5557(N9485,N9490,R3);
and and5558(N9486,R4,R5);
and and5563(N9496,N9500,N9501);
and and5564(N9497,N9502,N9503);
and and5565(N9498,N9504,R2);
and and5566(N9499,R3,R4);
and and5571(N9509,N9513,in0);
and and5572(N9510,N9514,in2);
and and5573(N9511,R2,R3);
and and5574(N9512,N9515,N9516);
and and5579(N9522,N9526,in0);
and and5580(N9523,in1,N9527);
and and5581(N9524,N9528,R2);
and and5582(N9525,R4,N9529);
and and5587(N9535,N9539,N9540);
and and5588(N9536,N9541,in2);
and and5589(N9537,N9542,R1);
and and5590(N9538,R2,N9543);
and and5595(N9548,N9552,in1);
and and5596(N9549,in2,R0);
and and5597(N9550,R2,N9553);
and and5598(N9551,N9554,N9555);
and and5603(N9561,N9565,N9566);
and and5604(N9562,in1,N9567);
and and5605(N9563,N9568,N9569);
and and5606(N9564,R3,R4);
and and5611(N9574,N9578,in0);
and and5612(N9575,in1,N9579);
and and5613(N9576,N9580,R3);
and and5614(N9577,R4,N9581);
and and5619(N9587,N9591,in0);
and and5620(N9588,N9592,in2);
and and5621(N9589,R1,N9593);
and and5622(N9590,N9594,R4);
and and5627(N9600,N9604,N9605);
and and5628(N9601,in2,N9606);
and and5629(N9602,R1,N9607);
and and5630(N9603,N9608,R4);
and and5635(N9613,N9617,in0);
and and5636(N9614,N9618,N9619);
and and5637(N9615,R0,R1);
and and5638(N9616,N9620,N9621);
and and5643(N9626,N9630,N9631);
and and5644(N9627,N9632,in2);
and and5645(N9628,R0,N9633);
and and5646(N9629,N9634,R3);
and and5651(N9639,N9643,in0);
and and5652(N9640,R0,N9644);
and and5653(N9641,R2,N9645);
and and5654(N9642,R4,N9646);
and and5659(N9651,N9655,N9656);
and and5660(N9652,N9657,R0);
and and5661(N9653,N9658,R2);
and and5662(N9654,R3,R5);
and and5667(N9663,N9667,in0);
and and5668(N9664,in1,R0);
and and5669(N9665,R1,N9668);
and and5670(N9666,N9669,N9670);
and and5675(N9675,N9679,N9680);
and and5676(N9676,in2,N9681);
and and5677(N9677,N9682,R2);
and and5678(N9678,R3,R5);
and and5683(N9687,N9691,N9692);
and and5684(N9688,N9693,N9694);
and and5685(N9689,R1,R2);
and and5686(N9690,R3,R4);
and and5691(N9699,N9703,N9704);
and and5692(N9700,N9705,R0);
and and5693(N9701,R1,R2);
and and5694(N9702,R3,N9706);
and and5699(N9711,N9715,in0);
and and5700(N9712,N9716,R1);
and and5701(N9713,R2,N9717);
and and5702(N9714,N9718,R5);
and and5707(N9723,N9727,in0);
and and5708(N9724,in2,N9728);
and and5709(N9725,N9729,R3);
and and5710(N9726,N9730,R5);
and and5715(N9735,N9739,in0);
and and5716(N9736,in1,N9740);
and and5717(N9737,N9741,R3);
and and5718(N9738,N9742,R5);
and and5723(N9747,N9751,in1);
and and5724(N9748,N9752,R0);
and and5725(N9749,N9753,R3);
and and5726(N9750,N9754,N9755);
and and5731(N9759,N9763,N9764);
and and5732(N9760,in2,N9765);
and and5733(N9761,N9766,R2);
and and5734(N9762,R3,R4);
and and5739(N9771,N9775,N9776);
and and5740(N9772,in1,N9777);
and and5741(N9773,R1,R3);
and and5742(N9774,N9778,R5);
and and5747(N9783,N9787,N9788);
and and5748(N9784,N9789,R1);
and and5749(N9785,N9790,R3);
and and5750(N9786,N9791,R5);
and and5755(N9795,N9799,in1);
and and5756(N9796,in2,N9800);
and and5757(N9797,R1,N9801);
and and5758(N9798,N9802,R5);
and and5763(N9807,N9811,in0);
and and5764(N9808,N9812,in2);
and and5765(N9809,R1,N9813);
and and5766(N9810,N9814,R5);
and and5771(N9819,N9823,in1);
and and5772(N9820,in2,R0);
and and5773(N9821,N9824,N9825);
and and5774(N9822,R4,R5);
and and5779(N9831,N9835,N9836);
and and5780(N9832,in2,N9837);
and and5781(N9833,N9838,R3);
and and5782(N9834,R4,N9839);
and and5787(N9843,N9847,N9848);
and and5788(N9844,in2,R0);
and and5789(N9845,R1,N9849);
and and5790(N9846,N9850,R4);
and and5795(N9855,N9859,in0);
and and5796(N9856,N9860,in2);
and and5797(N9857,R0,N9861);
and and5798(N9858,R3,R4);
and and5803(N9867,N9871,N9872);
and and5804(N9868,N9873,R0);
and and5805(N9869,R1,R2);
and and5806(N9870,N9874,R4);
and and5811(N9879,N9883,N9884);
and and5812(N9880,N9885,R1);
and and5813(N9881,R2,R3);
and and5814(N9882,R4,N9886);
and and5819(N9891,N9895,in1);
and and5820(N9892,N9896,N9897);
and and5821(N9893,R2,N9898);
and and5822(N9894,R4,N9899);
and and5827(N9903,N9907,in0);
and and5828(N9904,N9908,N9909);
and and5829(N9905,R2,R3);
and and5830(N9906,N9910,N9911);
and and5835(N9915,N9919,in0);
and and5836(N9916,in2,N9920);
and and5837(N9917,R1,R2);
and and5838(N9918,N9921,N9922);
and and5843(N9927,N9931,in1);
and and5844(N9928,in2,N9932);
and and5845(N9929,R1,R2);
and and5846(N9930,N9933,N9934);
and and5851(N9939,N9943,in0);
and and5852(N9940,N9944,R0);
and and5853(N9941,N9945,R2);
and and5854(N9942,R3,N9946);
and and5859(N9951,N9955,in1);
and and5860(N9952,R0,N9956);
and and5861(N9953,R2,R3);
and and5862(N9954,N9957,N9958);
and and5867(N9963,N9967,in0);
and and5868(N9964,in2,R0);
and and5869(N9965,R1,N9968);
and and5870(N9966,N9969,N9970);
and and5875(N9975,N9979,N9980);
and and5876(N9976,in1,R0);
and and5877(N9977,N9981,R2);
and and5878(N9978,N9982,R4);
and and5883(N9987,N9991,in0);
and and5884(N9988,N9992,R0);
and and5885(N9989,N9993,R2);
and and5886(N9990,N9994,R4);
and and5891(N9999,N10003,N10004);
and and5892(N10000,in2,R0);
and and5893(N10001,R1,R2);
and and5894(N10002,N10005,N10006);
and and5899(N10011,N10015,in0);
and and5900(N10012,N10016,N10017);
and and5901(N10013,N10018,R1);
and and5902(N10014,R2,N10019);
and and5907(N10023,N10027,in0);
and and5908(N10024,N10028,R0);
and and5909(N10025,N10029,R2);
and and5910(N10026,N10030,R4);
and and5915(N10035,N10039,in1);
and and5916(N10036,in2,N10040);
and and5917(N10037,N10041,R2);
and and5918(N10038,N10042,R4);
and and5923(N10047,N10051,in0);
and and5924(N10048,N10052,in2);
and and5925(N10049,N10053,R2);
and and5926(N10050,N10054,R4);
and and5931(N10059,N10063,in0);
and and5932(N10060,in1,N10064);
and and5933(N10061,N10065,R2);
and and5934(N10062,N10066,R4);
and and5939(N10071,N10075,in0);
and and5940(N10072,N10076,N10077);
and and5941(N10073,R0,N10078);
and and5942(N10074,R3,R4);
and and5947(N10083,N10087,in0);
and and5948(N10084,N10088,N10089);
and and5949(N10085,R2,R3);
and and5950(N10086,R4,N10090);
and and5955(N10095,N10099,in2);
and and5956(N10096,N10100,R1);
and and5957(N10097,N10101,N10102);
and and5958(N10098,R4,R5);
and and5963(N10107,N10111,in0);
and and5964(N10108,in1,in2);
and and5965(N10109,N10112,N10113);
and and5966(N10110,R3,N10114);
and and5971(N10119,N10123,in0);
and and5972(N10120,N10124,R0);
and and5973(N10121,R2,N10125);
and and5974(N10122,N10126,N10127);
and and5979(N10131,N10135,in0);
and and5980(N10132,N10136,R0);
and and5981(N10133,R2,N10137);
and and5982(N10134,N10138,N10139);
and and5987(N10143,N10147,in0);
and and5988(N10144,N10148,R0);
and and5989(N10145,R2,N10149);
and and5990(N10146,R4,N10150);
and and5995(N10155,N10159,in0);
and and5996(N10156,in1,in2);
and and5997(N10157,N10160,R1);
and and5998(N10158,N10161,N10162);
and and6003(N10167,N10171,in1);
and and6004(N10168,in2,N10172);
and and6005(N10169,N10173,R2);
and and6006(N10170,R3,N10174);
and and6011(N10179,N10183,in0);
and and6012(N10180,N10184,R0);
and and6013(N10181,R1,R2);
and and6014(N10182,N10185,R5);
and and6019(N10191,N10195,N10196);
and and6020(N10192,in1,in2);
and and6021(N10193,N10197,N10198);
and and6022(N10194,R2,R3);
and and6027(N10203,N10207,in0);
and and6028(N10204,in1,N10208);
and and6029(N10205,R0,R1);
and and6030(N10206,R2,R3);
and and6035(N10214,N10218,N10219);
and and6036(N10215,in2,N10220);
and and6037(N10216,R1,R2);
and and6038(N10217,R3,R5);
and and6043(N10225,N10229,in0);
and and6044(N10226,in1,in2);
and and6045(N10227,R1,N10230);
and and6046(N10228,R3,R5);
and and6051(N10236,N10240,in0);
and and6052(N10237,N10241,R1);
and and6053(N10238,N10242,R3);
and and6054(N10239,R4,N10243);
and and6059(N10247,N10251,in1);
and and6060(N10248,in2,R0);
and and6061(N10249,R1,N10252);
and and6062(N10250,R3,N10253);
and and6067(N10258,N10262,in0);
and and6068(N10259,in1,N10263);
and and6069(N10260,R0,R1);
and and6070(N10261,N10264,R3);
and and6075(N10269,N10273,N10274);
and and6076(N10270,in1,N10275);
and and6077(N10271,N10276,R2);
and and6078(N10272,R3,R4);
and and6083(N10280,N10284,in0);
and and6084(N10281,in1,N10285);
and and6085(N10282,R1,R2);
and and6086(N10283,R3,N10286);
and and6091(N10291,N10295,in0);
and and6092(N10292,R0,N10296);
and and6093(N10293,N10297,R3);
and and6094(N10294,R4,R5);
and and6099(N10302,N10306,in0);
and and6100(N10303,in2,N10307);
and and6101(N10304,R1,R2);
and and6102(N10305,R3,R5);
and and6107(N10313,N10317,N10318);
and and6108(N10314,in1,in2);
and and6109(N10315,R1,R2);
and and6110(N10316,N10319,R5);
and and6115(N10324,N10328,in0);
and and6116(N10325,in2,N10329);
and and6117(N10326,R1,N10330);
and and6118(N10327,R3,R5);
and and6123(N10335,N10339,in0);
and and6124(N10336,in1,in2);
and and6125(N10337,R0,N10340);
and and6126(N10338,N10341,R3);
and and6131(N10346,N10350,in1);
and and6132(N10347,R0,N10351);
and and6133(N10348,R2,R3);
and and6134(N10349,R4,N10352);
and and6139(N10357,N10361,N10362);
and and6140(N10358,in1,R0);
and and6141(N10359,R1,R2);
and and6142(N10360,R4,N10363);
and and6147(N10368,N10372,N10373);
and and6148(N10369,in2,N10374);
and and6149(N10370,R1,R2);
and and6150(N10371,R3,R4);
and and6155(N10379,N10383,in1);
and and6156(N10380,in2,N10384);
and and6157(N10381,R1,R3);
and and6158(N10382,R4,N10385);
and and6163(N10390,N10394,in0);
and and6164(N10391,in2,N10395);
and and6165(N10392,R1,R3);
and and6166(N10393,R4,N10396);
and and6171(N10401,N10405,in0);
and and6172(N10402,in1,in2);
and and6173(N10403,N10406,R1);
and and6174(N10404,N10407,R4);
and and6179(N10412,N10416,N10417);
and and6180(N10413,N10418,R1);
and and6181(N10414,R2,R3);
and and6182(N10415,N10419,R5);
and and6187(N10423,N10427,in0);
and and6188(N10424,in2,R0);
and and6189(N10425,R1,N10428);
and and6190(N10426,N10429,N10430);
and and6195(N10434,N10438,in0);
and and6196(N10435,in1,R0);
and and6197(N10436,R1,N10439);
and and6198(N10437,N10440,N10441);
and and6203(N10445,N10449,in1);
and and6204(N10446,in2,R1);
and and6205(N10447,N10450,N10451);
and and6206(N10448,R4,R5);
and and6211(N10456,N10460,in0);
and and6212(N10457,in2,R1);
and and6213(N10458,N10461,N10462);
and and6214(N10459,R4,R5);
and and6219(N10467,N10471,in0);
and and6220(N10468,in1,R1);
and and6221(N10469,N10472,N10473);
and and6222(N10470,R4,R5);
and and6227(N10478,N10482,in0);
and and6228(N10479,N10483,N10484);
and and6229(N10480,R1,R3);
and and6230(N10481,R4,R5);
and and6235(N10489,N10493,N10494);
and and6236(N10490,in2,N10495);
and and6237(N10491,R1,R3);
and and6238(N10492,R4,R5);
and and6243(N10500,N10504,in0);
and and6244(N10501,in2,R0);
and and6245(N10502,R1,N10505);
and and6246(N10503,R3,R5);
and and6251(N10511,N10515,in0);
and and6252(N10512,in2,N10516);
and and6253(N10513,R1,R2);
and and6254(N10514,N10517,R4);
and and6259(N10522,N10526,in0);
and and6260(N10523,N10527,R0);
and and6261(N10524,R1,R2);
and and6262(N10525,R4,R5);
and and6267(N10533,N10537,in0);
and and6268(N10534,N10538,in2);
and and6269(N10535,R0,R1);
and and6270(N10536,N10539,R4);
and and6275(N10544,N10548,in0);
and and6276(N10545,in1,N10549);
and and6277(N10546,R0,R1);
and and6278(N10547,R4,R5);
and and6283(N10555,N10559,in0);
and and6284(N10556,N10560,R0);
and and6285(N10557,N10561,R2);
and and6286(N10558,R3,R4);
and and6291(N10566,N10570,in1);
and and6292(N10567,in2,N10571);
and and6293(N10568,N10572,R2);
and and6294(N10569,R3,R5);
and and6299(N10577,N10581,in0);
and and6300(N10578,in2,R0);
and and6301(N10579,R1,N10582);
and and6302(N10580,N10583,R5);
and and6307(N10588,N10592,N10593);
and and6308(N10589,in1,in2);
and and6309(N10590,R0,R1);
and and6310(N10591,N10594,R4);
and and6315(N10599,N10603,in0);
and and6316(N10600,in1,R0);
and and6317(N10601,N10604,R2);
and and6318(N10602,N10605,R4);
and and6323(N10610,N10614,N10615);
and and6324(N10611,in2,N10616);
and and6325(N10612,R1,R2);
and and6326(N10613,R3,N10617);
and and6331(N10621,N10625,N10626);
and and6332(N10622,in2,N10627);
and and6333(N10623,R1,N10628);
and and6334(N10624,R3,R5);
and and6339(N10632,N10636,in0);
and and6340(N10633,in1,N10637);
and and6341(N10634,N10638,R1);
and and6342(N10635,R3,R5);
and and6347(N10643,N10647,N10648);
and and6348(N10644,in1,in2);
and and6349(N10645,R1,N10649);
and and6350(N10646,R4,R5);
and and6355(N10654,N10658,in0);
and and6356(N10655,in1,N10659);
and and6357(N10656,R0,R1);
and and6358(N10657,N10660,R3);
and and6363(N10665,N10669,in0);
and and6364(N10666,in2,N10670);
and and6365(N10667,R1,R2);
and and6366(N10668,R3,N10671);
and and6371(N10676,N10680,in0);
and and6372(N10677,in1,in2);
and and6373(N10678,R0,R1);
and and6374(N10679,R4,N10681);
and and6379(N10686,N10690,in1);
and and6380(N10687,in2,R0);
and and6381(N10688,R1,R2);
and and6382(N10689,N10691,N10692);
and and6387(N10696,N10700,in0);
and and6388(N10697,in1,R0);
and and6389(N10698,R2,N10701);
and and6390(N10699,R4,R5);
and and6395(N10706,N10710,in0);
and and6396(N10707,N10711,in2);
and and6397(N10708,R0,R3);
and and6398(N10709,R4,N10712);
and and6403(N10716,N10720,in0);
and and6404(N10717,in1,N10721);
and and6405(N10718,R0,R3);
and and6406(N10719,R4,N10722);
and and6411(N10726,N10730,in0);
and and6412(N10727,N10731,R0);
and and6413(N10728,R1,R2);
and and6414(N10729,R3,R4);
and and6419(N10736,N10740,in0);
and and6420(N10737,in2,R0);
and and6421(N10738,R1,R2);
and and6422(N10739,R3,N10741);
and and6427(N10746,N10750,in0);
and and6428(N10747,N10751,N10752);
and and6429(N10748,R2,R3);
and and6430(N10749,R4,R5);
and and6435(N10756,N10760,in0);
and and6436(N10757,in1,in2);
and and6437(N10758,R0,N10761);
and and6438(N10759,R2,N10762);
and and6443(N10766,N10770,N10771);
and and6444(N10767,in2,R0);
and and6445(N10768,R1,R2);
and and6446(N10769,R3,R5);
and and6451(N10776,N10780,in0);
and and6452(N10777,in1,in2);
and and6453(N10778,R0,R1);
and and6454(N10779,N10781,R4);
and and6459(N10786,N10790,in0);
and and6460(N10787,N10791,in2);
and and6461(N10788,R0,R1);
and and6462(N10789,R2,N10792);
and and6467(N10796,N10800,in0);
and and6468(N10797,N10801,N10802);
and and6469(N10798,R1,R2);
and and6470(N10799,R3,R4);
and and6475(N10806,N10810,in1);
and and6476(N10807,N10811,N10812);
and and6477(N10808,R1,R2);
and and6478(N10809,R3,R4);
and and6483(N10816,N10820,in0);
and and6484(N10817,N10821,in2);
and and6485(N10818,R0,R2);
and and6486(N10819,R3,R4);
and and6491(N10826,N10830,in0);
and and6492(N10827,N10831,R0);
and and6493(N10828,R1,R2);
and and6494(N10829,N10832,R4);
and and6499(N10836,N10840,N10841);
and and6500(N10837,in1,R0);
and and6501(N10838,R1,R2);
and and6502(N10839,N10842,R4);
and and6507(N10846,N10850,N10851);
and and6508(N10847,in2,R0);
and and6509(N10848,R1,R2);
and and6510(N10849,N10852,R4);
and and6515(N10856,N10860,in0);
and and6516(N10857,N10861,in2);
and and6517(N10858,R0,N10862);
and and6518(N10859,R2,R3);
and and6523(N10866,N10870,in0);
and and6524(N10867,N10871,N10872);
and and6525(N10868,R0,R1);
and and6526(N10869,R2,R3);
and and6531(N10876,N10880,in0);
and and6532(N10877,in1,N10881);
and and6533(N10878,R0,R1);
and and6534(N10879,R2,R3);
and and6539(N10886,N10890,in0);
and and6540(N10887,in1,in2);
and and6541(N10888,N10891,R1);
and and6542(N10889,R2,R4);
and and6547(N10896,N10900,in0);
and and6548(N10897,in1,in2);
and and6549(N10898,R1,N10901);
and and6550(N10899,R4,R5);
and and6555(N10906,N10910,in0);
and and6556(N10907,in1,in2);
and and6557(N10908,R0,R1);
and and6558(N10909,N10911,N10912);
and and6563(N10916,N10920,in0);
and and6564(N10917,in2,R0);
and and6565(N10918,R2,R3);
and and6566(N10919,R4,R5);
and and6571(N10926,N10930,in0);
and and6572(N10927,in1,in2);
and and6573(N10928,N10931,R1);
and and6574(N10929,R2,R3);
and and6579(N10935,N10939,in1);
and and6580(N10936,in2,N10940);
and and6581(N10937,R2,R3);
and and6582(N10938,R4,R5);
and and6587(N10944,N10948,in0);
and and6588(N10945,in1,R0);
and and6589(N10946,R1,R2);
and and6590(N10947,N10949,R5);
and and6595(N10953,N10957,in1);
and and6596(N10954,in2,R0);
and and6597(N10955,R1,R2);
and and6598(N10956,N10958,R5);
and and6603(N10962,N10966,in0);
and and6604(N10963,in1,in2);
and and6605(N10964,R1,N10967);
and and6606(N10965,R3,R4);
and and6611(N10971,N10975,N10976);
and and6612(N10972,N10977,R3);
and and6613(N10973,R4,N10978);
and and6614(N10974,N10979,N10980);
and and6618(N10984,in0,N10988);
and and6619(N10985,N10989,N10990);
and and6620(N10986,N10991,R4);
and and6621(N10987,N10992,N10993);
and and6625(N10997,in2,R0);
and and6626(N10998,N11001,N11002);
and and6627(N10999,N11003,N11004);
and and6628(N11000,N11005,N11006);
and and6632(N11010,in1,N11014);
and and6633(N11011,N11015,R1);
and and6634(N11012,R2,N11016);
and and6635(N11013,N11017,N11018);
and and6639(N11022,N11026,N11027);
and and6640(N11023,R2,N11028);
and and6641(N11024,R4,R5);
and and6642(N11025,N11029,N11030);
and and6646(N11034,in1,N11038);
and and6647(N11035,R2,N11039);
and and6648(N11036,N11040,N11041);
and and6649(N11037,N11042,R7);
and and6653(N11046,in1,R0);
and and6654(N11047,R1,N11050);
and and6655(N11048,N11051,N11052);
and and6656(N11049,N11053,N11054);
and and6660(N11058,in0,R0);
and and6661(N11059,R1,N11062);
and and6662(N11060,N11063,N11064);
and and6663(N11061,N11065,N11066);
and and6667(N11070,in0,N11074);
and and6668(N11071,N11075,R2);
and and6669(N11072,N11076,N11077);
and and6670(N11073,R6,N11078);
and and6674(N11082,in0,N11086);
and and6675(N11083,N11087,N11088);
and and6676(N11084,R1,N11089);
and and6677(N11085,N11090,R7);
and and6681(N11094,N11098,N11099);
and and6682(N11095,R0,N11100);
and and6683(N11096,R2,N11101);
and and6684(N11097,R5,N11102);
and and6688(N11106,N11110,N11111);
and and6689(N11107,N11112,R0);
and and6690(N11108,N11113,R2);
and and6691(N11109,R5,N11114);
and and6695(N11118,in0,in1);
and and6696(N11119,N11122,R3);
and and6697(N11120,N11123,N11124);
and and6698(N11121,R6,N11125);
and and6702(N11129,N11133,R0);
and and6703(N11130,R1,N11134);
and and6704(N11131,N11135,R5);
and and6705(N11132,N11136,R7);
and and6709(N11140,in0,in1);
and and6710(N11141,R1,N11144);
and and6711(N11142,N11145,N11146);
and and6712(N11143,R6,N11147);
and and6716(N11151,N11155,R0);
and and6717(N11152,N11156,R3);
and and6718(N11153,N11157,N11158);
and and6719(N11154,R6,R7);
and and6723(N11162,in1,N11166);
and and6724(N11163,R2,N11167);
and and6725(N11164,N11168,R5);
and and6726(N11165,N11169,R7);
and and6730(N11173,in0,in1);
and and6731(N11174,N11177,N11178);
and and6732(N11175,R3,N11179);
and and6733(N11176,R5,N11180);
and and6737(N11184,in0,N11188);
and and6738(N11185,N11189,R3);
and and6739(N11186,N11190,R5);
and and6740(N11187,R6,N11191);
and and6744(N11195,in0,N11199);
and and6745(N11196,N11200,R1);
and and6746(N11197,R2,N11201);
and and6747(N11198,N11202,R6);
and and6751(N11206,in0,in2);
and and6752(N11207,N11210,R1);
and and6753(N11208,N11211,N11212);
and and6754(N11209,N11213,R7);
and and6758(N11217,N11221,N11222);
and and6759(N11218,R2,R3);
and and6760(N11219,R4,N11223);
and and6761(N11220,R6,N11224);
and and6765(N11228,in0,N11232);
and and6766(N11229,R1,R2);
and and6767(N11230,N11233,R5);
and and6768(N11231,N11234,N11235);
and and6772(N11239,in1,N11243);
and and6773(N11240,R2,N11244);
and and6774(N11241,R4,R5);
and and6775(N11242,N11245,N11246);
and and6779(N11250,N11254,R0);
and and6780(N11251,R1,N11255);
and and6781(N11252,N11256,R5);
and and6782(N11253,N11257,R7);
and and6786(N11261,in0,N11265);
and and6787(N11262,N11266,R1);
and and6788(N11263,R4,N11267);
and and6789(N11264,N11268,R7);
and and6793(N11272,in0,N11276);
and and6794(N11273,R0,R1);
and and6795(N11274,N11277,R3);
and and6796(N11275,N11278,R7);
and and6800(N11282,in0,N11286);
and and6801(N11283,N11287,R2);
and and6802(N11284,R3,R5);
and and6803(N11285,R6,N11288);
and and6807(N11292,in0,R0);
and and6808(N11293,R1,R2);
and and6809(N11294,N11296,N11297);
and and6810(N11295,R6,N11298);
and and6814(N11302,in0,N11306);
and and6815(N11303,N11307,R2);
and and6816(N11304,R3,R4);
and and6817(N11305,R5,N11308);
and and6821(N11312,in0,in1);
and and6822(N11313,N11316,N11317);
and and6823(N11314,R3,R4);
and and6824(N11315,N11318,R7);
and and6828(N11322,in0,N11326);
and and6829(N11323,N11327,R3);
and and6830(N11324,R4,N11328);
and and6831(N11325,R6,R7);
and and6835(N11332,in0,in1);
and and6836(N11333,N11336,R1);
and and6837(N11334,N11337,R4);
and and6838(N11335,R6,N11338);
and and6842(N11342,in0,in2);
and and6843(N11343,R0,N11346);
and and6844(N11344,R2,N11347);
and and6845(N11345,R5,N11348);
and and6849(N11352,in0,in1);
and and6850(N11353,R0,N11356);
and and6851(N11354,R2,N11357);
and and6852(N11355,R5,N11358);
and and6856(N11362,in0,R0);
and and6857(N11363,R1,R2);
and and6858(N11364,N11366,N11367);
and and6859(N11365,N11368,R7);
and and6863(N11372,N11376,R1);
and and6864(N11373,R2,R3);
and and6865(N11374,N11377,R5);
and and6866(N11375,R6,N11378);
and and6870(N11382,in0,N11386);
and and6871(N11383,N11387,R2);
and and6872(N11384,R3,R5);
and and6873(N11385,R6,N11388);
and and6877(N11392,in0,in2);
and and6878(N11393,N11396,R1);
and and6879(N11394,R2,N11397);
and and6880(N11395,N11398,R6);
and and6884(N11402,in0,in1);
and and6885(N11403,R0,R2);
and and6886(N11404,R4,N11406);
and and6887(N11405,N11407,R7);
and and6891(N11411,N11414,N11415);
and and6892(N11412,N11416,N11417);
and and6893(N11413,N11418,N11419);
and and6897(N11423,N11426,R2);
and and6898(N11424,R3,N11427);
and and6899(N11425,N11428,N11429);
and and3309(N5938,N5945,N5946);
and and3310(N5939,N5947,N5948);
and and3318(N5956,N5963,N5964);
and and3319(N5957,N5965,N5966);
and and3327(N5974,R3,N5982);
and and3328(N5975,N5983,N5984);
and and3336(N5992,N5999,R5);
and and3337(N5993,N6000,N6001);
and and3345(N6009,N6015,N6016);
and and3346(N6010,N6017,N6018);
and and3354(N6026,R3,R5);
and and3355(N6027,N6034,N6035);
and and3363(N6043,R4,N6050);
and and3364(N6044,N6051,N6052);
and and3372(N6060,N6065,N6066);
and and3373(N6061,N6067,N6068);
and and3381(N6076,N6082,N6083);
and and3382(N6077,R6,N6084);
and and3390(N6092,N6098,N6099);
and and3391(N6093,N6100,R7);
and and3399(N6108,R4,N6114);
and and3400(N6109,N6115,N6116);
and and3408(N6124,N6130,N6131);
and and3409(N6125,N6132,R7);
and and3417(N6140,N6145,N6146);
and and3418(N6141,N6147,N6148);
and and3426(N6156,N6162,N6163);
and and3427(N6157,N6164,R7);
and and3435(N6172,N6178,N6179);
and and3436(N6173,N6180,R7);
and and3444(N6188,R4,N6195);
and and3445(N6189,R6,N6196);
and and3453(N6204,R4,N6211);
and and3454(N6205,R6,N6212);
and and3462(N6220,R4,N6227);
and and3463(N6221,N6228,R7);
and and3471(N6236,N6243,R5);
and and3472(N6237,R6,N6244);
and and3480(N6252,R3,N6259);
and and3481(N6253,R5,N6260);
and and3489(N6268,R3,N6274);
and and3490(N6269,N6275,N6276);
and and3498(N6284,N6290,N6291);
and and3499(N6285,N6292,R7);
and and3507(N6300,R4,N6305);
and and3508(N6301,N6306,N6307);
and and3516(N6315,N6319,N6320);
and and3517(N6316,N6321,N6322);
and and3525(N6330,R4,N6335);
and and3526(N6331,N6336,N6337);
and and3534(N6345,R4,R5);
and and3535(N6346,N6351,N6352);
and and3543(N6360,R3,N6366);
and and3544(N6361,R6,N6367);
and and3552(N6375,R4,R5);
and and3553(N6376,N6381,N6382);
and and3561(N6390,R4,N6397);
and and3562(N6391,R6,R7);
and and3570(N6405,N6411,N6412);
and and3571(N6406,R6,R7);
and and3579(N6420,N6425,R5);
and and3580(N6421,N6426,N6427);
and and3588(N6435,N6440,R5);
and and3589(N6436,N6441,N6442);
and and3597(N6450,N6456,N6457);
and and3598(N6451,R6,R7);
and and3606(N6465,N6471,N6472);
and and3607(N6466,R6,R7);
and and3615(N6480,R3,R4);
and and3616(N6481,R5,N6487);
and and3624(N6495,N6501,R5);
and and3625(N6496,N6502,R7);
and and3633(N6510,R4,N6515);
and and3634(N6511,N6516,N6517);
and and3642(N6525,R4,N6532);
and and3643(N6526,R6,R7);
and and3651(N6540,R4,N6545);
and and3652(N6541,N6546,N6547);
and and3660(N6555,N6561,R5);
and and3661(N6556,R6,N6562);
and and3669(N6570,R4,N6577);
and and3670(N6571,R6,R7);
and and3678(N6585,N6590,N6591);
and and3679(N6586,R6,N6592);
and and3687(N6600,R3,N6605);
and and3688(N6601,N6606,N6607);
and and3696(N6615,N6620,N6621);
and and3697(N6616,N6622,R7);
and and3705(N6630,R3,N6636);
and and3706(N6631,N6637,R7);
and and3714(N6645,N6650,R5);
and and3715(N6646,N6651,N6652);
and and3723(N6660,R4,R5);
and and3724(N6661,N6666,N6667);
and and3732(N6675,N6681,R4);
and and3733(N6676,N6682,R7);
and and3741(N6690,N6695,N6696);
and and3742(N6691,R5,N6697);
and and3750(N6705,R3,N6709);
and and3751(N6706,N6710,N6711);
and and3759(N6719,N6724,R5);
and and3760(N6720,N6725,R7);
and and3768(N6733,R4,N6737);
and and3769(N6734,N6738,N6739);
and and3777(N6747,R4,N6752);
and and3778(N6748,N6753,R7);
and and3786(N6761,N6766,R5);
and and3787(N6762,R6,N6767);
and and3795(N6775,R3,N6780);
and and3796(N6776,R6,N6781);
and and3804(N6789,R4,R5);
and and3805(N6790,N6794,N6795);
and and3813(N6803,R3,R4);
and and3814(N6804,N6809,R7);
and and3822(N6817,R3,N6822);
and and3823(N6818,R6,N6823);
and and3831(N6831,R3,N6836);
and and3832(N6832,R6,N6837);
and and3840(N6845,R3,N6850);
and and3841(N6846,N6851,R7);
and and3849(N6859,R3,N6864);
and and3850(N6860,N6865,R7);
and and3858(N6873,N6876,N6877);
and and3859(N6874,N6878,N6879);
and and3867(N6887,N6891,R5);
and and3868(N6888,N6892,N6893);
and and3876(N6901,R4,N6905);
and and3877(N6902,N6906,N6907);
and and3885(N6915,N6919,R4);
and and3886(N6916,N6920,N6921);
and and3894(N6929,R4,N6934);
and and3895(N6930,R6,N6935);
and and3903(N6943,R4,N6948);
and and3904(N6944,R6,N6949);
and and3912(N6957,R4,N6961);
and and3913(N6958,N6962,N6963);
and and3921(N6971,R4,R5);
and and3922(N6972,N6976,N6977);
and and3930(N6985,R3,N6990);
and and3931(N6986,R5,N6991);
and and3939(N6999,R4,N7004);
and and3940(N7000,R6,N7005);
and and3948(N7013,N7018,R4);
and and3949(N7014,N7019,R7);
and and3957(N7027,N7032,N7033);
and and3958(N7028,R6,R7);
and and3966(N7041,N7045,N7046);
and and3967(N7042,N7047,R7);
and and3975(N7055,N7059,N7060);
and and3976(N7056,N7061,R7);
and and3984(N7069,N7073,R5);
and and3985(N7070,N7074,N7075);
and and3993(N7083,N7087,R5);
and and3994(N7084,N7088,N7089);
and and4002(N7097,N7102,R4);
and and4003(N7098,R5,N7103);
and and4011(N7111,R4,N7116);
and and4012(N7112,N7117,R7);
and and4020(N7125,R4,N7128);
and and4021(N7126,N7129,N7130);
and and4029(N7138,R4,N7141);
and and4030(N7139,N7142,N7143);
and and4038(N7151,N7153,N7154);
and and4039(N7152,N7155,N7156);
and and4047(N7164,R4,N7167);
and and4048(N7165,N7168,N7169);
and and4056(N7177,R4,N7180);
and and4057(N7178,N7181,N7182);
and and4065(N7190,R4,N7193);
and and4066(N7191,N7194,N7195);
and and4074(N7203,N7207,R5);
and and4075(N7204,N7208,R7);
and and4083(N7216,N7220,N7221);
and and4084(N7217,R6,R7);
and and4092(N7229,R4,N7234);
and and4093(N7230,R6,R7);
and and4101(N7242,R3,R4);
and and4102(N7243,R5,N7247);
and and4110(N7255,R4,R5);
and and4111(N7256,R6,N7260);
and and4119(N7268,R4,R5);
and and4120(N7269,R6,N7273);
and and4128(N7281,R4,R5);
and and4129(N7282,R6,N7286);
and and4137(N7294,R4,R5);
and and4138(N7295,N7299,R7);
and and4146(N7307,R4,R5);
and and4147(N7308,N7311,N7312);
and and4155(N7320,R3,R5);
and and4156(N7321,R6,R7);
and and4164(N7333,R3,R4);
and and4165(N7334,N7338,R6);
and and4173(N7346,R4,N7351);
and and4174(N7347,R6,R7);
and and4182(N7359,R4,N7364);
and and4183(N7360,R6,R7);
and and4191(N7372,R4,N7377);
and and4192(N7373,R6,R7);
and and4200(N7385,N7390,R5);
and and4201(N7386,R6,R7);
and and4209(N7398,R4,R5);
and and4210(N7399,R6,N7403);
and and4218(N7411,R4,R5);
and and4219(N7412,R6,N7416);
and and4227(N7424,R4,N7429);
and and4228(N7425,R6,R7);
and and4236(N7437,R4,N7442);
and and4237(N7438,R6,R7);
and and4245(N7450,R4,N7455);
and and4246(N7451,R6,R7);
and and4254(N7463,N7467,N7468);
and and4255(N7464,R6,R7);
and and4263(N7476,R3,R4);
and and4264(N7477,R5,R7);
and and4272(N7489,R4,R5);
and and4273(N7490,R6,N7494);
and and4281(N7502,R4,R5);
and and4282(N7503,N7507,R7);
and and4290(N7515,R4,R5);
and and4291(N7516,N7520,R7);
and and4299(N7528,N7531,N7532);
and and4300(N7529,N7533,R7);
and and4308(N7541,R4,N7545);
and and4309(N7542,R6,N7546);
and and4317(N7554,R4,R5);
and and4318(N7555,N7558,N7559);
and and4326(N7567,N7571,N7572);
and and4327(N7568,R6,R7);
and and4335(N7580,N7583,R5);
and and4336(N7581,N7584,N7585);
and and4344(N7593,R4,R5);
and and4345(N7594,N7597,N7598);
and and4353(N7606,R4,N7610);
and and4354(N7607,N7611,R7);
and and4362(N7619,R4,N7621);
and and4363(N7620,N7622,N7623);
and and4371(N7631,R4,R5);
and and4372(N7632,N7635,R7);
and and4380(N7643,R4,R5);
and and4381(N7644,N7647,R7);
and and4389(N7655,N7658,R5);
and and4390(N7656,R6,N7659);
and and4398(N7667,R3,R5);
and and4399(N7668,R6,N7671);
and and4407(N7679,R4,N7683);
and and4408(N7680,R6,R7);
and and4416(N7691,N7694,R5);
and and4417(N7692,R6,N7695);
and and4425(N7703,R3,R4);
and and4426(N7704,R5,N7707);
and and4434(N7715,R4,R5);
and and4435(N7716,R6,R7);
and and4443(N7727,N7731,R5);
and and4444(N7728,R6,R7);
and and4452(N7739,N7743,R5);
and and4453(N7740,R6,R7);
and and4461(N7751,N7755,R5);
and and4462(N7752,R6,R7);
and and4470(N7763,N7767,R5);
and and4471(N7764,R6,R7);
and and4479(N7775,R4,N7779);
and and4480(N7776,R6,R7);
and and4488(N7787,N7790,N7791);
and and4489(N7788,R6,R7);
and and4497(N7799,R3,R4);
and and4498(N7800,R6,N7803);
and and4506(N7811,R4,N7814);
and and4507(N7812,R6,N7815);
and and4515(N7823,R4,R5);
and and4516(N7824,R6,R7);
and and4524(N7835,R4,R5);
and and4525(N7836,R6,R7);
and and4533(N7847,R4,R5);
and and4534(N7848,R6,N7851);
and and4542(N7859,N7863,R4);
and and4543(N7860,R5,R7);
and and4551(N7871,R4,R5);
and and4552(N7872,N7874,N7875);
and and4560(N7883,R4,R5);
and and4561(N7884,N7886,N7887);
and and4569(N7895,R3,R4);
and and4570(N7896,R5,N7899);
and and4578(N7907,R4,R5);
and and4579(N7908,R6,R7);
and and4587(N7918,R4,R5);
and and4588(N7919,R6,R7);
and and4596(N7929,N7931,R5);
and and4597(N7930,N7932,R7);
and and4605(N7940,R3,N7943);
and and4606(N7941,R5,R7);
and and4614(N7951,R4,R5);
and and4615(N7952,R6,N7954);
and and4623(N7962,R3,N7964);
and and4624(N7963,R5,N7965);
and and4632(N7973,N7976,R5);
and and4633(N7974,R6,R7);
and and4641(N7984,R4,R5);
and and4642(N7985,R6,N7987);
and and4650(N7995,R4,R5);
and and4651(N7996,R6,N7998);
and and4659(N8006,N8009,R5);
and and4660(N8007,R6,R7);
and and4668(N8017,R3,R4);
and and4669(N8018,R6,R7);
and and4677(N8028,R4,N8031);
and and4678(N8029,R6,R7);
and and4686(N8039,R3,R4);
and and4687(N8040,R5,R7);
and and4695(N8049,R4,R5);
and and4696(N8050,R6,R7);
and and4704(N8059,R4,R5);
and and4705(N8060,N8061,R7);
and and4713(N8069,R3,R4);
and and4714(N8070,R5,R7);
and and4722(N8079,N8081,R5);
and and4723(N8080,R6,R7);
and and4731(N8089,R4,R5);
and and4732(N8090,R6,R7);
and and4740(N8099,R3,R4);
and and4741(N8100,R5,R7);
and and4749(N8109,R4,N8111);
and and4750(N8110,R6,R7);
and and4758(N8119,R3,R4);
and and4759(N8120,R5,R6);
and and4767(N8128,N8136,R7);
and and4775(N8144,N8151,N8152);
and and4783(N8160,N8166,N8167);
and and4791(N8175,R6,N8182);
and and4799(N8190,N8196,N8197);
and and4807(N8205,N8211,N8212);
and and4815(N8220,R6,N8227);
and and4823(N8235,N8242,R6);
and and4831(N8250,N8256,N8257);
and and4839(N8265,N8271,N8272);
and and4847(N8280,N8286,N8287);
and and4855(N8295,N8302,R7);
and and4863(N8310,N8316,N8317);
and and4871(N8325,N8331,N8332);
and and4879(N8340,N8346,N8347);
and and4887(N8355,N8362,R7);
and and4895(N8370,N8375,N8376);
and and4903(N8384,N8390,R7);
and and4911(N8398,N8404,R7);
and and4919(N8412,N8418,R7);
and and4927(N8426,N8431,N8432);
and and4935(N8440,N8445,N8446);
and and4943(N8454,R6,N8460);
and and4951(N8468,R5,N8474);
and and4959(N8482,N8487,N8488);
and and4967(N8496,N8502,R6);
and and4975(N8510,N8515,N8516);
and and4983(N8524,N8529,N8530);
and and4991(N8538,R6,N8544);
and and4999(N8552,R6,N8558);
and and5007(N8566,R6,N8572);
and and5015(N8580,R6,N8586);
and and5023(N8594,N8599,N8600);
and and5031(N8608,N8613,N8614);
and and5039(N8622,N8627,N8628);
and and5047(N8636,N8641,N8642);
and and5055(N8650,R5,N8656);
and and5063(N8664,R5,N8670);
and and5071(N8678,R5,N8684);
and and5079(N8692,N8697,N8698);
and and5087(N8706,N8711,N8712);
and and5095(N8720,N8726,R7);
and and5103(N8734,N8739,N8740);
and and5111(N8748,N8754,R7);
and and5119(N8762,N8768,R7);
and and5127(N8776,N8782,R7);
and and5135(N8790,R6,N8796);
and and5143(N8804,N8809,N8810);
and and5151(N8818,N8824,R7);
and and5159(N8832,N8837,N8838);
and and5167(N8846,N8851,N8852);
and and5175(N8860,N8865,N8866);
and and5183(N8874,N8879,N8880);
and and5191(N8888,R6,N8894);
and and5199(N8902,N8906,N8907);
and and5207(N8915,R6,R7);
and and5215(N8928,N8932,N8933);
and and5223(N8941,N8946,R7);
and and5231(N8954,N8958,N8959);
and and5239(N8967,N8971,N8972);
and and5247(N8980,N8984,N8985);
and and5255(N8993,N8998,R7);
and and5263(N9006,R6,R7);
and and5271(N9019,N9023,N9024);
and and5279(N9032,R6,N9037);
and and5287(N9045,R6,N9050);
and and5295(N9058,R6,N9063);
and and5303(N9071,R6,N9076);
and and5311(N9084,R6,R7);
and and5319(N9097,N9102,R7);
and and5327(N9110,N9115,R7);
and and5335(N9123,R6,N9128);
and and5343(N9136,R6,N9141);
and and5351(N9149,R6,N9154);
and and5359(N9162,R6,N9167);
and and5367(N9175,R6,N9180);
and and5375(N9188,N9192,N9193);
and and5383(N9201,N9205,N9206);
and and5391(N9214,N9218,N9219);
and and5399(N9227,R5,N9232);
and and5407(N9240,R6,N9245);
and and5415(N9253,N9257,N9258);
and and5423(N9266,N9270,N9271);
and and5431(N9279,N9284,R7);
and and5439(N9292,R6,N9297);
and and5447(N9305,N9310,R7);
and and5455(N9318,N9323,R7);
and and5463(N9331,R6,R7);
and and5471(N9344,N9349,R7);
and and5479(N9357,N9361,N9362);
and and5487(N9370,N9374,N9375);
and and5495(N9383,N9387,N9388);
and and5503(N9396,N9401,R7);
and and5511(N9409,N9414,R7);
and and5519(N9422,N9427,R7);
and and5527(N9435,N9439,N9440);
and and5535(N9448,R5,N9453);
and and5543(N9461,N9466,R6);
and and5551(N9474,R6,N9479);
and and5559(N9487,N9491,N9492);
and and5567(N9500,N9505,R7);
and and5575(N9513,N9517,N9518);
and and5583(N9526,N9530,N9531);
and and5591(N9539,N9544,R7);
and and5599(N9552,N9556,N9557);
and and5607(N9565,N9570,R6);
and and5615(N9578,N9582,N9583);
and and5623(N9591,N9595,N9596);
and and5631(N9604,N9609,R6);
and and5639(N9617,R5,N9622);
and and5647(N9630,N9635,R7);
and and5655(N9643,R6,N9647);
and and5663(N9655,R6,N9659);
and and5671(N9667,R5,N9671);
and and5679(N9679,R6,N9683);
and and5687(N9691,R5,N9695);
and and5695(N9703,R6,N9707);
and and5703(N9715,R6,N9719);
and and5711(N9727,N9731,R7);
and and5719(N9739,N9743,R7);
and and5727(N9751,R6,R7);
and and5735(N9763,R5,N9767);
and and5743(N9775,N9779,R7);
and and5751(N9787,R6,R7);
and and5759(N9799,R6,N9803);
and and5767(N9811,R6,N9815);
and and5775(N9823,N9826,N9827);
and and5783(N9835,R6,R7);
and and5791(N9847,R6,N9851);
and and5799(N9859,N9862,N9863);
and and5807(N9871,N9875,R7);
and and5815(N9883,R6,N9887);
and and5823(N9895,R6,R7);
and and5831(N9907,R6,R7);
and and5839(N9919,N9923,R7);
and and5847(N9931,N9935,R7);
and and5855(N9943,N9947,R7);
and and5863(N9955,N9959,R7);
and and5871(N9967,R6,N9971);
and and5879(N9979,N9983,R7);
and and5887(N9991,N9995,R7);
and and5895(N10003,N10007,R7);
and and5903(N10015,R4,R6);
and and5911(N10027,R5,N10031);
and and5919(N10039,N10043,R7);
and and5927(N10051,N10055,R7);
and and5935(N10063,N10067,R7);
and and5943(N10075,N10079,R7);
and and5951(N10087,N10091,R7);
and and5959(N10099,R6,N10103);
and and5967(N10111,N10115,R6);
and and5975(N10123,R6,R7);
and and5983(N10135,R6,R7);
and and5991(N10147,R6,N10151);
and and5999(N10159,R6,N10163);
and and6007(N10171,N10175,R7);
and and6015(N10183,N10186,N10187);
and and6023(N10195,N10199,R7);
and and6031(N10207,N10209,N10210);
and and6039(N10218,N10221,R7);
and and6047(N10229,N10231,N10232);
and and6055(N10240,R6,R7);
and and6063(N10251,N10254,R7);
and and6071(N10262,N10265,R7);
and and6079(N10273,R5,R6);
and and6087(N10284,N10287,R6);
and and6095(N10295,N10298,R7);
and and6103(N10306,N10308,N10309);
and and6111(N10317,R6,N10320);
and and6119(N10328,N10331,R7);
and and6127(N10339,R4,N10342);
and and6135(N10350,R6,N10353);
and and6143(N10361,N10364,R7);
and and6151(N10372,N10375,R6);
and and6159(N10383,N10386,R7);
and and6167(N10394,N10397,R7);
and and6175(N10405,N10408,R7);
and and6183(N10416,R6,R7);
and and6191(N10427,R6,R7);
and and6199(N10438,R6,R7);
and and6207(N10449,N10452,R7);
and and6215(N10460,N10463,R7);
and and6223(N10471,N10474,R7);
and and6231(N10482,R6,N10485);
and and6239(N10493,R6,N10496);
and and6247(N10504,N10506,N10507);
and and6255(N10515,R6,N10518);
and and6263(N10526,N10528,N10529);
and and6271(N10537,R5,N10540);
and and6279(N10548,N10550,N10551);
and and6287(N10559,R5,N10562);
and and6295(N10570,R6,N10573);
and and6303(N10581,N10584,R7);
and and6311(N10592,R6,N10595);
and and6319(N10603,R6,N10606);
and and6327(N10614,R5,R7);
and and6335(N10625,R6,R7);
and and6343(N10636,N10639,R7);
and and6351(N10647,N10650,R7);
and and6359(N10658,N10661,R7);
and and6367(N10669,R5,N10672);
and and6375(N10680,N10682,R7);
and and6383(N10690,R6,R7);
and and6391(N10700,N10702,R7);
and and6399(N10710,R6,R7);
and and6407(N10720,R6,R7);
and and6415(N10730,N10732,R7);
and and6423(N10740,R6,N10742);
and and6431(N10750,R6,R7);
and and6439(N10760,R6,R7);
and and6447(N10770,R6,N10772);
and and6455(N10780,R6,N10782);
and and6463(N10790,R4,R7);
and and6471(N10800,R6,R7);
and and6479(N10810,R6,R7);
and and6487(N10820,R5,N10822);
and and6495(N10830,R6,R7);
and and6503(N10840,R6,R7);
and and6511(N10850,R6,R7);
and and6519(N10860,R5,R6);
and and6527(N10870,R4,R7);
and and6535(N10880,N10882,R6);
and and6543(N10890,R6,N10892);
and and6551(N10900,N10902,R7);
and and6559(N10910,R6,R7);
and and6567(N10920,N10921,N10922);
and and6575(N10930,R5,R7);
and and6583(N10939,R6,R7);
and and6591(N10948,R6,R7);
and and6599(N10957,R6,R7);
and and6607(N10966,R5,R6);
and and6900(N11882,N11883,N11884);
and and6909(N11900,N11901,N11902);
and and6918(N11918,N11919,N11920);
and and6927(N11935,N11936,N11937);
and and6936(N11952,N11953,N11954);
and and6945(N11969,N11970,N11971);
and and6954(N11986,N11987,N11988);
and and6963(N12002,N12003,N12004);
and and6972(N12018,N12019,N12020);
and and6981(N12034,N12035,N12036);
and and6990(N12050,N12051,N12052);
and and6999(N12066,N12067,N12068);
and and7008(N12082,N12083,N12084);
and and7017(N12098,N12099,N12100);
and and7026(N12114,N12115,N12116);
and and7035(N12130,N12131,N12132);
and and7044(N12146,N12147,N12148);
and and7053(N12162,N12163,N12164);
and and7062(N12178,N12179,N12180);
and and7071(N12194,N12195,N12196);
and and7080(N12209,N12210,N12211);
and and7089(N12224,N12225,N12226);
and and7098(N12239,N12240,N12241);
and and7107(N12254,N12255,N12256);
and and7116(N12269,N12270,N12271);
and and7125(N12284,N12285,N12286);
and and7134(N12299,N12300,N12301);
and and7143(N12314,N12315,N12316);
and and7152(N12329,N12330,N12331);
and and7161(N12344,N12345,N12346);
and and7170(N12359,N12360,N12361);
and and7179(N12374,N12375,N12376);
and and7188(N12389,N12390,N12391);
and and7197(N12404,N12405,N12406);
and and7206(N12419,N12420,N12421);
and and7215(N12434,N12435,N12436);
and and7224(N12449,N12450,N12451);
and and7233(N12464,N12465,N12466);
and and7242(N12479,N12480,N12481);
and and7251(N12494,N12495,N12496);
and and7260(N12509,N12510,N12511);
and and7269(N12524,N12525,N12526);
and and7278(N12539,N12540,N12541);
and and7287(N12554,N12555,N12556);
and and7296(N12569,N12570,N12571);
and and7305(N12584,N12585,N12586);
and and7314(N12599,N12600,N12601);
and and7323(N12614,N12615,N12616);
and and7332(N12629,N12630,N12631);
and and7341(N12644,N12645,N12646);
and and7350(N12659,N12660,N12661);
and and7359(N12674,N12675,N12676);
and and7368(N12689,N12690,N12691);
and and7377(N12704,N12705,N12706);
and and7386(N12719,N12720,N12721);
and and7395(N12734,N12735,N12736);
and and7404(N12749,N12750,N12751);
and and7413(N12763,N12764,N12765);
and and7422(N12777,N12778,N12779);
and and7431(N12791,N12792,N12793);
and and7440(N12805,N12806,N12807);
and and7449(N12819,N12820,N12821);
and and7458(N12833,N12834,N12835);
and and7467(N12847,N12848,N12849);
and and7476(N12861,N12862,N12863);
and and7485(N12875,N12876,N12877);
and and7494(N12889,N12890,N12891);
and and7503(N12903,N12904,N12905);
and and7512(N12917,N12918,N12919);
and and7521(N12931,N12932,N12933);
and and7530(N12945,N12946,N12947);
and and7539(N12959,N12960,N12961);
and and7548(N12973,N12974,N12975);
and and7557(N12987,N12988,N12989);
and and7566(N13001,N13002,N13003);
and and7575(N13015,N13016,N13017);
and and7584(N13029,N13030,N13031);
and and7593(N13043,N13044,N13045);
and and7602(N13057,N13058,N13059);
and and7611(N13071,N13072,N13073);
and and7620(N13085,N13086,N13087);
and and7629(N13099,N13100,N13101);
and and7638(N13113,N13114,N13115);
and and7647(N13127,N13128,N13129);
and and7656(N13141,N13142,N13143);
and and7665(N13155,N13156,N13157);
and and7674(N13169,N13170,N13171);
and and7683(N13183,N13184,N13185);
and and7692(N13197,N13198,N13199);
and and7701(N13211,N13212,N13213);
and and7710(N13225,N13226,N13227);
and and7719(N13239,N13240,N13241);
and and7728(N13253,N13254,N13255);
and and7737(N13267,N13268,N13269);
and and7746(N13281,N13282,N13283);
and and7755(N13295,N13296,N13297);
and and7764(N13309,N13310,N13311);
and and7773(N13323,N13324,N13325);
and and7782(N13336,N13337,N13338);
and and7791(N13349,N13350,N13351);
and and7800(N13362,N13363,N13364);
and and7809(N13375,N13376,N13377);
and and7818(N13388,N13389,N13390);
and and7827(N13401,N13402,N13403);
and and7836(N13414,N13415,N13416);
and and7845(N13427,N13428,N13429);
and and7854(N13440,N13441,N13442);
and and7863(N13453,N13454,N13455);
and and7872(N13466,N13467,N13468);
and and7881(N13479,N13480,N13481);
and and7890(N13492,N13493,N13494);
and and7899(N13505,N13506,N13507);
and and7908(N13518,N13519,N13520);
and and7917(N13531,N13532,N13533);
and and7926(N13544,N13545,N13546);
and and7935(N13557,N13558,N13559);
and and7944(N13570,N13571,N13572);
and and7953(N13583,N13584,N13585);
and and7962(N13596,N13597,N13598);
and and7971(N13609,N13610,N13611);
and and7980(N13622,N13623,N13624);
and and7989(N13635,N13636,N13637);
and and7998(N13648,N13649,N13650);
and and8007(N13661,N13662,N13663);
and and8016(N13674,N13675,N13676);
and and8025(N13687,N13688,N13689);
and and8034(N13700,N13701,N13702);
and and8043(N13713,N13714,N13715);
and and8052(N13726,N13727,N13728);
and and8061(N13739,N13740,N13741);
and and8070(N13752,N13753,N13754);
and and8079(N13765,N13766,N13767);
and and8088(N13778,N13779,N13780);
and and8097(N13791,N13792,N13793);
and and8106(N13804,N13805,N13806);
and and8115(N13817,N13818,N13819);
and and8124(N13830,N13831,N13832);
and and8133(N13843,N13844,N13845);
and and8142(N13856,N13857,N13858);
and and8151(N13869,N13870,N13871);
and and8160(N13882,N13883,N13884);
and and8169(N13895,N13896,N13897);
and and8178(N13908,N13909,N13910);
and and8187(N13921,N13922,N13923);
and and8196(N13933,N13934,N13935);
and and8205(N13945,N13946,N13947);
and and8214(N13957,N13958,N13959);
and and8223(N13969,N13970,N13971);
and and8232(N13981,N13982,N13983);
and and8241(N13993,N13994,N13995);
and and8250(N14005,N14006,N14007);
and and8259(N14017,N14018,N14019);
and and8268(N14029,N14030,N14031);
and and8277(N14041,N14042,N14043);
and and8286(N14053,N14054,N14055);
and and8295(N14065,N14066,N14067);
and and8304(N14077,N14078,N14079);
and and8313(N14089,N14090,N14091);
and and8322(N14101,N14102,N14103);
and and8331(N14113,N14114,N14115);
and and8340(N14125,N14126,N14127);
and and8349(N14137,N14138,N14139);
and and8358(N14149,N14150,N14151);
and and8367(N14161,N14162,N14163);
and and8376(N14173,N14174,N14175);
and and8385(N14185,N14186,N14187);
and and8394(N14197,N14198,N14199);
and and8403(N14209,N14210,N14211);
and and8412(N14221,N14222,N14223);
and and8421(N14233,N14234,N14235);
and and8430(N14245,N14246,N14247);
and and8439(N14257,N14258,N14259);
and and8448(N14268,N14269,N14270);
and and8457(N14279,N14280,N14281);
and and8466(N14290,N14291,N14292);
and and8475(N14301,N14302,N14303);
and and8484(N14312,N14313,N14314);
and and8493(N14323,N14324,N14325);
and and8502(N14334,N14335,N14336);
and and8511(N14345,N14346,N14347);
and and8520(N14356,N14357,N14358);
and and8529(N14367,N14368,N14369);
and and8538(N14378,N14379,N14380);
and and8547(N14389,N14390,N14391);
and and8556(N14400,N14401,N14402);
and and8565(N14411,N14412,N14413);
and and8574(N14422,N14423,N14424);
and and8583(N14433,N14434,N14435);
and and8592(N14443,N14444,N14445);
and and8601(N14453,N14454,N14455);
and and8610(N14463,N14464,N14465);
and and8619(N14473,N14474,N14475);
and and8628(N14483,N14484,N14485);
and and8637(N14493,N14494,N14495);
and and8646(N14502,N14503,N14504);
and and8654(N14518,N14519,N14520);
and and8662(N14534,N14535,N14536);
and and8670(N14550,N14551,N14552);
and and8678(N14565,N14566,N14567);
and and8686(N14580,N14581,N14582);
and and8694(N14595,N14596,N14597);
and and8702(N14610,N14611,N14612);
and and8710(N14625,N14626,N14627);
and and8718(N14640,N14641,N14642);
and and8726(N14655,N14656,N14657);
and and8734(N14670,N14671,N14672);
and and8742(N14685,N14686,N14687);
and and8750(N14700,N14701,N14702);
and and8758(N14714,N14715,N14716);
and and8766(N14728,N14729,N14730);
and and8774(N14742,N14743,N14744);
and and8782(N14756,N14757,N14758);
and and8790(N14770,N14771,N14772);
and and8798(N14784,N14785,N14786);
and and8806(N14798,N14799,N14800);
and and8814(N14812,N14813,N14814);
and and8822(N14826,N14827,N14828);
and and8830(N14840,N14841,N14842);
and and8838(N14854,N14855,N14856);
and and8846(N14868,N14869,N14870);
and and8854(N14882,N14883,N14884);
and and8862(N14896,N14897,N14898);
and and8870(N14910,N14911,N14912);
and and8878(N14924,N14925,N14926);
and and8886(N14938,N14939,N14940);
and and8894(N14952,N14953,N14954);
and and8902(N14966,N14967,N14968);
and and8910(N14980,N14981,N14982);
and and8918(N14994,N14995,N14996);
and and8926(N15008,N15009,N15010);
and and8934(N15022,N15023,N15024);
and and8942(N15036,N15037,N15038);
and and8950(N15050,N15051,N15052);
and and8958(N15064,N15065,N15066);
and and8966(N15078,N15079,N15080);
and and8974(N15092,N15093,N15094);
and and8982(N15106,N15107,N15108);
and and8990(N15120,N15121,N15122);
and and8998(N15134,N15135,N15136);
and and9006(N15148,N15149,N15150);
and and9014(N15162,N15163,N15164);
and and9022(N15176,N15177,N15178);
and and9030(N15190,N15191,N15192);
and and9038(N15203,N15204,N15205);
and and9046(N15216,N15217,N15218);
and and9054(N15229,N15230,N15231);
and and9062(N15242,N15243,N15244);
and and9070(N15255,N15256,N15257);
and and9078(N15268,N15269,N15270);
and and9086(N15281,N15282,N15283);
and and9094(N15294,N15295,N15296);
and and9102(N15307,N15308,N15309);
and and9110(N15320,N15321,N15322);
and and9118(N15333,N15334,N15335);
and and9126(N15346,N15347,N15348);
and and9134(N15359,N15360,N15361);
and and9142(N15372,N15373,N15374);
and and9150(N15385,N15386,N15387);
and and9158(N15398,N15399,N15400);
and and9166(N15411,N15412,N15413);
and and9174(N15424,N15425,N15426);
and and9182(N15437,N15438,N15439);
and and9190(N15450,N15451,N15452);
and and9198(N15463,N15464,N15465);
and and9206(N15476,N15477,N15478);
and and9214(N15489,N15490,N15491);
and and9222(N15502,N15503,N15504);
and and9230(N15515,N15516,N15517);
and and9238(N15528,N15529,N15530);
and and9246(N15541,N15542,N15543);
and and9254(N15554,N15555,N15556);
and and9262(N15567,N15568,N15569);
and and9270(N15580,N15581,N15582);
and and9278(N15593,N15594,N15595);
and and9286(N15606,N15607,N15608);
and and9294(N15619,N15620,N15621);
and and9302(N15632,N15633,N15634);
and and9310(N15645,N15646,N15647);
and and9318(N15658,N15659,N15660);
and and9326(N15671,N15672,N15673);
and and9334(N15684,N15685,N15686);
and and9342(N15697,N15698,N15699);
and and9350(N15710,N15711,N15712);
and and9358(N15723,N15724,N15725);
and and9366(N15736,N15737,N15738);
and and9374(N15749,N15750,N15751);
and and9382(N15762,N15763,N15764);
and and9390(N15775,N15776,N15777);
and and9398(N15788,N15789,N15790);
and and9406(N15801,N15802,N15803);
and and9414(N15814,N15815,N15816);
and and9422(N15826,N15827,N15828);
and and9430(N15838,N15839,N15840);
and and9438(N15850,N15851,N15852);
and and9446(N15862,N15863,N15864);
and and9454(N15874,N15875,N15876);
and and9462(N15886,N15887,N15888);
and and9470(N15898,N15899,N15900);
and and9478(N15910,N15911,N15912);
and and9486(N15922,N15923,N15924);
and and9494(N15934,N15935,N15936);
and and9502(N15946,N15947,N15948);
and and9510(N15958,N15959,N15960);
and and9518(N15970,N15971,N15972);
and and9526(N15982,N15983,N15984);
and and9534(N15994,N15995,N15996);
and and9542(N16006,N16007,N16008);
and and9550(N16018,N16019,N16020);
and and9558(N16030,N16031,N16032);
and and9566(N16042,N16043,N16044);
and and9574(N16054,N16055,N16056);
and and9582(N16066,N16067,N16068);
and and9590(N16078,N16079,N16080);
and and9598(N16090,N16091,N16092);
and and9606(N16102,N16103,N16104);
and and9614(N16114,N16115,N16116);
and and9622(N16126,N16127,N16128);
and and9630(N16138,N16139,N16140);
and and9638(N16150,N16151,N16152);
and and9646(N16162,N16163,N16164);
and and9654(N16174,N16175,N16176);
and and9662(N16186,N16187,N16188);
and and9670(N16198,N16199,N16200);
and and9678(N16210,N16211,N16212);
and and9686(N16222,N16223,N16224);
and and9694(N16234,N16235,N16236);
and and9702(N16246,N16247,N16248);
and and9710(N16258,N16259,N16260);
and and9718(N16270,N16271,N16272);
and and9726(N16282,N16283,N16284);
and and9734(N16294,N16295,N16296);
and and9742(N16306,N16307,N16308);
and and9750(N16318,N16319,N16320);
and and9758(N16330,N16331,N16332);
and and9766(N16342,N16343,N16344);
and and9774(N16354,N16355,N16356);
and and9782(N16366,N16367,N16368);
and and9790(N16378,N16379,N16380);
and and9798(N16390,N16391,N16392);
and and9806(N16402,N16403,N16404);
and and9814(N16414,N16415,N16416);
and and9822(N16426,N16427,N16428);
and and9830(N16438,N16439,N16440);
and and9838(N16450,N16451,N16452);
and and9846(N16461,N16462,N16463);
and and9854(N16472,N16473,N16474);
and and9862(N16483,N16484,N16485);
and and9870(N16494,N16495,N16496);
and and9878(N16505,N16506,N16507);
and and9886(N16516,N16517,N16518);
and and9894(N16527,N16528,N16529);
and and9902(N16538,N16539,N16540);
and and9910(N16549,N16550,N16551);
and and9918(N16560,N16561,N16562);
and and9926(N16571,N16572,N16573);
and and9934(N16582,N16583,N16584);
and and9942(N16593,N16594,N16595);
and and9950(N16604,N16605,N16606);
and and9958(N16615,N16616,N16617);
and and9966(N16626,N16627,N16628);
and and9974(N16637,N16638,N16639);
and and9982(N16648,N16649,N16650);
and and9990(N16659,N16660,N16661);
and and9998(N16670,N16671,N16672);
and and10006(N16681,N16682,N16683);
and and10014(N16692,N16693,N16694);
and and10022(N16703,N16704,N16705);
and and10030(N16714,N16715,N16716);
and and10038(N16725,N16726,N16727);
and and10046(N16736,N16737,N16738);
and and10054(N16747,N16748,N16749);
and and10062(N16758,N16759,N16760);
and and10070(N16769,N16770,N16771);
and and10078(N16780,N16781,N16782);
and and10086(N16791,N16792,N16793);
and and10094(N16802,N16803,N16804);
and and10102(N16813,N16814,N16815);
and and10110(N16824,N16825,N16826);
and and10118(N16835,N16836,N16837);
and and10126(N16846,N16847,N16848);
and and10134(N16857,N16858,N16859);
and and10142(N16868,N16869,N16870);
and and10150(N16879,N16880,N16881);
and and10158(N16890,N16891,N16892);
and and10166(N16900,N16901,N16902);
and and10174(N16910,N16911,N16912);
and and10182(N16920,N16921,N16922);
and and10190(N16930,N16931,N16932);
and and10198(N16940,N16941,N16942);
and and10206(N16950,N16951,N16952);
and and10214(N16960,N16961,N16962);
and and10222(N16970,N16971,N16972);
and and10230(N16980,N16981,N16982);
and and10238(N16990,N16991,N16992);
and and10246(N17000,N17001,N17002);
and and10254(N17010,N17011,N17012);
and and10262(N17020,N17021,N17022);
and and10270(N17030,N17031,N17032);
and and10278(N17040,N17041,N17042);
and and10286(N17050,N17051,N17052);
and and10294(N17060,N17061,N17062);
and and10302(N17069,N17070,N17071);
and and10310(N17078,N17079,N17080);
and and10318(N17087,N17088,N17089);
and and10326(N17096,N17097,N17098);
and and10334(N17105,N17106,N17107);
and and10342(N17114,N17115,N17116);
and and10350(N17123,N17124,N17125);
and and10358(N17132,N17133,N17134);
and and10366(N17141,N17142,N17143);
and and10374(N17150,N17151,N17152);
and and10382(N17158,N17159,N17160);
and and10389(N17172,N17173,N17174);
and and10396(N17186,N17187,N17188);
and and10403(N17200,N17201,N17202);
and and10410(N17214,N17215,N17216);
and and10417(N17227,N17228,N17229);
and and10424(N17240,N17241,N17242);
and and10431(N17253,N17254,N17255);
and and10438(N17266,N17267,N17268);
and and10445(N17279,N17280,N17281);
and and10452(N17291,N17292,N17293);
and and10459(N17303,N17304,N17305);
and and10466(N17315,N17316,N17317);
and and10473(N17327,N17328,N17329);
and and10480(N17339,N17340,N17341);
and and10487(N17351,N17352,N17353);
and and10494(N17363,N17364,N17365);
and and10501(N17375,N17376,N17377);
and and10508(N17387,N17388,N17389);
and and10515(N17398,N17399,N17400);
and and10522(N17409,N17410,N17411);
and and10529(N17420,N17421,N17422);
and and10536(N17431,N17432,N17433);
and and10543(N17442,N17443,N17444);
and and10550(N17453,N17454,N17455);
and and10557(N17464,N17465,N17466);
and and10564(N17475,N17476,N17477);
and and10571(N17486,N17487,N17488);
and and10578(N17497,N17498,N17499);
and and10585(N17508,N17509,N17510);
and and10592(N17519,N17520,N17521);
and and10599(N17530,N17531,N17532);
and and10606(N17541,N17542,N17543);
and and10613(N17552,N17553,N17554);
and and10620(N17563,N17564,N17565);
and and10627(N17574,N17575,N17576);
and and10634(N17584,N17585,N17586);
and and10641(N17594,N17595,N17596);
and and10648(N17604,N17605,N17606);
and and10655(N17614,N17615,N17616);
and and10662(N17624,N17625,N17626);
and and10669(N17634,N17635,N17636);
and and6901(N11883,N11885,N11886);
and and6902(N11884,N11887,N11888);
and and6910(N11901,N11903,N11904);
and and6911(N11902,N11905,N11906);
and and6919(N11919,N11921,N11922);
and and6920(N11920,N11923,N11924);
and and6928(N11936,N11938,N11939);
and and6929(N11937,N11940,N11941);
and and6937(N11953,N11955,N11956);
and and6938(N11954,N11957,N11958);
and and6946(N11970,N11972,N11973);
and and6947(N11971,N11974,N11975);
and and6955(N11987,N11989,N11990);
and and6956(N11988,N11991,N11992);
and and6964(N12003,N12005,N12006);
and and6965(N12004,N12007,N12008);
and and6973(N12019,N12021,N12022);
and and6974(N12020,N12023,N12024);
and and6982(N12035,N12037,N12038);
and and6983(N12036,N12039,N12040);
and and6991(N12051,N12053,N12054);
and and6992(N12052,N12055,N12056);
and and7000(N12067,N12069,N12070);
and and7001(N12068,N12071,N12072);
and and7009(N12083,N12085,N12086);
and and7010(N12084,N12087,N12088);
and and7018(N12099,N12101,N12102);
and and7019(N12100,N12103,N12104);
and and7027(N12115,N12117,N12118);
and and7028(N12116,N12119,N12120);
and and7036(N12131,N12133,N12134);
and and7037(N12132,N12135,N12136);
and and7045(N12147,N12149,N12150);
and and7046(N12148,N12151,N12152);
and and7054(N12163,N12165,N12166);
and and7055(N12164,N12167,N12168);
and and7063(N12179,N12181,N12182);
and and7064(N12180,N12183,N12184);
and and7072(N12195,N12197,N12198);
and and7073(N12196,N12199,N12200);
and and7081(N12210,N12212,N12213);
and and7082(N12211,N12214,N12215);
and and7090(N12225,N12227,N12228);
and and7091(N12226,N12229,N12230);
and and7099(N12240,N12242,N12243);
and and7100(N12241,N12244,N12245);
and and7108(N12255,N12257,N12258);
and and7109(N12256,N12259,N12260);
and and7117(N12270,N12272,N12273);
and and7118(N12271,N12274,N12275);
and and7126(N12285,N12287,N12288);
and and7127(N12286,N12289,N12290);
and and7135(N12300,N12302,N12303);
and and7136(N12301,N12304,N12305);
and and7144(N12315,N12317,N12318);
and and7145(N12316,N12319,N12320);
and and7153(N12330,N12332,N12333);
and and7154(N12331,N12334,N12335);
and and7162(N12345,N12347,N12348);
and and7163(N12346,N12349,N12350);
and and7171(N12360,N12362,N12363);
and and7172(N12361,N12364,N12365);
and and7180(N12375,N12377,N12378);
and and7181(N12376,N12379,N12380);
and and7189(N12390,N12392,N12393);
and and7190(N12391,N12394,N12395);
and and7198(N12405,N12407,N12408);
and and7199(N12406,N12409,N12410);
and and7207(N12420,N12422,N12423);
and and7208(N12421,N12424,N12425);
and and7216(N12435,N12437,N12438);
and and7217(N12436,N12439,N12440);
and and7225(N12450,N12452,N12453);
and and7226(N12451,N12454,N12455);
and and7234(N12465,N12467,N12468);
and and7235(N12466,N12469,N12470);
and and7243(N12480,N12482,N12483);
and and7244(N12481,N12484,N12485);
and and7252(N12495,N12497,N12498);
and and7253(N12496,N12499,N12500);
and and7261(N12510,N12512,N12513);
and and7262(N12511,N12514,N12515);
and and7270(N12525,N12527,N12528);
and and7271(N12526,N12529,N12530);
and and7279(N12540,N12542,N12543);
and and7280(N12541,N12544,N12545);
and and7288(N12555,N12557,N12558);
and and7289(N12556,N12559,N12560);
and and7297(N12570,N12572,N12573);
and and7298(N12571,N12574,N12575);
and and7306(N12585,N12587,N12588);
and and7307(N12586,N12589,N12590);
and and7315(N12600,N12602,N12603);
and and7316(N12601,N12604,N12605);
and and7324(N12615,N12617,N12618);
and and7325(N12616,N12619,N12620);
and and7333(N12630,N12632,N12633);
and and7334(N12631,N12634,N12635);
and and7342(N12645,N12647,N12648);
and and7343(N12646,N12649,N12650);
and and7351(N12660,N12662,N12663);
and and7352(N12661,N12664,N12665);
and and7360(N12675,N12677,N12678);
and and7361(N12676,N12679,N12680);
and and7369(N12690,N12692,N12693);
and and7370(N12691,N12694,N12695);
and and7378(N12705,N12707,N12708);
and and7379(N12706,N12709,N12710);
and and7387(N12720,N12722,N12723);
and and7388(N12721,N12724,N12725);
and and7396(N12735,N12737,N12738);
and and7397(N12736,N12739,N12740);
and and7405(N12750,N12752,N12753);
and and7406(N12751,N12754,N12755);
and and7414(N12764,N12766,N12767);
and and7415(N12765,N12768,N12769);
and and7423(N12778,N12780,N12781);
and and7424(N12779,N12782,N12783);
and and7432(N12792,N12794,N12795);
and and7433(N12793,N12796,N12797);
and and7441(N12806,N12808,N12809);
and and7442(N12807,N12810,N12811);
and and7450(N12820,N12822,N12823);
and and7451(N12821,N12824,N12825);
and and7459(N12834,N12836,N12837);
and and7460(N12835,N12838,N12839);
and and7468(N12848,N12850,N12851);
and and7469(N12849,N12852,N12853);
and and7477(N12862,N12864,N12865);
and and7478(N12863,N12866,N12867);
and and7486(N12876,N12878,N12879);
and and7487(N12877,N12880,N12881);
and and7495(N12890,N12892,N12893);
and and7496(N12891,N12894,N12895);
and and7504(N12904,N12906,N12907);
and and7505(N12905,N12908,N12909);
and and7513(N12918,N12920,N12921);
and and7514(N12919,N12922,N12923);
and and7522(N12932,N12934,N12935);
and and7523(N12933,N12936,N12937);
and and7531(N12946,N12948,N12949);
and and7532(N12947,N12950,N12951);
and and7540(N12960,N12962,N12963);
and and7541(N12961,N12964,N12965);
and and7549(N12974,N12976,N12977);
and and7550(N12975,N12978,N12979);
and and7558(N12988,N12990,N12991);
and and7559(N12989,N12992,N12993);
and and7567(N13002,N13004,N13005);
and and7568(N13003,N13006,N13007);
and and7576(N13016,N13018,N13019);
and and7577(N13017,N13020,N13021);
and and7585(N13030,N13032,N13033);
and and7586(N13031,N13034,N13035);
and and7594(N13044,N13046,N13047);
and and7595(N13045,N13048,N13049);
and and7603(N13058,N13060,N13061);
and and7604(N13059,N13062,N13063);
and and7612(N13072,N13074,N13075);
and and7613(N13073,N13076,N13077);
and and7621(N13086,N13088,N13089);
and and7622(N13087,N13090,N13091);
and and7630(N13100,N13102,N13103);
and and7631(N13101,N13104,N13105);
and and7639(N13114,N13116,N13117);
and and7640(N13115,N13118,N13119);
and and7648(N13128,N13130,N13131);
and and7649(N13129,N13132,N13133);
and and7657(N13142,N13144,N13145);
and and7658(N13143,N13146,N13147);
and and7666(N13156,N13158,N13159);
and and7667(N13157,N13160,N13161);
and and7675(N13170,N13172,N13173);
and and7676(N13171,N13174,N13175);
and and7684(N13184,N13186,N13187);
and and7685(N13185,N13188,N13189);
and and7693(N13198,N13200,N13201);
and and7694(N13199,N13202,N13203);
and and7702(N13212,N13214,N13215);
and and7703(N13213,N13216,N13217);
and and7711(N13226,N13228,N13229);
and and7712(N13227,N13230,N13231);
and and7720(N13240,N13242,N13243);
and and7721(N13241,N13244,N13245);
and and7729(N13254,N13256,N13257);
and and7730(N13255,N13258,N13259);
and and7738(N13268,N13270,N13271);
and and7739(N13269,N13272,N13273);
and and7747(N13282,N13284,N13285);
and and7748(N13283,N13286,N13287);
and and7756(N13296,N13298,N13299);
and and7757(N13297,N13300,N13301);
and and7765(N13310,N13312,N13313);
and and7766(N13311,N13314,N13315);
and and7774(N13324,N13326,N13327);
and and7775(N13325,N13328,N13329);
and and7783(N13337,N13339,N13340);
and and7784(N13338,N13341,N13342);
and and7792(N13350,N13352,N13353);
and and7793(N13351,N13354,N13355);
and and7801(N13363,N13365,N13366);
and and7802(N13364,N13367,N13368);
and and7810(N13376,N13378,N13379);
and and7811(N13377,N13380,N13381);
and and7819(N13389,N13391,N13392);
and and7820(N13390,N13393,N13394);
and and7828(N13402,N13404,N13405);
and and7829(N13403,N13406,N13407);
and and7837(N13415,N13417,N13418);
and and7838(N13416,N13419,N13420);
and and7846(N13428,N13430,N13431);
and and7847(N13429,N13432,N13433);
and and7855(N13441,N13443,N13444);
and and7856(N13442,N13445,N13446);
and and7864(N13454,N13456,N13457);
and and7865(N13455,N13458,N13459);
and and7873(N13467,N13469,N13470);
and and7874(N13468,N13471,N13472);
and and7882(N13480,N13482,N13483);
and and7883(N13481,N13484,N13485);
and and7891(N13493,N13495,N13496);
and and7892(N13494,N13497,N13498);
and and7900(N13506,N13508,N13509);
and and7901(N13507,N13510,N13511);
and and7909(N13519,N13521,N13522);
and and7910(N13520,N13523,N13524);
and and7918(N13532,N13534,N13535);
and and7919(N13533,N13536,N13537);
and and7927(N13545,N13547,N13548);
and and7928(N13546,N13549,N13550);
and and7936(N13558,N13560,N13561);
and and7937(N13559,N13562,N13563);
and and7945(N13571,N13573,N13574);
and and7946(N13572,N13575,N13576);
and and7954(N13584,N13586,N13587);
and and7955(N13585,N13588,N13589);
and and7963(N13597,N13599,N13600);
and and7964(N13598,N13601,N13602);
and and7972(N13610,N13612,N13613);
and and7973(N13611,N13614,N13615);
and and7981(N13623,N13625,N13626);
and and7982(N13624,N13627,N13628);
and and7990(N13636,N13638,N13639);
and and7991(N13637,N13640,N13641);
and and7999(N13649,N13651,N13652);
and and8000(N13650,N13653,N13654);
and and8008(N13662,N13664,N13665);
and and8009(N13663,N13666,N13667);
and and8017(N13675,N13677,N13678);
and and8018(N13676,N13679,N13680);
and and8026(N13688,N13690,N13691);
and and8027(N13689,N13692,N13693);
and and8035(N13701,N13703,N13704);
and and8036(N13702,N13705,N13706);
and and8044(N13714,N13716,N13717);
and and8045(N13715,N13718,N13719);
and and8053(N13727,N13729,N13730);
and and8054(N13728,N13731,N13732);
and and8062(N13740,N13742,N13743);
and and8063(N13741,N13744,N13745);
and and8071(N13753,N13755,N13756);
and and8072(N13754,N13757,N13758);
and and8080(N13766,N13768,N13769);
and and8081(N13767,N13770,N13771);
and and8089(N13779,N13781,N13782);
and and8090(N13780,N13783,N13784);
and and8098(N13792,N13794,N13795);
and and8099(N13793,N13796,N13797);
and and8107(N13805,N13807,N13808);
and and8108(N13806,N13809,N13810);
and and8116(N13818,N13820,N13821);
and and8117(N13819,N13822,N13823);
and and8125(N13831,N13833,N13834);
and and8126(N13832,N13835,N13836);
and and8134(N13844,N13846,N13847);
and and8135(N13845,N13848,N13849);
and and8143(N13857,N13859,N13860);
and and8144(N13858,N13861,N13862);
and and8152(N13870,N13872,N13873);
and and8153(N13871,N13874,N13875);
and and8161(N13883,N13885,N13886);
and and8162(N13884,N13887,N13888);
and and8170(N13896,N13898,N13899);
and and8171(N13897,N13900,N13901);
and and8179(N13909,N13911,N13912);
and and8180(N13910,N13913,N13914);
and and8188(N13922,N13924,N13925);
and and8189(N13923,N13926,N13927);
and and8197(N13934,N13936,N13937);
and and8198(N13935,N13938,N13939);
and and8206(N13946,N13948,N13949);
and and8207(N13947,N13950,N13951);
and and8215(N13958,N13960,N13961);
and and8216(N13959,N13962,N13963);
and and8224(N13970,N13972,N13973);
and and8225(N13971,N13974,N13975);
and and8233(N13982,N13984,N13985);
and and8234(N13983,N13986,N13987);
and and8242(N13994,N13996,N13997);
and and8243(N13995,N13998,N13999);
and and8251(N14006,N14008,N14009);
and and8252(N14007,N14010,N14011);
and and8260(N14018,N14020,N14021);
and and8261(N14019,N14022,N14023);
and and8269(N14030,N14032,N14033);
and and8270(N14031,N14034,N14035);
and and8278(N14042,N14044,N14045);
and and8279(N14043,N14046,N14047);
and and8287(N14054,N14056,N14057);
and and8288(N14055,N14058,N14059);
and and8296(N14066,N14068,N14069);
and and8297(N14067,N14070,N14071);
and and8305(N14078,N14080,N14081);
and and8306(N14079,N14082,N14083);
and and8314(N14090,N14092,N14093);
and and8315(N14091,N14094,N14095);
and and8323(N14102,N14104,N14105);
and and8324(N14103,N14106,N14107);
and and8332(N14114,N14116,N14117);
and and8333(N14115,N14118,N14119);
and and8341(N14126,N14128,N14129);
and and8342(N14127,N14130,N14131);
and and8350(N14138,N14140,N14141);
and and8351(N14139,N14142,N14143);
and and8359(N14150,N14152,N14153);
and and8360(N14151,N14154,N14155);
and and8368(N14162,N14164,N14165);
and and8369(N14163,N14166,N14167);
and and8377(N14174,N14176,N14177);
and and8378(N14175,N14178,N14179);
and and8386(N14186,N14188,N14189);
and and8387(N14187,N14190,N14191);
and and8395(N14198,N14200,N14201);
and and8396(N14199,N14202,N14203);
and and8404(N14210,N14212,N14213);
and and8405(N14211,N14214,N14215);
and and8413(N14222,N14224,N14225);
and and8414(N14223,N14226,N14227);
and and8422(N14234,N14236,N14237);
and and8423(N14235,N14238,N14239);
and and8431(N14246,N14248,N14249);
and and8432(N14247,N14250,N14251);
and and8440(N14258,N14260,N14261);
and and8441(N14259,N14262,N14263);
and and8449(N14269,N14271,N14272);
and and8450(N14270,N14273,N14274);
and and8458(N14280,N14282,N14283);
and and8459(N14281,N14284,N14285);
and and8467(N14291,N14293,N14294);
and and8468(N14292,N14295,N14296);
and and8476(N14302,N14304,N14305);
and and8477(N14303,N14306,N14307);
and and8485(N14313,N14315,N14316);
and and8486(N14314,N14317,N14318);
and and8494(N14324,N14326,N14327);
and and8495(N14325,N14328,N14329);
and and8503(N14335,N14337,N14338);
and and8504(N14336,N14339,N14340);
and and8512(N14346,N14348,N14349);
and and8513(N14347,N14350,N14351);
and and8521(N14357,N14359,N14360);
and and8522(N14358,N14361,N14362);
and and8530(N14368,N14370,N14371);
and and8531(N14369,N14372,N14373);
and and8539(N14379,N14381,N14382);
and and8540(N14380,N14383,N14384);
and and8548(N14390,N14392,N14393);
and and8549(N14391,N14394,N14395);
and and8557(N14401,N14403,N14404);
and and8558(N14402,N14405,N14406);
and and8566(N14412,N14414,N14415);
and and8567(N14413,N14416,N14417);
and and8575(N14423,N14425,N14426);
and and8576(N14424,N14427,N14428);
and and8584(N14434,N14436,N14437);
and and8585(N14435,N14438,N14439);
and and8593(N14444,N14446,N14447);
and and8594(N14445,N14448,N14449);
and and8602(N14454,N14456,N14457);
and and8603(N14455,N14458,N14459);
and and8611(N14464,N14466,N14467);
and and8612(N14465,N14468,N14469);
and and8620(N14474,N14476,N14477);
and and8621(N14475,N14478,N14479);
and and8629(N14484,N14486,N14487);
and and8630(N14485,N14488,N14489);
and and8638(N14494,N14496,N14497);
and and8639(N14495,N14498,N14499);
and and8647(N14503,N14505,N14506);
and and8648(N14504,N14507,N14508);
and and8655(N14519,N14521,N14522);
and and8656(N14520,N14523,N14524);
and and8663(N14535,N14537,N14538);
and and8664(N14536,N14539,N14540);
and and8671(N14551,N14553,N14554);
and and8672(N14552,N14555,N14556);
and and8679(N14566,N14568,N14569);
and and8680(N14567,N14570,N14571);
and and8687(N14581,N14583,N14584);
and and8688(N14582,N14585,N14586);
and and8695(N14596,N14598,N14599);
and and8696(N14597,N14600,N14601);
and and8703(N14611,N14613,N14614);
and and8704(N14612,N14615,N14616);
and and8711(N14626,N14628,N14629);
and and8712(N14627,N14630,N14631);
and and8719(N14641,N14643,N14644);
and and8720(N14642,N14645,N14646);
and and8727(N14656,N14658,N14659);
and and8728(N14657,N14660,N14661);
and and8735(N14671,N14673,N14674);
and and8736(N14672,N14675,N14676);
and and8743(N14686,N14688,N14689);
and and8744(N14687,N14690,N14691);
and and8751(N14701,N14703,N14704);
and and8752(N14702,N14705,N14706);
and and8759(N14715,N14717,N14718);
and and8760(N14716,N14719,N14720);
and and8767(N14729,N14731,N14732);
and and8768(N14730,N14733,N14734);
and and8775(N14743,N14745,N14746);
and and8776(N14744,N14747,N14748);
and and8783(N14757,N14759,N14760);
and and8784(N14758,N14761,N14762);
and and8791(N14771,N14773,N14774);
and and8792(N14772,N14775,N14776);
and and8799(N14785,N14787,N14788);
and and8800(N14786,N14789,N14790);
and and8807(N14799,N14801,N14802);
and and8808(N14800,N14803,N14804);
and and8815(N14813,N14815,N14816);
and and8816(N14814,N14817,N14818);
and and8823(N14827,N14829,N14830);
and and8824(N14828,N14831,N14832);
and and8831(N14841,N14843,N14844);
and and8832(N14842,N14845,N14846);
and and8839(N14855,N14857,N14858);
and and8840(N14856,N14859,N14860);
and and8847(N14869,N14871,N14872);
and and8848(N14870,N14873,N14874);
and and8855(N14883,N14885,N14886);
and and8856(N14884,N14887,N14888);
and and8863(N14897,N14899,N14900);
and and8864(N14898,N14901,N14902);
and and8871(N14911,N14913,N14914);
and and8872(N14912,N14915,N14916);
and and8879(N14925,N14927,N14928);
and and8880(N14926,N14929,N14930);
and and8887(N14939,N14941,N14942);
and and8888(N14940,N14943,N14944);
and and8895(N14953,N14955,N14956);
and and8896(N14954,N14957,N14958);
and and8903(N14967,N14969,N14970);
and and8904(N14968,N14971,N14972);
and and8911(N14981,N14983,N14984);
and and8912(N14982,N14985,N14986);
and and8919(N14995,N14997,N14998);
and and8920(N14996,N14999,N15000);
and and8927(N15009,N15011,N15012);
and and8928(N15010,N15013,N15014);
and and8935(N15023,N15025,N15026);
and and8936(N15024,N15027,N15028);
and and8943(N15037,N15039,N15040);
and and8944(N15038,N15041,N15042);
and and8951(N15051,N15053,N15054);
and and8952(N15052,N15055,N15056);
and and8959(N15065,N15067,N15068);
and and8960(N15066,N15069,N15070);
and and8967(N15079,N15081,N15082);
and and8968(N15080,N15083,N15084);
and and8975(N15093,N15095,N15096);
and and8976(N15094,N15097,N15098);
and and8983(N15107,N15109,N15110);
and and8984(N15108,N15111,N15112);
and and8991(N15121,N15123,N15124);
and and8992(N15122,N15125,N15126);
and and8999(N15135,N15137,N15138);
and and9000(N15136,N15139,N15140);
and and9007(N15149,N15151,N15152);
and and9008(N15150,N15153,N15154);
and and9015(N15163,N15165,N15166);
and and9016(N15164,N15167,N15168);
and and9023(N15177,N15179,N15180);
and and9024(N15178,N15181,N15182);
and and9031(N15191,N15193,N15194);
and and9032(N15192,N15195,N15196);
and and9039(N15204,N15206,N15207);
and and9040(N15205,N15208,N15209);
and and9047(N15217,N15219,N15220);
and and9048(N15218,N15221,N15222);
and and9055(N15230,N15232,N15233);
and and9056(N15231,N15234,N15235);
and and9063(N15243,N15245,N15246);
and and9064(N15244,N15247,N15248);
and and9071(N15256,N15258,N15259);
and and9072(N15257,N15260,N15261);
and and9079(N15269,N15271,N15272);
and and9080(N15270,N15273,N15274);
and and9087(N15282,N15284,N15285);
and and9088(N15283,N15286,N15287);
and and9095(N15295,N15297,N15298);
and and9096(N15296,N15299,N15300);
and and9103(N15308,N15310,N15311);
and and9104(N15309,N15312,N15313);
and and9111(N15321,N15323,N15324);
and and9112(N15322,N15325,N15326);
and and9119(N15334,N15336,N15337);
and and9120(N15335,N15338,N15339);
and and9127(N15347,N15349,N15350);
and and9128(N15348,N15351,N15352);
and and9135(N15360,N15362,N15363);
and and9136(N15361,N15364,N15365);
and and9143(N15373,N15375,N15376);
and and9144(N15374,N15377,N15378);
and and9151(N15386,N15388,N15389);
and and9152(N15387,N15390,N15391);
and and9159(N15399,N15401,N15402);
and and9160(N15400,N15403,N15404);
and and9167(N15412,N15414,N15415);
and and9168(N15413,N15416,N15417);
and and9175(N15425,N15427,N15428);
and and9176(N15426,N15429,N15430);
and and9183(N15438,N15440,N15441);
and and9184(N15439,N15442,N15443);
and and9191(N15451,N15453,N15454);
and and9192(N15452,N15455,N15456);
and and9199(N15464,N15466,N15467);
and and9200(N15465,N15468,N15469);
and and9207(N15477,N15479,N15480);
and and9208(N15478,N15481,N15482);
and and9215(N15490,N15492,N15493);
and and9216(N15491,N15494,N15495);
and and9223(N15503,N15505,N15506);
and and9224(N15504,N15507,N15508);
and and9231(N15516,N15518,N15519);
and and9232(N15517,N15520,N15521);
and and9239(N15529,N15531,N15532);
and and9240(N15530,N15533,N15534);
and and9247(N15542,N15544,N15545);
and and9248(N15543,N15546,N15547);
and and9255(N15555,N15557,N15558);
and and9256(N15556,N15559,N15560);
and and9263(N15568,N15570,N15571);
and and9264(N15569,N15572,N15573);
and and9271(N15581,N15583,N15584);
and and9272(N15582,N15585,N15586);
and and9279(N15594,N15596,N15597);
and and9280(N15595,N15598,N15599);
and and9287(N15607,N15609,N15610);
and and9288(N15608,N15611,N15612);
and and9295(N15620,N15622,N15623);
and and9296(N15621,N15624,N15625);
and and9303(N15633,N15635,N15636);
and and9304(N15634,N15637,N15638);
and and9311(N15646,N15648,N15649);
and and9312(N15647,N15650,N15651);
and and9319(N15659,N15661,N15662);
and and9320(N15660,N15663,N15664);
and and9327(N15672,N15674,N15675);
and and9328(N15673,N15676,N15677);
and and9335(N15685,N15687,N15688);
and and9336(N15686,N15689,N15690);
and and9343(N15698,N15700,N15701);
and and9344(N15699,N15702,N15703);
and and9351(N15711,N15713,N15714);
and and9352(N15712,N15715,N15716);
and and9359(N15724,N15726,N15727);
and and9360(N15725,N15728,N15729);
and and9367(N15737,N15739,N15740);
and and9368(N15738,N15741,N15742);
and and9375(N15750,N15752,N15753);
and and9376(N15751,N15754,N15755);
and and9383(N15763,N15765,N15766);
and and9384(N15764,N15767,N15768);
and and9391(N15776,N15778,N15779);
and and9392(N15777,N15780,N15781);
and and9399(N15789,N15791,N15792);
and and9400(N15790,N15793,N15794);
and and9407(N15802,N15804,N15805);
and and9408(N15803,N15806,N15807);
and and9415(N15815,N15817,N15818);
and and9416(N15816,N15819,N15820);
and and9423(N15827,N15829,N15830);
and and9424(N15828,N15831,N15832);
and and9431(N15839,N15841,N15842);
and and9432(N15840,N15843,N15844);
and and9439(N15851,N15853,N15854);
and and9440(N15852,N15855,N15856);
and and9447(N15863,N15865,N15866);
and and9448(N15864,N15867,N15868);
and and9455(N15875,N15877,N15878);
and and9456(N15876,N15879,N15880);
and and9463(N15887,N15889,N15890);
and and9464(N15888,N15891,N15892);
and and9471(N15899,N15901,N15902);
and and9472(N15900,N15903,N15904);
and and9479(N15911,N15913,N15914);
and and9480(N15912,N15915,N15916);
and and9487(N15923,N15925,N15926);
and and9488(N15924,N15927,N15928);
and and9495(N15935,N15937,N15938);
and and9496(N15936,N15939,N15940);
and and9503(N15947,N15949,N15950);
and and9504(N15948,N15951,N15952);
and and9511(N15959,N15961,N15962);
and and9512(N15960,N15963,N15964);
and and9519(N15971,N15973,N15974);
and and9520(N15972,N15975,N15976);
and and9527(N15983,N15985,N15986);
and and9528(N15984,N15987,N15988);
and and9535(N15995,N15997,N15998);
and and9536(N15996,N15999,N16000);
and and9543(N16007,N16009,N16010);
and and9544(N16008,N16011,N16012);
and and9551(N16019,N16021,N16022);
and and9552(N16020,N16023,N16024);
and and9559(N16031,N16033,N16034);
and and9560(N16032,N16035,N16036);
and and9567(N16043,N16045,N16046);
and and9568(N16044,N16047,N16048);
and and9575(N16055,N16057,N16058);
and and9576(N16056,N16059,N16060);
and and9583(N16067,N16069,N16070);
and and9584(N16068,N16071,N16072);
and and9591(N16079,N16081,N16082);
and and9592(N16080,N16083,N16084);
and and9599(N16091,N16093,N16094);
and and9600(N16092,N16095,N16096);
and and9607(N16103,N16105,N16106);
and and9608(N16104,N16107,N16108);
and and9615(N16115,N16117,N16118);
and and9616(N16116,N16119,N16120);
and and9623(N16127,N16129,N16130);
and and9624(N16128,N16131,N16132);
and and9631(N16139,N16141,N16142);
and and9632(N16140,N16143,N16144);
and and9639(N16151,N16153,N16154);
and and9640(N16152,N16155,N16156);
and and9647(N16163,N16165,N16166);
and and9648(N16164,N16167,N16168);
and and9655(N16175,N16177,N16178);
and and9656(N16176,N16179,N16180);
and and9663(N16187,N16189,N16190);
and and9664(N16188,N16191,N16192);
and and9671(N16199,N16201,N16202);
and and9672(N16200,N16203,N16204);
and and9679(N16211,N16213,N16214);
and and9680(N16212,N16215,N16216);
and and9687(N16223,N16225,N16226);
and and9688(N16224,N16227,N16228);
and and9695(N16235,N16237,N16238);
and and9696(N16236,N16239,N16240);
and and9703(N16247,N16249,N16250);
and and9704(N16248,N16251,N16252);
and and9711(N16259,N16261,N16262);
and and9712(N16260,N16263,N16264);
and and9719(N16271,N16273,N16274);
and and9720(N16272,N16275,N16276);
and and9727(N16283,N16285,N16286);
and and9728(N16284,N16287,N16288);
and and9735(N16295,N16297,N16298);
and and9736(N16296,N16299,N16300);
and and9743(N16307,N16309,N16310);
and and9744(N16308,N16311,N16312);
and and9751(N16319,N16321,N16322);
and and9752(N16320,N16323,N16324);
and and9759(N16331,N16333,N16334);
and and9760(N16332,N16335,N16336);
and and9767(N16343,N16345,N16346);
and and9768(N16344,N16347,N16348);
and and9775(N16355,N16357,N16358);
and and9776(N16356,N16359,N16360);
and and9783(N16367,N16369,N16370);
and and9784(N16368,N16371,N16372);
and and9791(N16379,N16381,N16382);
and and9792(N16380,N16383,N16384);
and and9799(N16391,N16393,N16394);
and and9800(N16392,N16395,N16396);
and and9807(N16403,N16405,N16406);
and and9808(N16404,N16407,N16408);
and and9815(N16415,N16417,N16418);
and and9816(N16416,N16419,N16420);
and and9823(N16427,N16429,N16430);
and and9824(N16428,N16431,N16432);
and and9831(N16439,N16441,N16442);
and and9832(N16440,N16443,N16444);
and and9839(N16451,N16453,N16454);
and and9840(N16452,N16455,N16456);
and and9847(N16462,N16464,N16465);
and and9848(N16463,N16466,N16467);
and and9855(N16473,N16475,N16476);
and and9856(N16474,N16477,N16478);
and and9863(N16484,N16486,N16487);
and and9864(N16485,N16488,N16489);
and and9871(N16495,N16497,N16498);
and and9872(N16496,N16499,N16500);
and and9879(N16506,N16508,N16509);
and and9880(N16507,N16510,N16511);
and and9887(N16517,N16519,N16520);
and and9888(N16518,N16521,N16522);
and and9895(N16528,N16530,N16531);
and and9896(N16529,N16532,N16533);
and and9903(N16539,N16541,N16542);
and and9904(N16540,N16543,N16544);
and and9911(N16550,N16552,N16553);
and and9912(N16551,N16554,N16555);
and and9919(N16561,N16563,N16564);
and and9920(N16562,N16565,N16566);
and and9927(N16572,N16574,N16575);
and and9928(N16573,N16576,N16577);
and and9935(N16583,N16585,N16586);
and and9936(N16584,N16587,N16588);
and and9943(N16594,N16596,N16597);
and and9944(N16595,N16598,N16599);
and and9951(N16605,N16607,N16608);
and and9952(N16606,N16609,N16610);
and and9959(N16616,N16618,N16619);
and and9960(N16617,N16620,N16621);
and and9967(N16627,N16629,N16630);
and and9968(N16628,N16631,N16632);
and and9975(N16638,N16640,N16641);
and and9976(N16639,N16642,N16643);
and and9983(N16649,N16651,N16652);
and and9984(N16650,N16653,N16654);
and and9991(N16660,N16662,N16663);
and and9992(N16661,N16664,N16665);
and and9999(N16671,N16673,N16674);
and and10000(N16672,N16675,N16676);
and and10007(N16682,N16684,N16685);
and and10008(N16683,N16686,N16687);
and and10015(N16693,N16695,N16696);
and and10016(N16694,N16697,N16698);
and and10023(N16704,N16706,N16707);
and and10024(N16705,N16708,N16709);
and and10031(N16715,N16717,N16718);
and and10032(N16716,N16719,N16720);
and and10039(N16726,N16728,N16729);
and and10040(N16727,N16730,N16731);
and and10047(N16737,N16739,N16740);
and and10048(N16738,N16741,N16742);
and and10055(N16748,N16750,N16751);
and and10056(N16749,N16752,N16753);
and and10063(N16759,N16761,N16762);
and and10064(N16760,N16763,N16764);
and and10071(N16770,N16772,N16773);
and and10072(N16771,N16774,N16775);
and and10079(N16781,N16783,N16784);
and and10080(N16782,N16785,N16786);
and and10087(N16792,N16794,N16795);
and and10088(N16793,N16796,N16797);
and and10095(N16803,N16805,N16806);
and and10096(N16804,N16807,N16808);
and and10103(N16814,N16816,N16817);
and and10104(N16815,N16818,N16819);
and and10111(N16825,N16827,N16828);
and and10112(N16826,N16829,N16830);
and and10119(N16836,N16838,N16839);
and and10120(N16837,N16840,N16841);
and and10127(N16847,N16849,N16850);
and and10128(N16848,N16851,N16852);
and and10135(N16858,N16860,N16861);
and and10136(N16859,N16862,N16863);
and and10143(N16869,N16871,N16872);
and and10144(N16870,N16873,N16874);
and and10151(N16880,N16882,N16883);
and and10152(N16881,N16884,N16885);
and and10159(N16891,N16893,N16894);
and and10160(N16892,N16895,N16896);
and and10167(N16901,N16903,N16904);
and and10168(N16902,N16905,N16906);
and and10175(N16911,N16913,N16914);
and and10176(N16912,N16915,N16916);
and and10183(N16921,N16923,N16924);
and and10184(N16922,N16925,N16926);
and and10191(N16931,N16933,N16934);
and and10192(N16932,N16935,N16936);
and and10199(N16941,N16943,N16944);
and and10200(N16942,N16945,N16946);
and and10207(N16951,N16953,N16954);
and and10208(N16952,N16955,N16956);
and and10215(N16961,N16963,N16964);
and and10216(N16962,N16965,N16966);
and and10223(N16971,N16973,N16974);
and and10224(N16972,N16975,N16976);
and and10231(N16981,N16983,N16984);
and and10232(N16982,N16985,N16986);
and and10239(N16991,N16993,N16994);
and and10240(N16992,N16995,N16996);
and and10247(N17001,N17003,N17004);
and and10248(N17002,N17005,N17006);
and and10255(N17011,N17013,N17014);
and and10256(N17012,N17015,N17016);
and and10263(N17021,N17023,N17024);
and and10264(N17022,N17025,N17026);
and and10271(N17031,N17033,N17034);
and and10272(N17032,N17035,N17036);
and and10279(N17041,N17043,N17044);
and and10280(N17042,N17045,N17046);
and and10287(N17051,N17053,N17054);
and and10288(N17052,N17055,N17056);
and and10295(N17061,N17063,N17064);
and and10296(N17062,N17065,N17066);
and and10303(N17070,N17072,N17073);
and and10304(N17071,N17074,N17075);
and and10311(N17079,N17081,N17082);
and and10312(N17080,N17083,N17084);
and and10319(N17088,N17090,N17091);
and and10320(N17089,N17092,N17093);
and and10327(N17097,N17099,N17100);
and and10328(N17098,N17101,N17102);
and and10335(N17106,N17108,N17109);
and and10336(N17107,N17110,N17111);
and and10343(N17115,N17117,N17118);
and and10344(N17116,N17119,N17120);
and and10351(N17124,N17126,N17127);
and and10352(N17125,N17128,N17129);
and and10359(N17133,N17135,N17136);
and and10360(N17134,N17137,N17138);
and and10367(N17142,N17144,N17145);
and and10368(N17143,N17146,N17147);
and and10375(N17151,N17153,N17154);
and and10376(N17152,N17155,N17156);
and and10383(N17159,N17161,N17162);
and and10384(N17160,N17163,N17164);
and and10390(N17173,N17175,N17176);
and and10391(N17174,N17177,N17178);
and and10397(N17187,N17189,N17190);
and and10398(N17188,N17191,N17192);
and and10404(N17201,N17203,N17204);
and and10405(N17202,N17205,N17206);
and and10411(N17215,N17217,N17218);
and and10412(N17216,N17219,N17220);
and and10418(N17228,N17230,N17231);
and and10419(N17229,N17232,N17233);
and and10425(N17241,N17243,N17244);
and and10426(N17242,N17245,N17246);
and and10432(N17254,N17256,N17257);
and and10433(N17255,N17258,N17259);
and and10439(N17267,N17269,N17270);
and and10440(N17268,N17271,N17272);
and and10446(N17280,N17282,N17283);
and and10447(N17281,N17284,N17285);
and and10453(N17292,N17294,N17295);
and and10454(N17293,N17296,N17297);
and and10460(N17304,N17306,N17307);
and and10461(N17305,N17308,N17309);
and and10467(N17316,N17318,N17319);
and and10468(N17317,N17320,N17321);
and and10474(N17328,N17330,N17331);
and and10475(N17329,N17332,N17333);
and and10481(N17340,N17342,N17343);
and and10482(N17341,N17344,N17345);
and and10488(N17352,N17354,N17355);
and and10489(N17353,N17356,N17357);
and and10495(N17364,N17366,N17367);
and and10496(N17365,N17368,N17369);
and and10502(N17376,N17378,N17379);
and and10503(N17377,N17380,N17381);
and and10509(N17388,N17390,N17391);
and and10510(N17389,N17392,N17393);
and and10516(N17399,N17401,N17402);
and and10517(N17400,N17403,N17404);
and and10523(N17410,N17412,N17413);
and and10524(N17411,N17414,N17415);
and and10530(N17421,N17423,N17424);
and and10531(N17422,N17425,N17426);
and and10537(N17432,N17434,N17435);
and and10538(N17433,N17436,N17437);
and and10544(N17443,N17445,N17446);
and and10545(N17444,N17447,N17448);
and and10551(N17454,N17456,N17457);
and and10552(N17455,N17458,N17459);
and and10558(N17465,N17467,N17468);
and and10559(N17466,N17469,N17470);
and and10565(N17476,N17478,N17479);
and and10566(N17477,N17480,N17481);
and and10572(N17487,N17489,N17490);
and and10573(N17488,N17491,N17492);
and and10579(N17498,N17500,N17501);
and and10580(N17499,N17502,N17503);
and and10586(N17509,N17511,N17512);
and and10587(N17510,N17513,N17514);
and and10593(N17520,N17522,N17523);
and and10594(N17521,N17524,N17525);
and and10600(N17531,N17533,N17534);
and and10601(N17532,N17535,N17536);
and and10607(N17542,N17544,N17545);
and and10608(N17543,N17546,N17547);
and and10614(N17553,N17555,N17556);
and and10615(N17554,N17557,N17558);
and and10621(N17564,N17566,N17567);
and and10622(N17565,N17568,N17569);
and and10628(N17575,N17577,N17578);
and and10629(N17576,N17579,N17580);
and and10635(N17585,N17587,N17588);
and and10636(N17586,N17589,N17590);
and and10642(N17595,N17597,N17598);
and and10643(N17596,N17599,N17600);
and and10649(N17605,N17607,N17608);
and and10650(N17606,N17609,N17610);
and and10656(N17615,N17617,N17618);
and and10657(N17616,N17619,N17620);
and and10663(N17625,N17627,N17628);
and and10664(N17626,N17629,N17630);
and and10670(N17635,N17637,N17638);
and and10671(N17636,N17639,N17640);
and and6903(N11885,N11889,N11890);
and and6904(N11886,N11891,in2);
and and6905(N11887,N11892,N11893);
and and6906(N11888,N11894,N11895);
and and6912(N11903,N11907,N11908);
and and6913(N11904,N11909,N11910);
and and6914(N11905,N11911,N11912);
and and6915(N11906,N11913,N11914);
and and6921(N11921,N11925,N11926);
and and6922(N11922,N11927,N11928);
and and6923(N11923,N11929,N11930);
and and6924(N11924,N11931,R3);
and and6930(N11938,N11942,N11943);
and and6931(N11939,N11944,N11945);
and and6932(N11940,N11946,R0);
and and6933(N11941,N11947,N11948);
and and6939(N11955,N11959,N11960);
and and6940(N11956,N11961,in1);
and and6941(N11957,N11962,N11963);
and and6942(N11958,N11964,N11965);
and and6948(N11972,N11976,N11977);
and and6949(N11973,N11978,N11979);
and and6950(N11974,N11980,N11981);
and and6951(N11975,R1,N11982);
and and6957(N11989,N11993,N11994);
and and6958(N11990,in0,in2);
and and6959(N11991,N11995,R1);
and and6960(N11992,N11996,N11997);
and and6966(N12005,N12009,N12010);
and and6967(N12006,N12011,in2);
and and6968(N12007,N12012,N12013);
and and6969(N12008,N12014,N12015);
and and6975(N12021,N12025,N12026);
and and6976(N12022,N12027,in1);
and and6977(N12023,N12028,N12029);
and and6978(N12024,N12030,R3);
and and6984(N12037,N12041,N12042);
and and6985(N12038,N12043,N12044);
and and6986(N12039,N12045,R0);
and and6987(N12040,N12046,N12047);
and and6993(N12053,N12057,N12058);
and and6994(N12054,N12059,N12060);
and and6995(N12055,N12061,N12062);
and and6996(N12056,N12063,R3);
and and7002(N12069,N12073,N12074);
and and7003(N12070,N12075,N12076);
and and7004(N12071,N12077,N12078);
and and7005(N12072,N12079,R3);
and and7011(N12085,N12089,N12090);
and and7012(N12086,N12091,N12092);
and and7013(N12087,R0,N12093);
and and7014(N12088,N12094,N12095);
and and7020(N12101,N12105,N12106);
and and7021(N12102,N12107,N12108);
and and7022(N12103,in2,N12109);
and and7023(N12104,R1,N12110);
and and7029(N12117,N12121,N12122);
and and7030(N12118,N12123,N12124);
and and7031(N12119,N12125,N12126);
and and7032(N12120,N12127,R3);
and and7038(N12133,N12137,N12138);
and and7039(N12134,N12139,N12140);
and and7040(N12135,in2,R0);
and and7041(N12136,N12141,N12142);
and and7047(N12149,N12153,N12154);
and and7048(N12150,N12155,N12156);
and and7049(N12151,N12157,R1);
and and7050(N12152,R2,N12158);
and and7056(N12165,N12169,N12170);
and and7057(N12166,N12171,N12172);
and and7058(N12167,in2,R0);
and and7059(N12168,N12173,N12174);
and and7065(N12181,N12185,N12186);
and and7066(N12182,N12187,N12188);
and and7067(N12183,N12189,N12190);
and and7068(N12184,R2,R3);
and and7074(N12197,N12201,N12202);
and and7075(N12198,N12203,N12204);
and and7076(N12199,N12205,R1);
and and7077(N12200,R2,R3);
and and7083(N12212,N12216,N12217);
and and7084(N12213,N12218,N12219);
and and7085(N12214,in2,N12220);
and and7086(N12215,R1,R3);
and and7092(N12227,N12231,N12232);
and and7093(N12228,N12233,N12234);
and and7094(N12229,R0,R1);
and and7095(N12230,N12235,R3);
and and7101(N12242,N12246,N12247);
and and7102(N12243,in0,in2);
and and7103(N12244,N12248,N12249);
and and7104(N12245,N12250,R3);
and and7110(N12257,N12261,N12262);
and and7111(N12258,N12263,N12264);
and and7112(N12259,N12265,R1);
and and7113(N12260,N12266,R3);
and and7119(N12272,N12276,N12277);
and and7120(N12273,in1,N12278);
and and7121(N12274,R0,N12279);
and and7122(N12275,R2,N12280);
and and7128(N12287,N12291,N12292);
and and7129(N12288,N12293,N12294);
and and7130(N12289,in2,R0);
and and7131(N12290,N12295,R3);
and and7137(N12302,N12306,N12307);
and and7138(N12303,in0,N12308);
and and7139(N12304,N12309,N12310);
and and7140(N12305,N12311,R3);
and and7146(N12317,N12321,N12322);
and and7147(N12318,N12323,in2);
and and7148(N12319,N12324,N12325);
and and7149(N12320,N12326,R3);
and and7155(N12332,N12336,N12337);
and and7156(N12333,in1,N12338);
and and7157(N12334,N12339,N12340);
and and7158(N12335,N12341,R3);
and and7164(N12347,N12351,N12352);
and and7165(N12348,N12353,N12354);
and and7166(N12349,R0,R1);
and and7167(N12350,N12355,R3);
and and7173(N12362,N12366,N12367);
and and7174(N12363,in0,in1);
and and7175(N12364,N12368,N12369);
and and7176(N12365,R2,N12370);
and and7182(N12377,N12381,N12382);
and and7183(N12378,in1,in2);
and and7184(N12379,N12383,N12384);
and and7185(N12380,R2,R3);
and and7191(N12392,N12396,N12397);
and and7192(N12393,in1,N12398);
and and7193(N12394,R0,N12399);
and and7194(N12395,N12400,R3);
and and7200(N12407,N12411,N12412);
and and7201(N12408,in0,N12413);
and and7202(N12409,N12414,N12415);
and and7203(N12410,R2,R3);
and and7209(N12422,N12426,N12427);
and and7210(N12423,in1,N12428);
and and7211(N12424,N12429,N12430);
and and7212(N12425,R2,R3);
and and7218(N12437,N12441,N12442);
and and7219(N12438,N12443,in2);
and and7220(N12439,N12444,N12445);
and and7221(N12440,R2,R3);
and and7227(N12452,N12456,N12457);
and and7228(N12453,N12458,N12459);
and and7229(N12454,N12460,N12461);
and and7230(N12455,R2,R3);
and and7236(N12467,N12471,N12472);
and and7237(N12468,N12473,N12474);
and and7238(N12469,N12475,N12476);
and and7239(N12470,R1,R2);
and and7245(N12482,N12486,N12487);
and and7246(N12483,N12488,N12489);
and and7247(N12484,N12490,R0);
and and7248(N12485,N12491,R2);
and and7254(N12497,N12501,N12502);
and and7255(N12498,in1,N12503);
and and7256(N12499,N12504,N12505);
and and7257(N12500,N12506,R3);
and and7263(N12512,N12516,N12517);
and and7264(N12513,N12518,N12519);
and and7265(N12514,N12520,N12521);
and and7266(N12515,R2,R3);
and and7272(N12527,N12531,N12532);
and and7273(N12528,N12533,N12534);
and and7274(N12529,N12535,R1);
and and7275(N12530,N12536,R3);
and and7281(N12542,N12546,N12547);
and and7282(N12543,N12548,in1);
and and7283(N12544,R0,N12549);
and and7284(N12545,N12550,N12551);
and and7290(N12557,N12561,N12562);
and and7291(N12558,in0,N12563);
and and7292(N12559,N12564,R0);
and and7293(N12560,N12565,N12566);
and and7299(N12572,N12576,N12577);
and and7300(N12573,N12578,in1);
and and7301(N12574,N12579,R0);
and and7302(N12575,N12580,R2);
and and7308(N12587,N12591,N12592);
and and7309(N12588,in0,N12593);
and and7310(N12589,N12594,N12595);
and and7311(N12590,N12596,R3);
and and7317(N12602,N12606,N12607);
and and7318(N12603,N12608,in1);
and and7319(N12604,R0,N12609);
and and7320(N12605,N12610,N12611);
and and7326(N12617,N12621,N12622);
and and7327(N12618,in0,N12623);
and and7328(N12619,R0,N12624);
and and7329(N12620,N12625,N12626);
and and7335(N12632,N12636,N12637);
and and7336(N12633,N12638,N12639);
and and7337(N12634,N12640,R0);
and and7338(N12635,R1,N12641);
and and7344(N12647,N12651,N12652);
and and7345(N12648,in0,N12653);
and and7346(N12649,R0,N12654);
and and7347(N12650,N12655,R3);
and and7353(N12662,N12666,N12667);
and and7354(N12663,N12668,N12669);
and and7355(N12664,in2,R0);
and and7356(N12665,N12670,R3);
and and7362(N12677,N12681,N12682);
and and7363(N12678,N12683,N12684);
and and7364(N12679,N12685,R1);
and and7365(N12680,N12686,R3);
and and7371(N12692,N12696,N12697);
and and7372(N12693,in0,in1);
and and7373(N12694,N12698,R0);
and and7374(N12695,N12699,N12700);
and and7380(N12707,N12711,N12712);
and and7381(N12708,in0,in1);
and and7382(N12709,N12713,N12714);
and and7383(N12710,R1,N12715);
and and7389(N12722,N12726,N12727);
and and7390(N12723,N12728,N12729);
and and7391(N12724,in2,R1);
and and7392(N12725,R2,N12730);
and and7398(N12737,N12741,N12742);
and and7399(N12738,in1,N12743);
and and7400(N12739,N12744,R1);
and and7401(N12740,R2,N12745);
and and7407(N12752,N12756,N12757);
and and7408(N12753,in1,N12758);
and and7409(N12754,R0,N12759);
and and7410(N12755,N12760,R3);
and and7416(N12766,N12770,N12771);
and and7417(N12767,N12772,in2);
and and7418(N12768,R0,N12773);
and and7419(N12769,R2,N12774);
and and7425(N12780,N12784,N12785);
and and7426(N12781,in1,N12786);
and and7427(N12782,R0,N12787);
and and7428(N12783,R2,N12788);
and and7434(N12794,N12798,N12799);
and and7435(N12795,in0,N12800);
and and7436(N12796,in2,R0);
and and7437(N12797,N12801,N12802);
and and7443(N12808,N12812,N12813);
and and7444(N12809,in0,in1);
and and7445(N12810,R0,N12814);
and and7446(N12811,N12815,R3);
and and7452(N12822,N12826,N12827);
and and7453(N12823,N12828,in1);
and and7454(N12824,in2,N12829);
and and7455(N12825,R1,N12830);
and and7461(N12836,N12840,N12841);
and and7462(N12837,N12842,N12843);
and and7463(N12838,in2,R0);
and and7464(N12839,N12844,R3);
and and7470(N12850,N12854,N12855);
and and7471(N12851,N12856,N12857);
and and7472(N12852,N12858,R0);
and and7473(N12853,N12859,R3);
and and7479(N12864,N12868,N12869);
and and7480(N12865,N12870,in1);
and and7481(N12866,N12871,R0);
and and7482(N12867,R1,N12872);
and and7488(N12878,N12882,N12883);
and and7489(N12879,N12884,N12885);
and and7490(N12880,in2,R0);
and and7491(N12881,R1,N12886);
and and7497(N12892,N12896,N12897);
and and7498(N12893,N12898,in2);
and and7499(N12894,N12899,N12900);
and and7500(N12895,R2,R3);
and and7506(N12906,N12910,N12911);
and and7507(N12907,in0,in1);
and and7508(N12908,in2,R0);
and and7509(N12909,N12912,N12913);
and and7515(N12920,N12924,N12925);
and and7516(N12921,N12926,in1);
and and7517(N12922,R0,N12927);
and and7518(N12923,N12928,R3);
and and7524(N12934,N12938,N12939);
and and7525(N12935,in1,N12940);
and and7526(N12936,N12941,N12942);
and and7527(N12937,R2,N12943);
and and7533(N12948,N12952,N12953);
and and7534(N12949,N12954,in2);
and and7535(N12950,N12955,N12956);
and and7536(N12951,R2,N12957);
and and7542(N12962,N12966,N12967);
and and7543(N12963,in0,in2);
and and7544(N12964,R0,N12968);
and and7545(N12965,N12969,N12970);
and and7551(N12976,N12980,N12981);
and and7552(N12977,N12982,in1);
and and7553(N12978,in2,R0);
and and7554(N12979,N12983,N12984);
and and7560(N12990,N12994,N12995);
and and7561(N12991,in1,in2);
and and7562(N12992,N12996,N12997);
and and7563(N12993,N12998,R3);
and and7569(N13004,N13008,N13009);
and and7570(N13005,in0,in1);
and and7571(N13006,N13010,N13011);
and and7572(N13007,N13012,N13013);
and and7578(N13018,N13022,N13023);
and and7579(N13019,N13024,in2);
and and7580(N13020,N13025,R1);
and and7581(N13021,R2,R3);
and and7587(N13032,N13036,N13037);
and and7588(N13033,N13038,in1);
and and7589(N13034,in2,R0);
and and7590(N13035,N13039,R3);
and and7596(N13046,N13050,N13051);
and and7597(N13047,N13052,N13053);
and and7598(N13048,N13054,R1);
and and7599(N13049,R2,R3);
and and7605(N13060,N13064,N13065);
and and7606(N13061,N13066,in1);
and and7607(N13062,R0,R1);
and and7608(N13063,N13067,N13068);
and and7614(N13074,N13078,N13079);
and and7615(N13075,in0,N13080);
and and7616(N13076,N13081,N13082);
and and7617(N13077,R2,N13083);
and and7623(N13088,N13092,N13093);
and and7624(N13089,N13094,N13095);
and and7625(N13090,in2,N13096);
and and7626(N13091,N13097,R2);
and and7632(N13102,N13106,N13107);
and and7633(N13103,in0,in2);
and and7634(N13104,N13108,R1);
and and7635(N13105,N13109,N13110);
and and7641(N13116,N13120,N13121);
and and7642(N13117,N13122,in1);
and and7643(N13118,in2,N13123);
and and7644(N13119,R1,N13124);
and and7650(N13130,N13134,N13135);
and and7651(N13131,in0,in2);
and and7652(N13132,N13136,R1);
and and7653(N13133,R2,N13137);
and and7659(N13144,N13148,N13149);
and and7660(N13145,in0,N13150);
and and7661(N13146,N13151,R0);
and and7662(N13147,N13152,R2);
and and7668(N13158,N13162,N13163);
and and7669(N13159,N13164,N13165);
and and7670(N13160,in2,R0);
and and7671(N13161,N13166,R2);
and and7677(N13172,N13176,N13177);
and and7678(N13173,N13178,N13179);
and and7679(N13174,N13180,R1);
and and7680(N13175,R2,N13181);
and and7686(N13186,N13190,N13191);
and and7687(N13187,N13192,in1);
and and7688(N13188,in2,R0);
and and7689(N13189,R1,N13193);
and and7695(N13200,N13204,N13205);
and and7696(N13201,in1,N13206);
and and7697(N13202,N13207,R1);
and and7698(N13203,R2,N13208);
and and7704(N13214,N13218,N13219);
and and7705(N13215,in0,N13220);
and and7706(N13216,N13221,R0);
and and7707(N13217,N13222,R2);
and and7713(N13228,N13232,N13233);
and and7714(N13229,in0,N13234);
and and7715(N13230,N13235,N13236);
and and7716(N13231,N13237,R2);
and and7722(N13242,N13246,N13247);
and and7723(N13243,N13248,in1);
and and7724(N13244,N13249,N13250);
and and7725(N13245,N13251,R2);
and and7731(N13256,N13260,N13261);
and and7732(N13257,N13262,N13263);
and and7733(N13258,in2,R0);
and and7734(N13259,N13264,N13265);
and and7740(N13270,N13274,N13275);
and and7741(N13271,N13276,in1);
and and7742(N13272,N13277,R0);
and and7743(N13273,R1,N13278);
and and7749(N13284,N13288,N13289);
and and7750(N13285,in0,in1);
and and7751(N13286,N13290,N13291);
and and7752(N13287,R2,N13292);
and and7758(N13298,N13302,N13303);
and and7759(N13299,N13304,in1);
and and7760(N13300,N13305,R0);
and and7761(N13301,N13306,R3);
and and7767(N13312,N13316,N13317);
and and7768(N13313,in1,N13318);
and and7769(N13314,N13319,N13320);
and and7770(N13315,R2,R3);
and and7776(N13326,N13330,N13331);
and and7777(N13327,in1,in2);
and and7778(N13328,N13332,R1);
and and7779(N13329,R2,R3);
and and7785(N13339,N13343,N13344);
and and7786(N13340,in0,in2);
and and7787(N13341,R0,R1);
and and7788(N13342,N13345,R3);
and and7794(N13352,N13356,N13357);
and and7795(N13353,in1,in2);
and and7796(N13354,R0,N13358);
and and7797(N13355,N13359,R3);
and and7803(N13365,N13369,N13370);
and and7804(N13366,in0,in2);
and and7805(N13367,R0,N13371);
and and7806(N13368,R2,R3);
and and7812(N13378,N13382,N13383);
and and7813(N13379,in0,in1);
and and7814(N13380,N13384,R0);
and and7815(N13381,N13385,R2);
and and7821(N13391,N13395,N13396);
and and7822(N13392,N13397,in1);
and and7823(N13393,N13398,R1);
and and7824(N13394,R2,R3);
and and7830(N13404,N13408,N13409);
and and7831(N13405,in0,in2);
and and7832(N13406,R0,N13410);
and and7833(N13407,R2,R3);
and and7839(N13417,N13421,N13422);
and and7840(N13418,in0,in1);
and and7841(N13419,in2,N13423);
and and7842(N13420,N13424,R3);
and and7848(N13430,N13434,N13435);
and and7849(N13431,in0,in1);
and and7850(N13432,in2,R0);
and and7851(N13433,R1,R2);
and and7857(N13443,N13447,N13448);
and and7858(N13444,in1,N13449);
and and7859(N13445,R0,N13450);
and and7860(N13446,N13451,R3);
and and7866(N13456,N13460,N13461);
and and7867(N13457,in0,in1);
and and7868(N13458,in2,N13462);
and and7869(N13459,N13463,R2);
and and7875(N13469,N13473,N13474);
and and7876(N13470,in0,in1);
and and7877(N13471,N13475,N13476);
and and7878(N13472,R1,R2);
and and7884(N13482,N13486,N13487);
and and7885(N13483,in1,in2);
and and7886(N13484,R0,R1);
and and7887(N13485,N13488,N13489);
and and7893(N13495,N13499,N13500);
and and7894(N13496,in1,N13501);
and and7895(N13497,N13502,R1);
and and7896(N13498,R2,R3);
and and7902(N13508,N13512,N13513);
and and7903(N13509,in1,in2);
and and7904(N13510,N13514,R1);
and and7905(N13511,R2,N13515);
and and7911(N13521,N13525,N13526);
and and7912(N13522,in0,in1);
and and7913(N13523,N13527,N13528);
and and7914(N13524,R1,R2);
and and7920(N13534,N13538,N13539);
and and7921(N13535,in0,in1);
and and7922(N13536,N13540,R1);
and and7923(N13537,N13541,N13542);
and and7929(N13547,N13551,N13552);
and and7930(N13548,in0,in1);
and and7931(N13549,N13553,N13554);
and and7932(N13550,N13555,R2);
and and7938(N13560,N13564,N13565);
and and7939(N13561,N13566,in1);
and and7940(N13562,in2,N13567);
and and7941(N13563,R2,R3);
and and7947(N13573,N13577,N13578);
and and7948(N13574,N13579,in1);
and and7949(N13575,N13580,R0);
and and7950(N13576,R1,N13581);
and and7956(N13586,N13590,N13591);
and and7957(N13587,N13592,N13593);
and and7958(N13588,R0,R1);
and and7959(N13589,R2,R3);
and and7965(N13599,N13603,N13604);
and and7966(N13600,in0,in1);
and and7967(N13601,in2,N13605);
and and7968(N13602,N13606,R3);
and and7974(N13612,N13616,N13617);
and and7975(N13613,N13618,in2);
and and7976(N13614,R0,R1);
and and7977(N13615,R2,N13619);
and and7983(N13625,N13629,N13630);
and and7984(N13626,N13631,in1);
and and7985(N13627,in2,R1);
and and7986(N13628,R2,R3);
and and7992(N13638,N13642,N13643);
and and7993(N13639,N13644,in2);
and and7994(N13640,R0,R1);
and and7995(N13641,N13645,N13646);
and and8001(N13651,N13655,N13656);
and and8002(N13652,in0,in1);
and and8003(N13653,in2,R0);
and and8004(N13654,N13657,N13658);
and and8010(N13664,N13668,N13669);
and and8011(N13665,in0,N13670);
and and8012(N13666,N13671,R0);
and and8013(N13667,R2,R3);
and and8019(N13677,N13681,N13682);
and and8020(N13678,N13683,in2);
and and8021(N13679,R0,N13684);
and and8022(N13680,R2,R3);
and and8028(N13690,N13694,N13695);
and and8029(N13691,N13696,in1);
and and8030(N13692,N13697,R0);
and and8031(N13693,R1,R2);
and and8037(N13703,N13707,N13708);
and and8038(N13704,in0,in1);
and and8039(N13705,N13709,N13710);
and and8040(N13706,N13711,R2);
and and8046(N13716,N13720,N13721);
and and8047(N13717,in0,N13722);
and and8048(N13718,N13723,N13724);
and and8049(N13719,R1,R3);
and and8055(N13729,N13733,N13734);
and and8056(N13730,N13735,N13736);
and and8057(N13731,in2,N13737);
and and8058(N13732,R1,N13738);
and and8064(N13742,N13746,N13747);
and and8065(N13743,in0,in1);
and and8066(N13744,N13748,R0);
and and8067(N13745,R2,R3);
and and8073(N13755,N13759,N13760);
and and8074(N13756,N13761,in1);
and and8075(N13757,in2,R0);
and and8076(N13758,N13762,R2);
and and8082(N13768,N13772,N13773);
and and8083(N13769,in0,in1);
and and8084(N13770,in2,N13774);
and and8085(N13771,R2,R3);
and and8091(N13781,N13785,N13786);
and and8092(N13782,in0,N13787);
and and8093(N13783,in2,R0);
and and8094(N13784,N13788,R2);
and and8100(N13794,N13798,N13799);
and and8101(N13795,in0,in1);
and and8102(N13796,N13800,R0);
and and8103(N13797,R1,R2);
and and8109(N13807,N13811,N13812);
and and8110(N13808,N13813,in1);
and and8111(N13809,in2,R1);
and and8112(N13810,R2,N13814);
and and8118(N13820,N13824,N13825);
and and8119(N13821,in0,in2);
and and8120(N13822,N13826,N13827);
and and8121(N13823,R2,R3);
and and8127(N13833,N13837,N13838);
and and8128(N13834,in0,in1);
and and8129(N13835,N13839,N13840);
and and8130(N13836,R2,R3);
and and8136(N13846,N13850,N13851);
and and8137(N13847,N13852,in1);
and and8138(N13848,in2,N13853);
and and8139(N13849,R2,R3);
and and8145(N13859,N13863,N13864);
and and8146(N13860,N13865,in1);
and and8147(N13861,N13866,R0);
and and8148(N13862,R1,R2);
and and8154(N13872,N13876,N13877);
and and8155(N13873,N13878,in1);
and and8156(N13874,in2,R0);
and and8157(N13875,R1,N13879);
and and8163(N13885,N13889,N13890);
and and8164(N13886,in0,N13891);
and and8165(N13887,R0,N13892);
and and8166(N13888,R2,R3);
and and8172(N13898,N13902,N13903);
and and8173(N13899,in0,in2);
and and8174(N13900,N13904,N13905);
and and8175(N13901,R2,R3);
and and8181(N13911,N13915,N13916);
and and8182(N13912,N13917,in1);
and and8183(N13913,in2,N13918);
and and8184(N13914,R2,R3);
and and8190(N13924,N13928,N13929);
and and8191(N13925,in0,in1);
and and8192(N13926,N13930,N13931);
and and8193(N13927,R1,R2);
and and8199(N13936,N13940,N13941);
and and8200(N13937,in0,in2);
and and8201(N13938,N13942,R1);
and and8202(N13939,R2,R3);
and and8208(N13948,N13952,N13953);
and and8209(N13949,in0,in1);
and and8210(N13950,in2,N13954);
and and8211(N13951,R1,R3);
and and8217(N13960,N13964,N13965);
and and8218(N13961,in0,in1);
and and8219(N13962,in2,R0);
and and8220(N13963,R2,N13966);
and and8226(N13972,N13976,N13977);
and and8227(N13973,in0,in1);
and and8228(N13974,in2,R1);
and and8229(N13975,R2,R3);
and and8235(N13984,N13988,N13989);
and and8236(N13985,in0,N13990);
and and8237(N13986,R0,R1);
and and8238(N13987,R2,N13991);
and and8244(N13996,N14000,N14001);
and and8245(N13997,in1,in2);
and and8246(N13998,R0,N14002);
and and8247(N13999,N14003,R3);
and and8253(N14008,N14012,N14013);
and and8254(N14009,N14014,in2);
and and8255(N14010,R0,R1);
and and8256(N14011,R2,R3);
and and8262(N14020,N14024,N14025);
and and8263(N14021,in1,N14026);
and and8264(N14022,R0,R1);
and and8265(N14023,R2,R3);
and and8271(N14032,N14036,N14037);
and and8272(N14033,in0,N14038);
and and8273(N14034,N14039,R0);
and and8274(N14035,R1,R2);
and and8280(N14044,N14048,N14049);
and and8281(N14045,in1,N14050);
and and8282(N14046,N14051,N14052);
and and8283(N14047,R2,R3);
and and8289(N14056,N14060,N14061);
and and8290(N14057,in0,N14062);
and and8291(N14058,N14063,R0);
and and8292(N14059,R2,R3);
and and8298(N14068,N14072,N14073);
and and8299(N14069,N14074,N14075);
and and8300(N14070,R0,R1);
and and8301(N14071,R2,N14076);
and and8307(N14080,N14084,N14085);
and and8308(N14081,in0,N14086);
and and8309(N14082,R0,R1);
and and8310(N14083,R2,R3);
and and8316(N14092,N14096,N14097);
and and8317(N14093,N14098,in1);
and and8318(N14094,in2,N14099);
and and8319(N14095,R1,R2);
and and8325(N14104,N14108,N14109);
and and8326(N14105,in0,in1);
and and8327(N14106,N14110,N14111);
and and8328(N14107,R1,R2);
and and8334(N14116,N14120,N14121);
and and8335(N14117,in0,N14122);
and and8336(N14118,in2,R0);
and and8337(N14119,R1,R3);
and and8343(N14128,N14132,N14133);
and and8344(N14129,in1,in2);
and and8345(N14130,R0,R1);
and and8346(N14131,N14134,R3);
and and8352(N14140,N14144,N14145);
and and8353(N14141,in0,N14146);
and and8354(N14142,R0,R1);
and and8355(N14143,R2,N14147);
and and8361(N14152,N14156,N14157);
and and8362(N14153,in1,N14158);
and and8363(N14154,R0,R1);
and and8364(N14155,R2,N14159);
and and8370(N14164,N14168,N14169);
and and8371(N14165,in0,in2);
and and8372(N14166,R0,N14170);
and and8373(N14167,R2,N14171);
and and8379(N14176,N14180,N14181);
and and8380(N14177,in0,in1);
and and8381(N14178,N14182,R0);
and and8382(N14179,N14183,R2);
and and8388(N14188,N14192,N14193);
and and8389(N14189,in1,N14194);
and and8390(N14190,R0,N14195);
and and8391(N14191,R2,R3);
and and8397(N14200,N14204,N14205);
and and8398(N14201,in0,in1);
and and8399(N14202,N14206,N14207);
and and8400(N14203,R1,N14208);
and and8406(N14212,N14216,N14217);
and and8407(N14213,in1,N14218);
and and8408(N14214,N14219,R1);
and and8409(N14215,R2,R3);
and and8415(N14224,N14228,N14229);
and and8416(N14225,in0,in1);
and and8417(N14226,in2,R0);
and and8418(N14227,R1,N14230);
and and8424(N14236,N14240,N14241);
and and8425(N14237,N14242,in1);
and and8426(N14238,in2,N14243);
and and8427(N14239,R1,R2);
and and8433(N14248,N14252,N14253);
and and8434(N14249,N14254,N14255);
and and8435(N14250,in2,R0);
and and8436(N14251,R1,R2);
and and8442(N14260,N14264,N14265);
and and8443(N14261,in0,in1);
and and8444(N14262,in2,R0);
and and8445(N14263,R1,R2);
and and8451(N14271,N14275,N14276);
and and8452(N14272,in0,in1);
and and8453(N14273,in2,N14277);
and and8454(N14274,R1,R2);
and and8460(N14282,N14286,N14287);
and and8461(N14283,in0,in1);
and and8462(N14284,R0,R1);
and and8463(N14285,R2,R3);
and and8469(N14293,N14297,N14298);
and and8470(N14294,in0,in1);
and and8471(N14295,in2,N14299);
and and8472(N14296,R2,R3);
and and8478(N14304,N14308,N14309);
and and8479(N14305,in0,in1);
and and8480(N14306,in2,R0);
and and8481(N14307,R2,R3);
and and8487(N14315,N14319,N14320);
and and8488(N14316,in0,in1);
and and8489(N14317,in2,N14321);
and and8490(N14318,N14322,R2);
and and8496(N14326,N14330,N14331);
and and8497(N14327,in0,in1);
and and8498(N14328,in2,R0);
and and8499(N14329,N14332,R3);
and and8505(N14337,N14341,N14342);
and and8506(N14338,in0,in1);
and and8507(N14339,in2,R1);
and and8508(N14340,R2,R3);
and and8514(N14348,N14352,N14353);
and and8515(N14349,in1,in2);
and and8516(N14350,R0,R1);
and and8517(N14351,R2,R3);
and and8523(N14359,N14363,N14364);
and and8524(N14360,in0,N14365);
and and8525(N14361,R0,R1);
and and8526(N14362,R2,R3);
and and8532(N14370,N14374,N14375);
and and8533(N14371,in0,in1);
and and8534(N14372,in2,R0);
and and8535(N14373,R1,N14376);
and and8541(N14381,N14385,N14386);
and and8542(N14382,in0,in1);
and and8543(N14383,in2,R0);
and and8544(N14384,N14387,R2);
and and8550(N14392,N14396,N14397);
and and8551(N14393,N14398,in1);
and and8552(N14394,in2,R0);
and and8553(N14395,R1,R2);
and and8559(N14403,N14407,N14408);
and and8560(N14404,in0,in1);
and and8561(N14405,N14409,R0);
and and8562(N14406,N14410,R2);
and and8568(N14414,N14418,N14419);
and and8569(N14415,in0,in1);
and and8570(N14416,in2,R0);
and and8571(N14417,R1,R2);
and and8577(N14425,N14429,N14430);
and and8578(N14426,in0,in1);
and and8579(N14427,in2,R0);
and and8580(N14428,N14431,R2);
and and8586(N14436,N14440,N14441);
and and8587(N14437,in0,in2);
and and8588(N14438,R0,R1);
and and8589(N14439,R2,R3);
and and8595(N14446,N14450,N14451);
and and8596(N14447,in0,N14452);
and and8597(N14448,in2,R0);
and and8598(N14449,R1,R2);
and and8604(N14456,N14460,N14461);
and and8605(N14457,in0,in1);
and and8606(N14458,R0,R1);
and and8607(N14459,R2,N14462);
and and8613(N14466,N14470,N14471);
and and8614(N14467,in0,in1);
and and8615(N14468,in2,R0);
and and8616(N14469,R1,R2);
and and8622(N14476,N14480,N14481);
and and8623(N14477,N14482,in1);
and and8624(N14478,in2,R1);
and and8625(N14479,R2,R3);
and and8631(N14486,N14490,N14491);
and and8632(N14487,in0,in1);
and and8633(N14488,in2,R1);
and and8634(N14489,R2,R3);
and and8640(N14496,N14500,N14501);
and and8641(N14497,in0,in1);
and and8642(N14498,in2,R0);
and and8643(N14499,R1,R2);
and and8649(N14505,N14509,in0);
and and8650(N14506,N14510,N14511);
and and8651(N14507,N14512,N14513);
and and8652(N14508,N14514,N14515);
and and8657(N14521,N14525,in1);
and and8658(N14522,N14526,N14527);
and and8659(N14523,N14528,N14529);
and and8660(N14524,N14530,N14531);
and and8665(N14537,N14541,N14542);
and and8666(N14538,N14543,N14544);
and and8667(N14539,N14545,R3);
and and8668(N14540,N14546,N14547);
and and8673(N14553,N14557,in0);
and and8674(N14554,N14558,N14559);
and and8675(N14555,N14560,N14561);
and and8676(N14556,N14562,N14563);
and and8681(N14568,N14572,N14573);
and and8682(N14569,in2,N14574);
and and8683(N14570,N14575,N14576);
and and8684(N14571,N14577,N14578);
and and8689(N14583,N14587,N14588);
and and8690(N14584,N14589,N14590);
and and8691(N14585,R1,N14591);
and and8692(N14586,N14592,N14593);
and and8697(N14598,N14602,N14603);
and and8698(N14599,N14604,R0);
and and8699(N14600,R1,N14605);
and and8700(N14601,N14606,N14607);
and and8705(N14613,N14617,N14618);
and and8706(N14614,N14619,N14620);
and and8707(N14615,N14621,N14622);
and and8708(N14616,R4,N14623);
and and8713(N14628,N14632,N14633);
and and8714(N14629,N14634,N14635);
and and8715(N14630,R1,N14636);
and and8716(N14631,N14637,R5);
and and8721(N14643,N14647,N14648);
and and8722(N14644,N14649,N14650);
and and8723(N14645,N14651,R3);
and and8724(N14646,N14652,R5);
and and8729(N14658,N14662,N14663);
and and8730(N14659,N14664,R0);
and and8731(N14660,N14665,N14666);
and and8732(N14661,N14667,R4);
and and8737(N14673,N14677,in0);
and and8738(N14674,N14678,N14679);
and and8739(N14675,N14680,N14681);
and and8740(N14676,R3,N14682);
and and8745(N14688,N14692,N14693);
and and8746(N14689,N14694,N14695);
and and8747(N14690,N14696,R1);
and and8748(N14691,N14697,R5);
and and8753(N14703,N14707,N14708);
and and8754(N14704,in2,N14709);
and and8755(N14705,N14710,N14711);
and and8756(N14706,R4,R5);
and and8761(N14717,N14721,in0);
and and8762(N14718,in1,N14722);
and and8763(N14719,N14723,N14724);
and and8764(N14720,N14725,N14726);
and and8769(N14731,N14735,N14736);
and and8770(N14732,N14737,N14738);
and and8771(N14733,R0,N14739);
and and8772(N14734,N14740,R3);
and and8777(N14745,N14749,N14750);
and and8778(N14746,in2,N14751);
and and8779(N14747,R2,N14752);
and and8780(N14748,N14753,N14754);
and and8785(N14759,N14763,in0);
and and8786(N14760,N14764,N14765);
and and8787(N14761,R2,N14766);
and and8788(N14762,N14767,N14768);
and and8793(N14773,N14777,N14778);
and and8794(N14774,in1,N14779);
and and8795(N14775,R2,R3);
and and8796(N14776,N14780,N14781);
and and8801(N14787,N14791,in0);
and and8802(N14788,N14792,N14793);
and and8803(N14789,N14794,N14795);
and and8804(N14790,R3,N14796);
and and8809(N14801,N14805,in0);
and and8810(N14802,in1,in2);
and and8811(N14803,N14806,N14807);
and and8812(N14804,N14808,N14809);
and and8817(N14815,N14819,in0);
and and8818(N14816,in1,N14820);
and and8819(N14817,N14821,N14822);
and and8820(N14818,N14823,N14824);
and and8825(N14829,N14833,N14834);
and and8826(N14830,in1,N14835);
and and8827(N14831,N14836,R1);
and and8828(N14832,N14837,N14838);
and and8833(N14843,N14847,N14848);
and and8834(N14844,N14849,in2);
and and8835(N14845,N14850,R1);
and and8836(N14846,N14851,N14852);
and and8841(N14857,N14861,in0);
and and8842(N14858,N14862,R0);
and and8843(N14859,N14863,R3);
and and8844(N14860,N14864,N14865);
and and8849(N14871,N14875,in0);
and and8850(N14872,N14876,R0);
and and8851(N14873,N14877,N14878);
and and8852(N14874,N14879,N14880);
and and8857(N14885,N14889,N14890);
and and8858(N14886,in1,R0);
and and8859(N14887,R1,N14891);
and and8860(N14888,N14892,N14893);
and and8865(N14899,N14903,in0);
and and8866(N14900,N14904,N14905);
and and8867(N14901,N14906,N14907);
and and8868(N14902,R4,N14908);
and and8873(N14913,N14917,in0);
and and8874(N14914,N14918,R0);
and and8875(N14915,R2,N14919);
and and8876(N14916,N14920,N14921);
and and8881(N14927,N14931,N14932);
and and8882(N14928,in1,N14933);
and and8883(N14929,N14934,R3);
and and8884(N14930,N14935,R5);
and and8889(N14941,N14945,N14946);
and and8890(N14942,N14947,in2);
and and8891(N14943,N14948,N14949);
and and8892(N14944,R3,N14950);
and and8897(N14955,N14959,N14960);
and and8898(N14956,in1,in2);
and and8899(N14957,N14961,N14962);
and and8900(N14958,R4,N14963);
and and8905(N14969,N14973,in0);
and and8906(N14970,N14974,N14975);
and and8907(N14971,R1,N14976);
and and8908(N14972,R4,N14977);
and and8913(N14983,N14987,in0);
and and8914(N14984,N14988,R0);
and and8915(N14985,N14989,N14990);
and and8916(N14986,N14991,N14992);
and and8921(N14997,N15001,N15002);
and and8922(N14998,N15003,N15004);
and and8923(N14999,R1,R2);
and and8924(N15000,N15005,N15006);
and and8929(N15011,N15015,in0);
and and8930(N15012,in1,N15016);
and and8931(N15013,N15017,N15018);
and and8932(N15014,R3,N15019);
and and8937(N15025,N15029,in0);
and and8938(N15026,N15030,N15031);
and and8939(N15027,N15032,R1);
and and8940(N15028,N15033,N15034);
and and8945(N15039,N15043,N15044);
and and8946(N15040,in1,N15045);
and and8947(N15041,N15046,R1);
and and8948(N15042,N15047,N15048);
and and8953(N15053,N15057,N15058);
and and8954(N15054,in1,in2);
and and8955(N15055,R0,N15059);
and and8956(N15056,N15060,N15061);
and and8961(N15067,N15071,N15072);
and and8962(N15068,N15073,N15074);
and and8963(N15069,N15075,R2);
and and8964(N15070,R4,N15076);
and and8969(N15081,N15085,in1);
and and8970(N15082,N15086,N15087);
and and8971(N15083,R2,R3);
and and8972(N15084,N15088,N15089);
and and8977(N15095,N15099,in0);
and and8978(N15096,N15100,R0);
and and8979(N15097,N15101,N15102);
and and8980(N15098,N15103,N15104);
and and8985(N15109,N15113,N15114);
and and8986(N15110,in2,N15115);
and and8987(N15111,N15116,N15117);
and and8988(N15112,R4,N15118);
and and8993(N15123,N15127,in0);
and and8994(N15124,N15128,N15129);
and and8995(N15125,N15130,R2);
and and8996(N15126,R4,N15131);
and and9001(N15137,N15141,N15142);
and and9002(N15138,in1,N15143);
and and9003(N15139,N15144,R1);
and and9004(N15140,N15145,N15146);
and and9009(N15151,N15155,N15156);
and and9010(N15152,in1,N15157);
and and9011(N15153,R1,N15158);
and and9012(N15154,N15159,R5);
and and9017(N15165,N15169,N15170);
and and9018(N15166,in1,in2);
and and9019(N15167,N15171,N15172);
and and9020(N15168,R4,N15173);
and and9025(N15179,N15183,in0);
and and9026(N15180,in2,R0);
and and9027(N15181,N15184,N15185);
and and9028(N15182,N15186,N15187);
and and9033(N15193,N15197,N15198);
and and9034(N15194,in1,N15199);
and and9035(N15195,R1,R3);
and and9036(N15196,R4,N15200);
and and9041(N15206,N15210,in0);
and and9042(N15207,in1,N15211);
and and9043(N15208,N15212,R3);
and and9044(N15209,R4,N15213);
and and9049(N15219,N15223,N15224);
and and9050(N15220,R0,N15225);
and and9051(N15221,R2,R3);
and and9052(N15222,N15226,N15227);
and and9057(N15232,N15236,in0);
and and9058(N15233,in1,N15237);
and and9059(N15234,N15238,R2);
and and9060(N15235,R4,N15239);
and and9065(N15245,N15249,N15250);
and and9066(N15246,N15251,N15252);
and and9067(N15247,R1,N15253);
and and9068(N15248,R4,N15254);
and and9073(N15258,N15262,in1);
and and9074(N15259,in2,N15263);
and and9075(N15260,R1,R2);
and and9076(N15261,N15264,N15265);
and and9081(N15271,N15275,in0);
and and9082(N15272,in1,N15276);
and and9083(N15273,N15277,R1);
and and9084(N15274,R2,N15278);
and and9089(N15284,N15288,N15289);
and and9090(N15285,N15290,in2);
and and9091(N15286,N15291,R2);
and and9092(N15287,R4,R5);
and and9097(N15297,N15301,N15302);
and and9098(N15298,in1,in2);
and and9099(N15299,N15303,N15304);
and and9100(N15300,R3,N15305);
and and9105(N15310,N15314,in0);
and and9106(N15311,N15315,N15316);
and and9107(N15312,R2,R3);
and and9108(N15313,N15317,N15318);
and and9113(N15323,N15327,N15328);
and and9114(N15324,in1,N15329);
and and9115(N15325,R0,R1);
and and9116(N15326,R4,N15330);
and and9121(N15336,N15340,in0);
and and9122(N15337,in2,N15341);
and and9123(N15338,R1,N15342);
and and9124(N15339,N15343,N15344);
and and9129(N15349,N15353,in0);
and and9130(N15350,in1,N15354);
and and9131(N15351,N15355,R1);
and and9132(N15352,N15356,N15357);
and and9137(N15362,N15366,in0);
and and9138(N15363,in1,N15367);
and and9139(N15364,R0,N15368);
and and9140(N15365,R3,N15369);
and and9145(N15375,N15379,N15380);
and and9146(N15376,N15381,N15382);
and and9147(N15377,R1,N15383);
and and9148(N15378,R4,R5);
and and9153(N15388,N15392,in0);
and and9154(N15389,N15393,N15394);
and and9155(N15390,N15395,R3);
and and9156(N15391,N15396,R5);
and and9161(N15401,N15405,in0);
and and9162(N15402,N15406,N15407);
and and9163(N15403,N15408,R3);
and and9164(N15404,R4,N15409);
and and9169(N15414,N15418,in0);
and and9170(N15415,in1,N15419);
and and9171(N15416,R0,R2);
and and9172(N15417,N15420,N15421);
and and9177(N15427,N15431,N15432);
and and9178(N15428,in2,R0);
and and9179(N15429,R2,N15433);
and and9180(N15430,R4,N15434);
and and9185(N15440,N15444,N15445);
and and9186(N15441,in2,R1);
and and9187(N15442,N15446,N15447);
and and9188(N15443,N15448,R5);
and and9193(N15453,N15457,in0);
and and9194(N15454,N15458,N15459);
and and9195(N15455,R1,N15460);
and and9196(N15456,N15461,R5);
and and9201(N15466,N15470,in0);
and and9202(N15467,in1,N15471);
and and9203(N15468,N15472,N15473);
and and9204(N15469,R3,N15474);
and and9209(N15479,N15483,N15484);
and and9210(N15480,N15485,R0);
and and9211(N15481,R2,R3);
and and9212(N15482,N15486,R5);
and and9217(N15492,N15496,in0);
and and9218(N15493,in1,R1);
and and9219(N15494,N15497,N15498);
and and9220(N15495,R4,N15499);
and and9225(N15505,N15509,in1);
and and9226(N15506,N15510,N15511);
and and9227(N15507,N15512,R3);
and and9228(N15508,N15513,R5);
and and9233(N15518,N15522,N15523);
and and9234(N15519,in1,N15524);
and and9235(N15520,R1,N15525);
and and9236(N15521,R4,N15526);
and and9241(N15531,N15535,N15536);
and and9242(N15532,N15537,R0);
and and9243(N15533,R1,N15538);
and and9244(N15534,N15539,N15540);
and and9249(N15544,N15548,in0);
and and9250(N15545,N15549,N15550);
and and9251(N15546,R1,N15551);
and and9252(N15547,N15552,R4);
and and9257(N15557,N15561,N15562);
and and9258(N15558,in1,in2);
and and9259(N15559,R0,N15563);
and and9260(N15560,R4,N15564);
and and9265(N15570,N15574,in0);
and and9266(N15571,N15575,in2);
and and9267(N15572,R0,N15576);
and and9268(N15573,N15577,R4);
and and9273(N15583,N15587,in0);
and and9274(N15584,N15588,N15589);
and and9275(N15585,N15590,R2);
and and9276(N15586,R3,N15591);
and and9281(N15596,N15600,N15601);
and and9282(N15597,in2,R0);
and and9283(N15598,N15602,R2);
and and9284(N15599,N15603,N15604);
and and9289(N15609,N15613,N15614);
and and9290(N15610,in2,R0);
and and9291(N15611,R1,N15615);
and and9292(N15612,N15616,N15617);
and and9297(N15622,N15626,N15627);
and and9298(N15623,N15628,N15629);
and and9299(N15624,R0,R1);
and and9300(N15625,R2,N15630);
and and9305(N15635,N15639,N15640);
and and9306(N15636,N15641,R0);
and and9307(N15637,R1,N15642);
and and9308(N15638,R4,R5);
and and9313(N15648,N15652,in0);
and and9314(N15649,N15653,N15654);
and and9315(N15650,N15655,R2);
and and9316(N15651,N15656,R4);
and and9321(N15661,N15665,N15666);
and and9322(N15662,N15667,N15668);
and and9323(N15663,R1,N15669);
and and9324(N15664,R4,N15670);
and and9329(N15674,N15678,N15679);
and and9330(N15675,N15680,in2);
and and9331(N15676,R1,R2);
and and9332(N15677,N15681,N15682);
and and9337(N15687,N15691,in0);
and and9338(N15688,in1,N15692);
and and9339(N15689,N15693,N15694);
and and9340(N15690,R3,R4);
and and9345(N15700,N15704,in0);
and and9346(N15701,in2,R0);
and and9347(N15702,N15705,N15706);
and and9348(N15703,N15707,N15708);
and and9353(N15713,N15717,in0);
and and9354(N15714,N15718,in2);
and and9355(N15715,N15719,R2);
and and9356(N15716,N15720,N15721);
and and9361(N15726,N15730,N15731);
and and9362(N15727,N15732,in2);
and and9363(N15728,R0,R2);
and and9364(N15729,N15733,R4);
and and9369(N15739,N15743,in0);
and and9370(N15740,N15744,N15745);
and and9371(N15741,R1,R2);
and and9372(N15742,N15746,N15747);
and and9377(N15752,N15756,N15757);
and and9378(N15753,in1,N15758);
and and9379(N15754,R1,R2);
and and9380(N15755,N15759,N15760);
and and9385(N15765,N15769,in0);
and and9386(N15766,N15770,N15771);
and and9387(N15767,R1,R2);
and and9388(N15768,N15772,R4);
and and9393(N15778,N15782,N15783);
and and9394(N15779,N15784,R0);
and and9395(N15780,R1,N15785);
and and9396(N15781,R4,R5);
and and9401(N15791,N15795,N15796);
and and9402(N15792,N15797,N15798);
and and9403(N15793,R0,N15799);
and and9404(N15794,R3,N15800);
and and9409(N15804,N15808,in0);
and and9410(N15805,N15809,N15810);
and and9411(N15806,N15811,N15812);
and and9412(N15807,R2,R3);
and and9417(N15817,N15821,N15822);
and and9418(N15818,in2,N15823);
and and9419(N15819,R1,N15824);
and and9420(N15820,R3,N15825);
and and9425(N15829,N15833,in0);
and and9426(N15830,in1,in2);
and and9427(N15831,N15834,N15835);
and and9428(N15832,R4,R5);
and and9433(N15841,N15845,in1);
and and9434(N15842,in2,R0);
and and9435(N15843,N15846,R2);
and and9436(N15844,N15847,N15848);
and and9441(N15853,N15857,in0);
and and9442(N15854,R0,R1);
and and9443(N15855,N15858,N15859);
and and9444(N15856,R4,N15860);
and and9449(N15865,N15869,in0);
and and9450(N15866,N15870,R0);
and and9451(N15867,N15871,R2);
and and9452(N15868,N15872,R4);
and and9457(N15877,N15881,in2);
and and9458(N15878,N15882,R1);
and and9459(N15879,N15883,R3);
and and9460(N15880,N15884,R5);
and and9465(N15889,N15893,in1);
and and9466(N15890,in2,N15894);
and and9467(N15891,R1,N15895);
and and9468(N15892,N15896,N15897);
and and9473(N15901,N15905,in0);
and and9474(N15902,in2,N15906);
and and9475(N15903,R1,N15907);
and and9476(N15904,N15908,N15909);
and and9481(N15913,N15917,in0);
and and9482(N15914,N15918,R0);
and and9483(N15915,R1,N15919);
and and9484(N15916,N15920,R5);
and and9489(N15925,N15929,in1);
and and9490(N15926,N15930,R0);
and and9491(N15927,R1,R2);
and and9492(N15928,N15931,N15932);
and and9497(N15937,N15941,in0);
and and9498(N15938,N15942,R0);
and and9499(N15939,R1,R2);
and and9500(N15940,N15943,N15944);
and and9505(N15949,N15953,in0);
and and9506(N15950,in1,in2);
and and9507(N15951,R0,R3);
and and9508(N15952,N15954,N15955);
and and9513(N15961,N15965,N15966);
and and9514(N15962,N15967,R0);
and and9515(N15963,R1,R2);
and and9516(N15964,R3,N15968);
and and9521(N15973,N15977,N15978);
and and9522(N15974,in1,N15979);
and and9523(N15975,R2,R3);
and and9524(N15976,N15980,R5);
and and9529(N15985,N15989,in0);
and and9530(N15986,N15990,R0);
and and9531(N15987,R2,N15991);
and and9532(N15988,N15992,N15993);
and and9537(N15997,N16001,in2);
and and9538(N15998,R0,N16002);
and and9539(N15999,R2,N16003);
and and9540(N16000,N16004,N16005);
and and9545(N16009,N16013,in0);
and and9546(N16010,N16014,N16015);
and and9547(N16011,R1,R3);
and and9548(N16012,N16016,R5);
and and9553(N16021,N16025,in1);
and and9554(N16022,N16026,N16027);
and and9555(N16023,R1,N16028);
and and9556(N16024,R3,N16029);
and and9561(N16033,N16037,in0);
and and9562(N16034,in1,N16038);
and and9563(N16035,R2,N16039);
and and9564(N16036,N16040,R5);
and and9569(N16045,N16049,N16050);
and and9570(N16046,in1,in2);
and and9571(N16047,N16051,R2);
and and9572(N16048,N16052,R5);
and and9577(N16057,N16061,N16062);
and and9578(N16058,N16063,R1);
and and9579(N16059,N16064,R3);
and and9580(N16060,N16065,R5);
and and9585(N16069,N16073,in0);
and and9586(N16070,in1,in2);
and and9587(N16071,R0,N16074);
and and9588(N16072,R2,N16075);
and and9593(N16081,N16085,in0);
and and9594(N16082,in1,in2);
and and9595(N16083,N16086,R1);
and and9596(N16084,N16087,R5);
and and9601(N16093,N16097,N16098);
and and9602(N16094,in1,N16099);
and and9603(N16095,R0,R2);
and and9604(N16096,R3,N16100);
and and9609(N16105,N16109,N16110);
and and9610(N16106,N16111,in2);
and and9611(N16107,R0,R1);
and and9612(N16108,N16112,R4);
and and9617(N16117,N16121,N16122);
and and9618(N16118,in1,N16123);
and and9619(N16119,R1,N16124);
and and9620(N16120,R3,R4);
and and9625(N16129,N16133,N16134);
and and9626(N16130,R0,N16135);
and and9627(N16131,R2,N16136);
and and9628(N16132,R4,N16137);
and and9633(N16141,N16145,in2);
and and9634(N16142,N16146,N16147);
and and9635(N16143,R2,N16148);
and and9636(N16144,R4,N16149);
and and9641(N16153,N16157,in1);
and and9642(N16154,N16158,N16159);
and and9643(N16155,R2,N16160);
and and9644(N16156,R4,N16161);
and and9649(N16165,N16169,in1);
and and9650(N16166,in2,N16170);
and and9651(N16167,R1,R2);
and and9652(N16168,N16171,N16172);
and and9657(N16177,N16181,in0);
and and9658(N16178,N16182,in2);
and and9659(N16179,N16183,R1);
and and9660(N16180,R2,N16184);
and and9665(N16189,N16193,N16194);
and and9666(N16190,N16195,N16196);
and and9667(N16191,R1,R3);
and and9668(N16192,R4,R5);
and and9673(N16201,N16205,in0);
and and9674(N16202,in1,in2);
and and9675(N16203,R0,N16206);
and and9676(N16204,N16207,R4);
and and9681(N16213,N16217,N16218);
and and9682(N16214,N16219,N16220);
and and9683(N16215,R1,N16221);
and and9684(N16216,R3,R4);
and and9689(N16225,N16229,N16230);
and and9690(N16226,in2,R0);
and and9691(N16227,R1,N16231);
and and9692(N16228,R3,R5);
and and9697(N16237,N16241,in2);
and and9698(N16238,R0,R1);
and and9699(N16239,R2,N16242);
and and9700(N16240,N16243,N16244);
and and9705(N16249,N16253,N16254);
and and9706(N16250,in1,R0);
and and9707(N16251,N16255,R2);
and and9708(N16252,N16256,R4);
and and9713(N16261,N16265,in1);
and and9714(N16262,N16266,R0);
and and9715(N16263,N16267,R3);
and and9716(N16264,R4,R5);
and and9721(N16273,N16277,in0);
and and9722(N16274,in2,N16278);
and and9723(N16275,N16279,R2);
and and9724(N16276,N16280,R4);
and and9729(N16285,N16289,N16290);
and and9730(N16286,in1,in2);
and and9731(N16287,N16291,R3);
and and9732(N16288,N16292,R5);
and and9737(N16297,N16301,in0);
and and9738(N16298,N16302,R0);
and and9739(N16299,R1,N16303);
and and9740(N16300,N16304,R5);
and and9745(N16309,N16313,in0);
and and9746(N16310,N16314,R0);
and and9747(N16311,N16315,R3);
and and9748(N16312,N16316,N16317);
and and9753(N16321,N16325,in1);
and and9754(N16322,in2,R1);
and and9755(N16323,N16326,N16327);
and and9756(N16324,N16328,R5);
and and9761(N16333,N16337,N16338);
and and9762(N16334,in1,N16339);
and and9763(N16335,R0,R1);
and and9764(N16336,R3,R4);
and and9769(N16345,N16349,in0);
and and9770(N16346,in1,in2);
and and9771(N16347,N16350,R1);
and and9772(N16348,N16351,N16352);
and and9777(N16357,N16361,in0);
and and9778(N16358,N16362,R0);
and and9779(N16359,R1,N16363);
and and9780(N16360,N16364,N16365);
and and9785(N16369,N16373,in0);
and and9786(N16370,in1,in2);
and and9787(N16371,R1,N16374);
and and9788(N16372,N16375,N16376);
and and9793(N16381,N16385,in0);
and and9794(N16382,N16386,in2);
and and9795(N16383,R0,N16387);
and and9796(N16384,R2,N16388);
and and9801(N16393,N16397,in0);
and and9802(N16394,in1,N16398);
and and9803(N16395,R0,N16399);
and and9804(N16396,R2,N16400);
and and9809(N16405,N16409,N16410);
and and9810(N16406,in1,R0);
and and9811(N16407,N16411,R3);
and and9812(N16408,R4,R5);
and and9817(N16417,N16421,in0);
and and9818(N16418,N16422,R0);
and and9819(N16419,R1,R2);
and and9820(N16420,N16423,R5);
and and9825(N16429,N16433,in0);
and and9826(N16430,N16434,R0);
and and9827(N16431,R1,N16435);
and and9828(N16432,R4,R5);
and and9833(N16441,N16445,in0);
and and9834(N16442,N16446,N16447);
and and9835(N16443,N16448,R1);
and and9836(N16444,R2,R3);
and and9841(N16453,N16457,in0);
and and9842(N16454,in1,N16458);
and and9843(N16455,R1,N16459);
and and9844(N16456,R3,N16460);
and and9849(N16464,N16468,in0);
and and9850(N16465,in1,N16469);
and and9851(N16466,R0,R1);
and and9852(N16467,R2,R3);
and and9857(N16475,N16479,N16480);
and and9858(N16476,in1,in2);
and and9859(N16477,R0,R1);
and and9860(N16478,R2,R3);
and and9865(N16486,N16490,in1);
and and9866(N16487,in2,N16491);
and and9867(N16488,R1,N16492);
and and9868(N16489,R3,R4);
and and9873(N16497,N16501,N16502);
and and9874(N16498,R0,R1);
and and9875(N16499,R2,R3);
and and9876(N16500,N16503,R5);
and and9881(N16508,N16512,in0);
and and9882(N16509,N16513,N16514);
and and9883(N16510,R1,R3);
and and9884(N16511,R4,N16515);
and and9889(N16519,N16523,in1);
and and9890(N16520,in2,R0);
and and9891(N16521,R1,N16524);
and and9892(N16522,R3,N16525);
and and9897(N16530,N16534,in0);
and and9898(N16531,in1,N16535);
and and9899(N16532,R0,R1);
and and9900(N16533,N16536,R3);
and and9905(N16541,N16545,in0);
and and9906(N16542,N16546,R0);
and and9907(N16543,N16547,R2);
and and9908(N16544,R3,R5);
and and9913(N16552,N16556,in1);
and and9914(N16553,R0,N16557);
and and9915(N16554,N16558,R3);
and and9916(N16555,R4,R5);
and and9921(N16563,N16567,in0);
and and9922(N16564,R0,N16568);
and and9923(N16565,N16569,R3);
and and9924(N16566,R4,R5);
and and9929(N16574,N16578,N16579);
and and9930(N16575,in2,R0);
and and9931(N16576,N16580,R3);
and and9932(N16577,R4,N16581);
and and9937(N16585,N16589,in0);
and and9938(N16586,N16590,in2);
and and9939(N16587,N16591,R2);
and and9940(N16588,R3,R5);
and and9945(N16596,N16600,in0);
and and9946(N16597,in1,N16601);
and and9947(N16598,N16602,R2);
and and9948(N16599,R3,R5);
and and9953(N16607,N16611,in0);
and and9954(N16608,in1,in2);
and and9955(N16609,N16612,R1);
and and9956(N16610,R2,N16613);
and and9961(N16618,N16622,in0);
and and9962(N16619,N16623,N16624);
and and9963(N16620,R1,R2);
and and9964(N16621,R3,R4);
and and9969(N16629,N16633,N16634);
and and9970(N16630,N16635,N16636);
and and9971(N16631,R2,R3);
and and9972(N16632,R4,R5);
and and9977(N16640,N16644,in0);
and and9978(N16641,in1,in2);
and and9979(N16642,N16645,R3);
and and9980(N16643,N16646,R5);
and and9985(N16651,N16655,in0);
and and9986(N16652,in1,in2);
and and9987(N16653,N16656,R3);
and and9988(N16654,N16657,N16658);
and and9993(N16662,N16666,in0);
and and9994(N16663,N16667,in2);
and and9995(N16664,N16668,R2);
and and9996(N16665,R3,R4);
and and10001(N16673,N16677,in0);
and and10002(N16674,N16678,R0);
and and10003(N16675,R1,R2);
and and10004(N16676,N16679,R4);
and and10009(N16684,N16688,in0);
and and10010(N16685,N16689,N16690);
and and10011(N16686,R1,R2);
and and10012(N16687,R3,R4);
and and10017(N16695,N16699,in0);
and and10018(N16696,in2,R0);
and and10019(N16697,R1,N16700);
and and10020(N16698,N16701,N16702);
and and10025(N16706,N16710,in0);
and and10026(N16707,N16711,N16712);
and and10027(N16708,R1,N16713);
and and10028(N16709,R3,R4);
and and10033(N16717,N16721,in1);
and and10034(N16718,N16722,R1);
and and10035(N16719,N16723,R3);
and and10036(N16720,R4,R5);
and and10041(N16728,N16732,in0);
and and10042(N16729,N16733,N16734);
and and10043(N16730,R1,R2);
and and10044(N16731,N16735,R4);
and and10049(N16739,N16743,in0);
and and10050(N16740,in2,R0);
and and10051(N16741,R1,N16744);
and and10052(N16742,R3,N16745);
and and10057(N16750,N16754,N16755);
and and10058(N16751,R0,N16756);
and and10059(N16752,R2,R3);
and and10060(N16753,R4,R5);
and and10065(N16761,N16765,N16766);
and and10066(N16762,in1,R0);
and and10067(N16763,R1,N16767);
and and10068(N16764,R3,N16768);
and and10073(N16772,N16776,N16777);
and and10074(N16773,in1,N16778);
and and10075(N16774,R1,R2);
and and10076(N16775,R3,R5);
and and10081(N16783,N16787,in0);
and and10082(N16784,in2,R0);
and and10083(N16785,N16788,R3);
and and10084(N16786,R4,N16789);
and and10089(N16794,N16798,in0);
and and10090(N16795,in2,R0);
and and10091(N16796,R1,R2);
and and10092(N16797,N16799,N16800);
and and10097(N16805,N16809,in1);
and and10098(N16806,in2,N16810);
and and10099(N16807,R1,N16811);
and and10100(N16808,R3,N16812);
and and10105(N16816,N16820,in0);
and and10106(N16817,in1,N16821);
and and10107(N16818,R0,R1);
and and10108(N16819,R2,N16822);
and and10113(N16827,N16831,in0);
and and10114(N16828,in1,R0);
and and10115(N16829,R1,N16832);
and and10116(N16830,N16833,R4);
and and10121(N16838,N16842,in0);
and and10122(N16839,R0,N16843);
and and10123(N16840,R2,N16844);
and and10124(N16841,R4,N16845);
and and10129(N16849,N16853,in0);
and and10130(N16850,N16854,R0);
and and10131(N16851,N16855,R2);
and and10132(N16852,R4,N16856);
and and10137(N16860,N16864,in0);
and and10138(N16861,N16865,in2);
and and10139(N16862,R0,R1);
and and10140(N16863,R2,R5);
and and10145(N16871,N16875,in0);
and and10146(N16872,in1,N16876);
and and10147(N16873,R0,R3);
and and10148(N16874,R4,R5);
and and10153(N16882,N16886,in0);
and and10154(N16883,N16887,R0);
and and10155(N16884,R2,N16888);
and and10156(N16885,R4,N16889);
and and10161(N16893,N16897,in0);
and and10162(N16894,in2,R0);
and and10163(N16895,R1,R2);
and and10164(N16896,R3,N16898);
and and10169(N16903,N16907,N16908);
and and10170(N16904,in2,N16909);
and and10171(N16905,R2,R3);
and and10172(N16906,R4,R5);
and and10177(N16913,N16917,N16918);
and and10178(N16914,N16919,R0);
and and10179(N16915,R1,R2);
and and10180(N16916,R3,R5);
and and10185(N16923,N16927,in0);
and and10186(N16924,in1,in2);
and and10187(N16925,R0,R2);
and and10188(N16926,R3,N16928);
and and10193(N16933,N16937,N16938);
and and10194(N16934,N16939,in2);
and and10195(N16935,R0,R1);
and and10196(N16936,R3,R5);
and and10201(N16943,N16947,N16948);
and and10202(N16944,N16949,R1);
and and10203(N16945,R2,R3);
and and10204(N16946,R4,R5);
and and10209(N16953,N16957,in0);
and and10210(N16954,N16958,in2);
and and10211(N16955,R1,R3);
and and10212(N16956,R4,R5);
and and10217(N16963,N16967,in0);
and and10218(N16964,in1,in2);
and and10219(N16965,R0,R2);
and and10220(N16966,R3,N16968);
and and10225(N16973,N16977,in0);
and and10226(N16974,in1,N16978);
and and10227(N16975,R1,R2);
and and10228(N16976,R4,R5);
and and10233(N16983,N16987,in0);
and and10234(N16984,in1,in2);
and and10235(N16985,R0,R2);
and and10236(N16986,N16988,R4);
and and10241(N16993,N16997,in0);
and and10242(N16994,in1,in2);
and and10243(N16995,R0,R1);
and and10244(N16996,R2,N16998);
and and10249(N17003,N17007,in0);
and and10250(N17004,in1,N17008);
and and10251(N17005,R1,R2);
and and10252(N17006,R3,N17009);
and and10257(N17013,N17017,in1);
and and10258(N17014,R0,R1);
and and10259(N17015,R2,N17018);
and and10260(N17016,R4,N17019);
and and10265(N17023,N17027,in0);
and and10266(N17024,in1,in2);
and and10267(N17025,N17028,R1);
and and10268(N17026,R2,N17029);
and and10273(N17033,N17037,in0);
and and10274(N17034,in1,N17038);
and and10275(N17035,R0,R1);
and and10276(N17036,R2,R3);
and and10281(N17043,N17047,in0);
and and10282(N17044,N17048,in2);
and and10283(N17045,R1,R2);
and and10284(N17046,R3,N17049);
and and10289(N17053,N17057,in0);
and and10290(N17054,in1,in2);
and and10291(N17055,R1,N17058);
and and10292(N17056,R4,R5);
and and10297(N17063,N17067,in0);
and and10298(N17064,in1,R0);
and and10299(N17065,R1,N17068);
and and10300(N17066,R3,R4);
and and10305(N17072,N17076,in1);
and and10306(N17073,R0,R1);
and and10307(N17074,N17077,R3);
and and10308(N17075,R4,R5);
and and10313(N17081,N17085,in0);
and and10314(N17082,R0,R1);
and and10315(N17083,N17086,R3);
and and10316(N17084,R4,R5);
and and10321(N17090,N17094,in0);
and and10322(N17091,in2,R0);
and and10323(N17092,N17095,R2);
and and10324(N17093,R3,R5);
and and10329(N17099,N17103,in0);
and and10330(N17100,in1,R0);
and and10331(N17101,N17104,R2);
and and10332(N17102,R3,R5);
and and10337(N17108,N17112,in0);
and and10338(N17109,N17113,R0);
and and10339(N17110,R1,R2);
and and10340(N17111,R3,R4);
and and10345(N17117,N17121,in0);
and and10346(N17118,in1,in2);
and and10347(N17119,R1,N17122);
and and10348(N17120,R3,R4);
and and10353(N17126,N17130,in0);
and and10354(N17127,in1,in2);
and and10355(N17128,R0,R1);
and and10356(N17129,R3,N17131);
and and10361(N17135,N17139,in0);
and and10362(N17136,in1,in2);
and and10363(N17137,N17140,R1);
and and10364(N17138,R2,R3);
and and10369(N17144,N17148,in0);
and and10370(N17145,in1,N17149);
and and10371(N17146,R1,R2);
and and10372(N17147,R3,R4);
and and10377(N17153,N17157,in0);
and and10378(N17154,in1,R0);
and and10379(N17155,R1,R2);
and and10380(N17156,R3,R4);
and and10385(N17161,N17165,N17166);
and and10386(N17162,N17167,N17168);
and and10387(N17163,N17169,R4);
and and10388(N17164,N17170,N17171);
and and10392(N17175,N17179,N17180);
and and10393(N17176,N17181,R2);
and and10394(N17177,N17182,N17183);
and and10395(N17178,N17184,N17185);
and and10399(N17189,N17193,R0);
and and10400(N17190,N17194,N17195);
and and10401(N17191,N17196,N17197);
and and10402(N17192,N17198,N17199);
and and10406(N17203,N17207,R0);
and and10407(N17204,N17208,N17209);
and and10408(N17205,N17210,N17211);
and and10409(N17206,N17212,N17213);
and and10413(N17217,N17221,N17222);
and and10414(N17218,N17223,R2);
and and10415(N17219,R4,N17224);
and and10416(N17220,N17225,N17226);
and and10420(N17230,N17234,N17235);
and and10421(N17231,R1,R2);
and and10422(N17232,N17236,N17237);
and and10423(N17233,N17238,N17239);
and and10427(N17243,N17247,N17248);
and and10428(N17244,R2,R3);
and and10429(N17245,N17249,N17250);
and and10430(N17246,N17251,N17252);
and and10434(N17256,in2,N17260);
and and10435(N17257,N17261,R3);
and and10436(N17258,N17262,N17263);
and and10437(N17259,N17264,N17265);
and and10441(N17269,in0,N17273);
and and10442(N17270,N17274,R2);
and and10443(N17271,N17275,N17276);
and and10444(N17272,N17277,N17278);
and and10448(N17282,in0,R0);
and and10449(N17283,R1,N17286);
and and10450(N17284,N17287,N17288);
and and10451(N17285,N17289,N17290);
and and10455(N17294,N17298,N17299);
and and10456(N17295,R2,N17300);
and and10457(N17296,N17301,R5);
and and10458(N17297,N17302,R7);
and and10462(N17306,in0,N17310);
and and10463(N17307,N17311,R2);
and and10464(N17308,N17312,N17313);
and and10465(N17309,R6,N17314);
and and10469(N17318,in0,N17322);
and and10470(N17319,N17323,R1);
and and10471(N17320,N17324,R5);
and and10472(N17321,N17325,N17326);
and and10476(N17330,in0,N17334);
and and10477(N17331,in2,N17335);
and and10478(N17332,R4,N17336);
and and10479(N17333,N17337,N17338);
and and10483(N17342,N17346,N17347);
and and10484(N17343,R1,N17348);
and and10485(N17344,N17349,R4);
and and10486(N17345,N17350,R7);
and and10490(N17354,in2,N17358);
and and10491(N17355,R1,N17359);
and and10492(N17356,N17360,N17361);
and and10493(N17357,N17362,R7);
and and10497(N17366,N17370,R0);
and and10498(N17367,R1,N17371);
and and10499(N17368,N17372,N17373);
and and10500(N17369,R6,N17374);
and and10504(N17378,in0,N17382);
and and10505(N17379,N17383,R1);
and and10506(N17380,N17384,R5);
and and10507(N17381,N17385,N17386);
and and10511(N17390,N17394,R0);
and and10512(N17391,R1,R2);
and and10513(N17392,R3,N17395);
and and10514(N17393,N17396,N17397);
and and10518(N17401,in0,N17405);
and and10519(N17402,R2,N17406);
and and10520(N17403,R4,R5);
and and10521(N17404,N17407,N17408);
and and10525(N17412,in0,R0);
and and10526(N17413,R1,N17416);
and and10527(N17414,N17417,N17418);
and and10528(N17415,R5,N17419);
and and10532(N17423,N17427,N17428);
and and10533(N17424,R1,R2);
and and10534(N17425,N17429,R5);
and and10535(N17426,R6,N17430);
and and10539(N17434,in0,N17438);
and and10540(N17435,N17439,R3);
and and10541(N17436,N17440,N17441);
and and10542(N17437,R6,R7);
and and10546(N17445,in0,in2);
and and10547(N17446,N17449,N17450);
and and10548(N17447,R3,N17451);
and and10549(N17448,R5,N17452);
and and10553(N17456,N17460,N17461);
and and10554(N17457,N17462,R3);
and and10555(N17458,R4,N17463);
and and10556(N17459,R6,R7);
and and10560(N17467,in0,N17471);
and and10561(N17468,N17472,R1);
and and10562(N17469,R4,N17473);
and and10563(N17470,N17474,R7);
and and10567(N17478,in0,N17482);
and and10568(N17479,N17483,R1);
and and10569(N17480,R2,N17484);
and and10570(N17481,N17485,R6);
and and10574(N17489,N17493,R0);
and and10575(N17490,R1,N17494);
and and10576(N17491,R3,N17495);
and and10577(N17492,R5,N17496);
and and10581(N17500,in0,N17504);
and and10582(N17501,R0,N17505);
and and10583(N17502,R2,N17506);
and and10584(N17503,R5,N17507);
and and10588(N17511,N17515,N17516);
and and10589(N17512,R0,N17517);
and and10590(N17513,R3,R4);
and and10591(N17514,R5,N17518);
and and10595(N17522,in0,N17526);
and and10596(N17523,R1,R2);
and and10597(N17524,N17527,R5);
and and10598(N17525,N17528,N17529);
and and10602(N17533,in0,N17537);
and and10603(N17534,in2,R1);
and and10604(N17535,N17538,N17539);
and and10605(N17536,R5,N17540);
and and10609(N17544,in0,in1);
and and10610(N17545,N17548,N17549);
and and10611(N17546,R1,R2);
and and10612(N17547,N17550,N17551);
and and10616(N17555,in0,N17559);
and and10617(N17556,N17560,R1);
and and10618(N17557,R4,N17561);
and and10619(N17558,N17562,R7);
and and10623(N17566,in0,N17570);
and and10624(N17567,R0,N17571);
and and10625(N17568,R2,N17572);
and and10626(N17569,R5,N17573);
and and10630(N17577,in0,N17581);
and and10631(N17578,R0,R1);
and and10632(N17579,N17582,R3);
and and10633(N17580,N17583,R7);
and and10637(N17587,N17591,in2);
and and10638(N17588,R1,R2);
and and10639(N17589,R3,N17592);
and and10640(N17590,R6,N17593);
and and10644(N17597,in0,N17601);
and and10645(N17598,R0,R1);
and and10646(N17599,N17602,R4);
and and10647(N17600,R6,N17603);
and and10651(N17607,in0,R1);
and and10652(N17608,N17611,N17612);
and and10653(N17609,R4,R5);
and and10654(N17610,N17613,R7);
and and10658(N17617,in0,N17621);
and and10659(N17618,R0,N17622);
and and10660(N17619,R3,R4);
and and10661(N17620,N17623,R7);
and and10665(N17627,in2,N17631);
and and10666(N17628,N17632,R3);
and and10667(N17629,R4,N17633);
and and10668(N17630,R6,R7);
and and10672(N17637,in0,N17641);
and and10673(N17638,R0,N17642);
and and10674(N17639,R3,R4);
and and10675(N17640,R5,N17643);
and and6907(N11889,N11896,N11897);
and and6908(N11890,N11898,N11899);
and and6916(N11907,N11915,N11916);
and and6917(N11908,R6,N11917);
and and6925(N11925,N11932,N11933);
and and6926(N11926,N11934,R7);
and and6934(N11942,N11949,N11950);
and and6935(N11943,N11951,R7);
and and6943(N11959,R3,N11966);
and and6944(N11960,N11967,N11968);
and and6952(N11976,N11983,N11984);
and and6953(N11977,N11985,R7);
and and6961(N11993,N11998,N11999);
and and6962(N11994,N12000,N12001);
and and6970(N12009,R4,N12016);
and and6971(N12010,N12017,R7);
and and6979(N12025,N12031,N12032);
and and6980(N12026,R6,N12033);
and and6988(N12041,R3,N12048);
and and6989(N12042,N12049,R7);
and and6997(N12057,N12064,R5);
and and6998(N12058,N12065,R7);
and and7006(N12073,N12080,N12081);
and and7007(N12074,R6,R7);
and and7015(N12089,R4,N12096);
and and7016(N12090,R6,N12097);
and and7024(N12105,N12111,R5);
and and7025(N12106,N12112,N12113);
and and7033(N12121,N12128,R5);
and and7034(N12122,R6,N12129);
and and7042(N12137,N12143,N12144);
and and7043(N12138,N12145,R7);
and and7051(N12153,N12159,N12160);
and and7052(N12154,R6,N12161);
and and7060(N12169,N12175,R4);
and and7061(N12170,N12176,N12177);
and and7069(N12185,N12191,N12192);
and and7070(N12186,N12193,R7);
and and7078(N12201,R4,N12206);
and and7079(N12202,N12207,N12208);
and and7087(N12216,R4,N12221);
and and7088(N12217,N12222,N12223);
and and7096(N12231,R4,N12236);
and and7097(N12232,N12237,N12238);
and and7105(N12246,N12251,N12252);
and and7106(N12247,N12253,R7);
and and7114(N12261,R4,R5);
and and7115(N12262,N12267,N12268);
and and7123(N12276,N12281,N12282);
and and7124(N12277,N12283,R7);
and and7132(N12291,N12296,N12297);
and and7133(N12292,R6,N12298);
and and7141(N12306,R4,R5);
and and7142(N12307,N12312,N12313);
and and7150(N12321,R4,R5);
and and7151(N12322,N12327,N12328);
and and7159(N12336,R4,R5);
and and7160(N12337,N12342,N12343);
and and7168(N12351,N12356,N12357);
and and7169(N12352,N12358,R7);
and and7177(N12366,N12371,N12372);
and and7178(N12367,N12373,R7);
and and7186(N12381,N12385,N12386);
and and7187(N12382,N12387,N12388);
and and7195(N12396,N12401,N12402);
and and7196(N12397,N12403,R7);
and and7204(N12411,N12416,R5);
and and7205(N12412,N12417,N12418);
and and7213(N12426,N12431,R5);
and and7214(N12427,N12432,N12433);
and and7222(N12441,N12446,R5);
and and7223(N12442,N12447,N12448);
and and7231(N12456,N12462,R5);
and and7232(N12457,R6,N12463);
and and7240(N12471,R3,N12477);
and and7241(N12472,R5,N12478);
and and7249(N12486,N12492,R5);
and and7250(N12487,N12493,R7);
and and7258(N12501,N12507,N12508);
and and7259(N12502,R6,R7);
and and7267(N12516,R4,R5);
and and7268(N12517,N12522,N12523);
and and7276(N12531,N12537,R5);
and and7277(N12532,N12538,R7);
and and7285(N12546,R4,N12552);
and and7286(N12547,N12553,R7);
and and7294(N12561,R4,N12567);
and and7295(N12562,R6,N12568);
and and7303(N12576,R4,N12581);
and and7304(N12577,N12582,N12583);
and and7312(N12591,R4,N12597);
and and7313(N12592,N12598,R7);
and and7321(N12606,R4,R5);
and and7322(N12607,N12612,N12613);
and and7330(N12621,R4,R5);
and and7331(N12622,N12627,N12628);
and and7339(N12636,R4,N12642);
and and7340(N12637,R6,N12643);
and and7348(N12651,R4,N12656);
and and7349(N12652,N12657,N12658);
and and7357(N12666,R4,N12671);
and and7358(N12667,N12672,N12673);
and and7366(N12681,R4,N12687);
and and7367(N12682,N12688,R7);
and and7375(N12696,N12701,R4);
and and7376(N12697,N12702,N12703);
and and7384(N12711,N12716,N12717);
and and7385(N12712,N12718,R7);
and and7393(N12726,N12731,R5);
and and7394(N12727,N12732,N12733);
and and7402(N12741,N12746,R5);
and and7403(N12742,N12747,N12748);
and and7411(N12756,R4,N12761);
and and7412(N12757,R6,N12762);
and and7420(N12770,R4,N12775);
and and7421(N12771,R6,N12776);
and and7429(N12784,R4,N12789);
and and7430(N12785,R6,N12790);
and and7438(N12798,R3,N12803);
and and7439(N12799,R6,N12804);
and and7447(N12812,N12816,N12817);
and and7448(N12813,R6,N12818);
and and7456(N12826,R3,N12831);
and and7457(N12827,R6,N12832);
and and7465(N12840,N12845,R5);
and and7466(N12841,R6,N12846);
and and7474(N12854,R4,R5);
and and7475(N12855,R6,N12860);
and and7483(N12868,N12873,R5);
and and7484(N12869,N12874,R7);
and and7492(N12882,N12887,R5);
and and7493(N12883,N12888,R7);
and and7501(N12896,N12901,R5);
and and7502(N12897,N12902,R7);
and and7510(N12910,N12914,N12915);
and and7511(N12911,R6,N12916);
and and7519(N12924,N12929,N12930);
and and7520(N12925,R6,R7);
and and7528(N12938,R4,R5);
and and7529(N12939,N12944,R7);
and and7537(N12952,R4,R5);
and and7538(N12953,N12958,R7);
and and7546(N12966,R4,N12971);
and and7547(N12967,N12972,R7);
and and7555(N12980,R4,N12985);
and and7556(N12981,R6,N12986);
and and7564(N12994,R4,N12999);
and and7565(N12995,N13000,R7);
and and7573(N13008,R3,R4);
and and7574(N13009,N13014,R7);
and and7582(N13022,N13026,N13027);
and and7583(N13023,N13028,R7);
and and7591(N13036,R4,N13040);
and and7592(N13037,N13041,N13042);
and and7600(N13050,R4,N13055);
and and7601(N13051,R6,N13056);
and and7609(N13064,N13069,N13070);
and and7610(N13065,R6,R7);
and and7618(N13078,R4,N13084);
and and7619(N13079,R6,R7);
and and7627(N13092,R3,N13098);
and and7628(N13093,R6,R7);
and and7636(N13106,R4,N13111);
and and7637(N13107,R6,N13112);
and and7645(N13120,N13125,R4);
and and7646(N13121,R6,N13126);
and and7654(N13134,N13138,N13139);
and and7655(N13135,N13140,R7);
and and7663(N13148,R3,N13153);
and and7664(N13149,N13154,R7);
and and7672(N13162,R3,N13167);
and and7673(N13163,N13168,R7);
and and7681(N13176,R4,R5);
and and7682(N13177,N13182,R7);
and and7690(N13190,N13194,N13195);
and and7691(N13191,R6,N13196);
and and7699(N13204,R4,N13209);
and and7700(N13205,R6,N13210);
and and7708(N13218,N13223,R4);
and and7709(N13219,R5,N13224);
and and7717(N13232,R3,R4);
and and7718(N13233,R6,N13238);
and and7726(N13246,R3,R4);
and and7727(N13247,R6,N13252);
and and7735(N13260,R3,R4);
and and7736(N13261,R5,N13266);
and and7744(N13274,N13279,R4);
and and7745(N13275,R5,N13280);
and and7753(N13288,R4,N13293);
and and7754(N13289,N13294,R7);
and and7762(N13302,R4,N13307);
and and7763(N13303,N13308,R7);
and and7771(N13316,R4,N13321);
and and7772(N13317,N13322,R7);
and and7780(N13330,R4,N13333);
and and7781(N13331,N13334,N13335);
and and7789(N13343,R4,N13346);
and and7790(N13344,N13347,N13348);
and and7798(N13356,N13360,R5);
and and7799(N13357,N13361,R7);
and and7807(N13369,R4,N13372);
and and7808(N13370,N13373,N13374);
and and7816(N13382,R3,R4);
and and7817(N13383,N13386,N13387);
and and7825(N13395,N13399,N13400);
and and7826(N13396,R6,R7);
and and7834(N13408,N13411,N13412);
and and7835(N13409,R6,N13413);
and and7843(N13421,R4,R5);
and and7844(N13422,N13425,N13426);
and and7852(N13434,N13436,N13437);
and and7853(N13435,N13438,N13439);
and and7861(N13447,R4,R5);
and and7862(N13448,N13452,R7);
and and7870(N13460,R3,N13464);
and and7871(N13461,R5,N13465);
and and7879(N13473,R3,N13477);
and and7880(N13474,R5,N13478);
and and7888(N13486,N13490,R5);
and and7889(N13487,N13491,R7);
and and7897(N13499,R4,R5);
and and7898(N13500,N13503,N13504);
and and7906(N13512,N13516,R5);
and and7907(N13513,R6,N13517);
and and7915(N13525,N13529,R5);
and and7916(N13526,R6,N13530);
and and7924(N13538,R4,R5);
and and7925(N13539,R6,N13543);
and and7933(N13551,R3,R4);
and and7934(N13552,R5,N13556);
and and7942(N13564,R4,R5);
and and7943(N13565,N13568,N13569);
and and7951(N13577,R4,R5);
and and7952(N13578,R6,N13582);
and and7960(N13590,R4,R5);
and and7961(N13591,N13594,N13595);
and and7969(N13603,R4,N13607);
and and7970(N13604,R6,N13608);
and and7978(N13616,R4,N13620);
and and7979(N13617,R6,N13621);
and and7987(N13629,N13632,N13633);
and and7988(N13630,N13634,R7);
and and7996(N13642,R4,N13647);
and and7997(N13643,R6,R7);
and and8005(N13655,R3,R4);
and and8006(N13656,N13659,N13660);
and and8014(N13668,R4,N13672);
and and8015(N13669,R6,N13673);
and and8023(N13681,R4,N13685);
and and8024(N13682,R6,N13686);
and and8032(N13694,N13698,R4);
and and8033(N13695,N13699,R7);
and and8041(N13707,R3,N13712);
and and8042(N13708,R6,R7);
and and8050(N13720,R4,R5);
and and8051(N13721,R6,N13725);
and and8059(N13733,R3,R4);
and and8060(N13734,R5,R6);
and and8068(N13746,N13749,N13750);
and and8069(N13747,N13751,R7);
and and8077(N13759,R3,N13763);
and and8078(N13760,N13764,R7);
and and8086(N13772,N13775,N13776);
and and8087(N13773,N13777,R7);
and and8095(N13785,R4,N13789);
and and8096(N13786,N13790,R7);
and and8104(N13798,N13801,N13802);
and and8105(N13799,N13803,R7);
and and8113(N13811,R4,N13815);
and and8114(N13812,R6,N13816);
and and8122(N13824,R4,N13828);
and and8123(N13825,R6,N13829);
and and8131(N13837,R4,N13841);
and and8132(N13838,R6,N13842);
and and8140(N13850,R4,N13854);
and and8141(N13851,R6,N13855);
and and8149(N13863,R4,R5);
and and8150(N13864,N13867,N13868);
and and8158(N13876,N13880,R4);
and and8159(N13877,R5,N13881);
and and8167(N13889,R4,R5);
and and8168(N13890,N13893,N13894);
and and8176(N13902,R4,N13906);
and and8177(N13903,N13907,R7);
and and8185(N13915,R4,N13919);
and and8186(N13916,N13920,R7);
and and8194(N13928,N13932,R4);
and and8195(N13929,R6,R7);
and and8203(N13940,N13943,N13944);
and and8204(N13941,R6,R7);
and and8212(N13952,R4,N13955);
and and8213(N13953,R6,N13956);
and and8221(N13964,R4,N13967);
and and8222(N13965,R6,N13968);
and and8230(N13976,N13978,N13979);
and and8231(N13977,R6,N13980);
and and8239(N13988,R4,R5);
and and8240(N13989,R6,N13992);
and and8248(N14000,R4,N14004);
and and8249(N14001,R6,R7);
and and8257(N14012,R4,N14015);
and and8258(N14013,N14016,R7);
and and8266(N14024,R4,N14027);
and and8267(N14025,N14028,R7);
and and8275(N14036,R3,R4);
and and8276(N14037,N14040,R7);
and and8284(N14048,R4,R5);
and and8285(N14049,R6,R7);
and and8293(N14060,N14064,R5);
and and8294(N14061,R6,R7);
and and8302(N14072,R4,R5);
and and8303(N14073,R6,R7);
and and8311(N14084,N14087,N14088);
and and8312(N14085,R6,R7);
and and8320(N14096,R3,R4);
and and8321(N14097,N14100,R6);
and and8329(N14108,R3,R4);
and and8330(N14109,R6,N14112);
and and8338(N14120,R4,N14123);
and and8339(N14121,R6,N14124);
and and8347(N14132,R4,N14135);
and and8348(N14133,R6,N14136);
and and8356(N14144,N14148,R5);
and and8357(N14145,R6,R7);
and and8365(N14156,N14160,R5);
and and8366(N14157,R6,R7);
and and8374(N14168,R4,R5);
and and8375(N14169,R6,N14172);
and and8383(N14180,R4,R5);
and and8384(N14181,R6,N14184);
and and8392(N14192,R4,N14196);
and and8393(N14193,R6,R7);
and and8401(N14204,R3,R4);
and and8402(N14205,R5,R6);
and and8410(N14216,R4,N14220);
and and8411(N14217,R6,R7);
and and8419(N14228,R4,R5);
and and8420(N14229,N14231,N14232);
and and8428(N14240,R3,N14244);
and and8429(N14241,R5,R6);
and and8437(N14252,N14256,R4);
and and8438(N14253,R6,R7);
and and8446(N14264,R3,R4);
and and8447(N14265,N14266,N14267);
and and8455(N14275,R3,R4);
and and8456(N14276,N14278,R7);
and and8464(N14286,N14288,R5);
and and8465(N14287,N14289,R7);
and and8473(N14297,R4,R5);
and and8474(N14298,R6,N14300);
and and8482(N14308,N14310,R5);
and and8483(N14309,R6,N14311);
and and8491(N14319,R3,R4);
and and8492(N14320,R5,R7);
and and8500(N14330,R4,R5);
and and8501(N14331,N14333,R7);
and and8509(N14341,R4,R5);
and and8510(N14342,N14343,N14344);
and and8518(N14352,R4,R5);
and and8519(N14353,N14354,N14355);
and and8527(N14363,R4,R5);
and and8528(N14364,N14366,R7);
and and8536(N14374,R4,N14377);
and and8537(N14375,R6,R7);
and and8545(N14385,R3,R4);
and and8546(N14386,N14388,R6);
and and8554(N14396,N14399,R5);
and and8555(N14397,R6,R7);
and and8563(N14407,R3,R4);
and and8564(N14408,R5,R7);
and and8572(N14418,N14420,R4);
and and8573(N14419,R5,N14421);
and and8581(N14429,R3,R4);
and and8582(N14430,R5,N14432);
and and8590(N14440,R4,N14442);
and and8591(N14441,R6,R7);
and and8599(N14450,R4,R5);
and and8600(N14451,R6,R7);
and and8608(N14460,R4,R5);
and and8609(N14461,R6,R7);
and and8617(N14470,N14472,R5);
and and8618(N14471,R6,R7);
and and8626(N14480,R4,R5);
and and8627(N14481,R6,R7);
and and8635(N14490,R4,N14492);
and and8636(N14491,R6,R7);
and and8644(N14500,R3,R4);
and and8645(N14501,R5,R7);
and and8653(N14509,N14516,N14517);
and and8661(N14525,N14532,N14533);
and and8669(N14541,N14548,N14549);
and and8677(N14557,N14564,R7);
and and8685(N14572,R6,N14579);
and and8693(N14587,R6,N14594);
and and8701(N14602,N14608,N14609);
and and8709(N14617,R6,N14624);
and and8717(N14632,N14638,N14639);
and and8725(N14647,N14653,N14654);
and and8733(N14662,N14668,N14669);
and and8741(N14677,N14683,N14684);
and and8749(N14692,N14698,N14699);
and and8757(N14707,N14712,N14713);
and and8765(N14721,N14727,R7);
and and8773(N14735,N14741,R6);
and and8781(N14749,N14755,R7);
and and8789(N14763,N14769,R7);
and and8797(N14777,N14782,N14783);
and and8805(N14791,R6,N14797);
and and8813(N14805,N14810,N14811);
and and8821(N14819,R6,N14825);
and and8829(N14833,N14839,R6);
and and8837(N14847,N14853,R6);
and and8845(N14861,N14866,N14867);
and and8853(N14875,R6,N14881);
and and8861(N14889,N14894,N14895);
and and8869(N14903,R6,N14909);
and and8877(N14917,N14922,N14923);
and and8885(N14931,N14936,N14937);
and and8893(N14945,R5,N14951);
and and8901(N14959,N14964,N14965);
and and8909(N14973,N14978,N14979);
and and8917(N14987,N14993,R7);
and and8925(N15001,N15007,R7);
and and8933(N15015,N15020,N15021);
and and8941(N15029,N15035,R7);
and and8949(N15043,N15049,R7);
and and8957(N15057,N15062,N15063);
and and8965(N15071,N15077,R7);
and and8973(N15085,N15090,N15091);
and and8981(N15099,R6,N15105);
and and8989(N15113,R6,N15119);
and and8997(N15127,N15132,N15133);
and and9005(N15141,R5,N15147);
and and9013(N15155,N15160,N15161);
and and9021(N15169,N15174,N15175);
and and9029(N15183,N15188,N15189);
and and9037(N15197,N15201,N15202);
and and9045(N15210,N15214,N15215);
and and9053(N15223,R6,N15228);
and and9061(N15236,N15240,N15241);
and and9069(N15249,R6,R7);
and and9077(N15262,N15266,N15267);
and and9085(N15275,N15279,N15280);
and and9093(N15288,N15292,N15293);
and and9101(N15301,R6,N15306);
and and9109(N15314,R6,N15319);
and and9117(N15327,N15331,N15332);
and and9125(N15340,R6,N15345);
and and9133(N15353,R6,N15358);
and and9141(N15366,N15370,N15371);
and and9149(N15379,R6,N15384);
and and9157(N15392,N15397,R7);
and and9165(N15405,R6,N15410);
and and9173(N15418,N15422,N15423);
and and9181(N15431,N15435,N15436);
and and9189(N15444,R6,N15449);
and and9197(N15457,R6,N15462);
and and9205(N15470,R5,N15475);
and and9213(N15483,N15487,N15488);
and and9221(N15496,N15500,N15501);
and and9229(N15509,R6,N15514);
and and9237(N15522,N15527,R7);
and and9245(N15535,R6,R7);
and and9253(N15548,N15553,R6);
and and9261(N15561,N15565,N15566);
and and9269(N15574,N15578,N15579);
and and9277(N15587,N15592,R7);
and and9285(N15600,R5,N15605);
and and9293(N15613,R6,N15618);
and and9301(N15626,N15631,R7);
and and9309(N15639,N15643,N15644);
and and9317(N15652,N15657,R7);
and and9325(N15665,R6,R7);
and and9333(N15678,N15683,R6);
and and9341(N15691,N15695,N15696);
and and9349(N15704,N15709,R7);
and and9357(N15717,N15722,R7);
and and9365(N15730,N15734,N15735);
and and9373(N15743,N15748,R7);
and and9381(N15756,N15761,R7);
and and9389(N15769,N15773,N15774);
and and9397(N15782,N15786,N15787);
and and9405(N15795,R6,R7);
and and9413(N15808,N15813,R7);
and and9421(N15821,R6,R7);
and and9429(N15833,N15836,N15837);
and and9437(N15845,N15849,R6);
and and9445(N15857,N15861,R7);
and and9453(N15869,N15873,R6);
and and9461(N15881,R6,N15885);
and and9469(N15893,R6,R7);
and and9477(N15905,R6,R7);
and and9485(N15917,N15921,R7);
and and9493(N15929,R6,N15933);
and and9501(N15941,R6,N15945);
and and9509(N15953,N15956,N15957);
and and9517(N15965,R6,N15969);
and and9525(N15977,N15981,R7);
and and9533(N15989,R6,R7);
and and9541(N16001,R6,R7);
and and9549(N16013,N16017,R7);
and and9557(N16025,R5,R7);
and and9565(N16037,N16041,R7);
and and9573(N16049,N16053,R7);
and and9581(N16061,R6,R7);
and and9589(N16073,N16076,N16077);
and and9597(N16085,N16088,N16089);
and and9605(N16097,R5,N16101);
and and9613(N16109,R6,N16113);
and and9621(N16121,N16125,R7);
and and9629(N16133,R6,R7);
and and9637(N16145,R6,R7);
and and9645(N16157,R6,R7);
and and9653(N16169,N16173,R6);
and and9661(N16181,N16185,R6);
and and9669(N16193,N16197,R7);
and and9677(N16205,N16208,N16209);
and and9685(N16217,R5,R6);
and and9693(N16229,N16232,N16233);
and and9701(N16241,N16245,R7);
and and9709(N16253,R5,N16257);
and and9717(N16265,N16268,N16269);
and and9725(N16277,N16281,R7);
and and9733(N16289,R6,N16293);
and and9741(N16301,N16305,R7);
and and9749(N16313,R6,R7);
and and9757(N16325,R6,N16329);
and and9765(N16337,N16340,N16341);
and and9773(N16349,N16353,R7);
and and9781(N16361,R6,R7);
and and9789(N16373,R6,N16377);
and and9797(N16385,R5,N16389);
and and9805(N16397,R5,N16401);
and and9813(N16409,N16412,N16413);
and and9821(N16421,N16424,N16425);
and and9829(N16433,N16436,N16437);
and and9837(N16445,N16449,R6);
and and9845(N16457,R6,R7);
and and9853(N16468,N16470,N16471);
and and9861(N16479,N16481,N16482);
and and9869(N16490,R5,N16493);
and and9877(N16501,N16504,R7);
and and9885(N16512,R6,R7);
and and9893(N16523,N16526,R7);
and and9901(N16534,N16537,R7);
and and9909(N16545,R6,N16548);
and and9917(N16556,R6,N16559);
and and9925(N16567,R6,N16570);
and and9933(N16578,R6,R7);
and and9941(N16589,R6,N16592);
and and9949(N16600,R6,N16603);
and and9957(N16611,R4,N16614);
and and9965(N16622,R5,N16625);
and and9973(N16633,R6,R7);
and and9981(N16644,N16647,R7);
and and9989(N16655,R6,R7);
and and9997(N16666,R5,N16669);
and and10005(N16677,N16680,R7);
and and10013(N16688,N16691,R6);
and and10021(N16699,R6,R7);
and and10029(N16710,R5,R7);
and and10037(N16721,N16724,R7);
and and10045(N16732,R5,R7);
and and10053(N16743,R5,N16746);
and and10061(N16754,N16757,R7);
and and10069(N16765,R6,R7);
and and10077(N16776,R6,N16779);
and and10085(N16787,N16790,R7);
and and10093(N16798,R6,N16801);
and and10101(N16809,R5,R6);
and and10109(N16820,R6,N16823);
and and10117(N16831,R6,N16834);
and and10125(N16842,R6,R7);
and and10133(N16853,R6,R7);
and and10141(N16864,N16866,N16867);
and and10149(N16875,N16877,N16878);
and and10157(N16886,R6,R7);
and and10165(N16897,N16899,R7);
and and10173(N16907,R6,R7);
and and10181(N16917,R6,R7);
and and10189(N16927,R5,N16929);
and and10197(N16937,R6,R7);
and and10205(N16947,R6,R7);
and and10213(N16957,R6,N16959);
and and10221(N16967,N16969,R7);
and and10229(N16977,N16979,R7);
and and10237(N16987,N16989,R7);
and and10245(N16997,R5,N16999);
and and10253(N17007,R5,R6);
and and10261(N17017,R6,R7);
and and10269(N17027,R4,R6);
and and10277(N17037,N17039,R6);
and and10285(N17047,R5,R6);
and and10293(N17057,N17059,R7);
and and10301(N17067,R5,R7);
and and10309(N17076,R6,R7);
and and10317(N17085,R6,R7);
and and10325(N17094,R6,R7);
and and10333(N17103,R6,R7);
and and10341(N17112,R5,R6);
and and10349(N17121,R5,R6);
and and10357(N17130,R6,R7);
and and10365(N17139,R5,R6);
and and10373(N17148,R5,R7);
and and10381(N17157,R5,R6);
and and10676(N18110,N18111,N18112);
and and10685(N18128,N18129,N18130);
and and10694(N18145,N18146,N18147);
and and10703(N18162,N18163,N18164);
and and10712(N18179,N18180,N18181);
and and10721(N18196,N18197,N18198);
and and10730(N18213,N18214,N18215);
and and10739(N18230,N18231,N18232);
and and10748(N18246,N18247,N18248);
and and10757(N18262,N18263,N18264);
and and10766(N18278,N18279,N18280);
and and10775(N18294,N18295,N18296);
and and10784(N18310,N18311,N18312);
and and10793(N18326,N18327,N18328);
and and10802(N18342,N18343,N18344);
and and10811(N18358,N18359,N18360);
and and10820(N18374,N18375,N18376);
and and10829(N18390,N18391,N18392);
and and10838(N18406,N18407,N18408);
and and10847(N18422,N18423,N18424);
and and10856(N18438,N18439,N18440);
and and10865(N18454,N18455,N18456);
and and10874(N18470,N18471,N18472);
and and10883(N18486,N18487,N18488);
and and10892(N18502,N18503,N18504);
and and10901(N18518,N18519,N18520);
and and10910(N18534,N18535,N18536);
and and10919(N18550,N18551,N18552);
and and10928(N18565,N18566,N18567);
and and10937(N18580,N18581,N18582);
and and10946(N18595,N18596,N18597);
and and10955(N18610,N18611,N18612);
and and10964(N18625,N18626,N18627);
and and10973(N18640,N18641,N18642);
and and10982(N18655,N18656,N18657);
and and10991(N18670,N18671,N18672);
and and11000(N18685,N18686,N18687);
and and11009(N18700,N18701,N18702);
and and11018(N18715,N18716,N18717);
and and11027(N18730,N18731,N18732);
and and11036(N18745,N18746,N18747);
and and11045(N18760,N18761,N18762);
and and11054(N18775,N18776,N18777);
and and11063(N18790,N18791,N18792);
and and11072(N18805,N18806,N18807);
and and11081(N18820,N18821,N18822);
and and11090(N18835,N18836,N18837);
and and11099(N18850,N18851,N18852);
and and11108(N18865,N18866,N18867);
and and11117(N18880,N18881,N18882);
and and11126(N18895,N18896,N18897);
and and11135(N18910,N18911,N18912);
and and11144(N18924,N18925,N18926);
and and11153(N18938,N18939,N18940);
and and11162(N18952,N18953,N18954);
and and11171(N18966,N18967,N18968);
and and11180(N18980,N18981,N18982);
and and11189(N18994,N18995,N18996);
and and11198(N19008,N19009,N19010);
and and11207(N19022,N19023,N19024);
and and11216(N19036,N19037,N19038);
and and11225(N19050,N19051,N19052);
and and11234(N19064,N19065,N19066);
and and11243(N19078,N19079,N19080);
and and11252(N19092,N19093,N19094);
and and11261(N19106,N19107,N19108);
and and11270(N19120,N19121,N19122);
and and11279(N19134,N19135,N19136);
and and11288(N19148,N19149,N19150);
and and11297(N19162,N19163,N19164);
and and11306(N19176,N19177,N19178);
and and11315(N19190,N19191,N19192);
and and11324(N19204,N19205,N19206);
and and11333(N19218,N19219,N19220);
and and11342(N19232,N19233,N19234);
and and11351(N19246,N19247,N19248);
and and11360(N19260,N19261,N19262);
and and11369(N19274,N19275,N19276);
and and11378(N19288,N19289,N19290);
and and11387(N19302,N19303,N19304);
and and11396(N19316,N19317,N19318);
and and11405(N19330,N19331,N19332);
and and11414(N19344,N19345,N19346);
and and11423(N19358,N19359,N19360);
and and11432(N19372,N19373,N19374);
and and11441(N19386,N19387,N19388);
and and11450(N19400,N19401,N19402);
and and11459(N19414,N19415,N19416);
and and11468(N19428,N19429,N19430);
and and11477(N19442,N19443,N19444);
and and11486(N19456,N19457,N19458);
and and11495(N19470,N19471,N19472);
and and11504(N19484,N19485,N19486);
and and11513(N19498,N19499,N19500);
and and11522(N19512,N19513,N19514);
and and11531(N19526,N19527,N19528);
and and11540(N19540,N19541,N19542);
and and11549(N19554,N19555,N19556);
and and11558(N19568,N19569,N19570);
and and11567(N19582,N19583,N19584);
and and11576(N19596,N19597,N19598);
and and11585(N19610,N19611,N19612);
and and11594(N19624,N19625,N19626);
and and11603(N19638,N19639,N19640);
and and11612(N19652,N19653,N19654);
and and11621(N19666,N19667,N19668);
and and11630(N19680,N19681,N19682);
and and11639(N19694,N19695,N19696);
and and11648(N19708,N19709,N19710);
and and11657(N19722,N19723,N19724);
and and11666(N19735,N19736,N19737);
and and11675(N19748,N19749,N19750);
and and11684(N19761,N19762,N19763);
and and11693(N19774,N19775,N19776);
and and11702(N19787,N19788,N19789);
and and11711(N19800,N19801,N19802);
and and11720(N19813,N19814,N19815);
and and11729(N19826,N19827,N19828);
and and11738(N19839,N19840,N19841);
and and11747(N19852,N19853,N19854);
and and11756(N19865,N19866,N19867);
and and11765(N19878,N19879,N19880);
and and11774(N19891,N19892,N19893);
and and11783(N19904,N19905,N19906);
and and11792(N19917,N19918,N19919);
and and11801(N19930,N19931,N19932);
and and11810(N19943,N19944,N19945);
and and11819(N19956,N19957,N19958);
and and11828(N19969,N19970,N19971);
and and11837(N19982,N19983,N19984);
and and11846(N19995,N19996,N19997);
and and11855(N20008,N20009,N20010);
and and11864(N20021,N20022,N20023);
and and11873(N20034,N20035,N20036);
and and11882(N20047,N20048,N20049);
and and11891(N20060,N20061,N20062);
and and11900(N20073,N20074,N20075);
and and11909(N20086,N20087,N20088);
and and11918(N20099,N20100,N20101);
and and11927(N20112,N20113,N20114);
and and11936(N20125,N20126,N20127);
and and11945(N20138,N20139,N20140);
and and11954(N20151,N20152,N20153);
and and11963(N20164,N20165,N20166);
and and11972(N20177,N20178,N20179);
and and11981(N20190,N20191,N20192);
and and11990(N20203,N20204,N20205);
and and11999(N20216,N20217,N20218);
and and12008(N20229,N20230,N20231);
and and12017(N20242,N20243,N20244);
and and12026(N20254,N20255,N20256);
and and12035(N20266,N20267,N20268);
and and12044(N20278,N20279,N20280);
and and12053(N20290,N20291,N20292);
and and12062(N20302,N20303,N20304);
and and12071(N20314,N20315,N20316);
and and12080(N20326,N20327,N20328);
and and12089(N20338,N20339,N20340);
and and12098(N20350,N20351,N20352);
and and12107(N20362,N20363,N20364);
and and12116(N20374,N20375,N20376);
and and12125(N20386,N20387,N20388);
and and12134(N20398,N20399,N20400);
and and12143(N20410,N20411,N20412);
and and12152(N20422,N20423,N20424);
and and12161(N20434,N20435,N20436);
and and12170(N20446,N20447,N20448);
and and12179(N20458,N20459,N20460);
and and12188(N20470,N20471,N20472);
and and12197(N20482,N20483,N20484);
and and12206(N20494,N20495,N20496);
and and12215(N20506,N20507,N20508);
and and12224(N20518,N20519,N20520);
and and12233(N20530,N20531,N20532);
and and12242(N20542,N20543,N20544);
and and12251(N20554,N20555,N20556);
and and12260(N20566,N20567,N20568);
and and12269(N20578,N20579,N20580);
and and12278(N20590,N20591,N20592);
and and12287(N20602,N20603,N20604);
and and12296(N20614,N20615,N20616);
and and12305(N20626,N20627,N20628);
and and12314(N20638,N20639,N20640);
and and12323(N20650,N20651,N20652);
and and12332(N20662,N20663,N20664);
and and12341(N20673,N20674,N20675);
and and12350(N20684,N20685,N20686);
and and12359(N20695,N20696,N20697);
and and12368(N20706,N20707,N20708);
and and12377(N20717,N20718,N20719);
and and12386(N20728,N20729,N20730);
and and12395(N20738,N20739,N20740);
and and12404(N20748,N20749,N20750);
and and12413(N20758,N20759,N20760);
and and12422(N20768,N20769,N20770);
and and12431(N20778,N20779,N20780);
and and12440(N20788,N20789,N20790);
and and12449(N20798,N20799,N20800);
and and12458(N20808,N20809,N20810);
and and12467(N20818,N20819,N20820);
and and12476(N20828,N20829,N20830);
and and12485(N20838,N20839,N20840);
and and12494(N20848,N20849,N20850);
and and12502(N20864,N20865,N20866);
and and12510(N20880,N20881,N20882);
and and12518(N20895,N20896,N20897);
and and12526(N20910,N20911,N20912);
and and12534(N20925,N20926,N20927);
and and12542(N20940,N20941,N20942);
and and12550(N20955,N20956,N20957);
and and12558(N20970,N20971,N20972);
and and12566(N20985,N20986,N20987);
and and12574(N21000,N21001,N21002);
and and12582(N21015,N21016,N21017);
and and12590(N21030,N21031,N21032);
and and12598(N21045,N21046,N21047);
and and12606(N21060,N21061,N21062);
and and12614(N21075,N21076,N21077);
and and12622(N21089,N21090,N21091);
and and12630(N21103,N21104,N21105);
and and12638(N21117,N21118,N21119);
and and12646(N21131,N21132,N21133);
and and12654(N21145,N21146,N21147);
and and12662(N21159,N21160,N21161);
and and12670(N21173,N21174,N21175);
and and12678(N21187,N21188,N21189);
and and12686(N21201,N21202,N21203);
and and12694(N21215,N21216,N21217);
and and12702(N21229,N21230,N21231);
and and12710(N21243,N21244,N21245);
and and12718(N21257,N21258,N21259);
and and12726(N21271,N21272,N21273);
and and12734(N21285,N21286,N21287);
and and12742(N21299,N21300,N21301);
and and12750(N21313,N21314,N21315);
and and12758(N21327,N21328,N21329);
and and12766(N21341,N21342,N21343);
and and12774(N21355,N21356,N21357);
and and12782(N21369,N21370,N21371);
and and12790(N21383,N21384,N21385);
and and12798(N21397,N21398,N21399);
and and12806(N21411,N21412,N21413);
and and12814(N21425,N21426,N21427);
and and12822(N21439,N21440,N21441);
and and12830(N21453,N21454,N21455);
and and12838(N21467,N21468,N21469);
and and12846(N21481,N21482,N21483);
and and12854(N21495,N21496,N21497);
and and12862(N21509,N21510,N21511);
and and12870(N21523,N21524,N21525);
and and12878(N21536,N21537,N21538);
and and12886(N21549,N21550,N21551);
and and12894(N21562,N21563,N21564);
and and12902(N21575,N21576,N21577);
and and12910(N21588,N21589,N21590);
and and12918(N21601,N21602,N21603);
and and12926(N21614,N21615,N21616);
and and12934(N21627,N21628,N21629);
and and12942(N21640,N21641,N21642);
and and12950(N21653,N21654,N21655);
and and12958(N21666,N21667,N21668);
and and12966(N21679,N21680,N21681);
and and12974(N21692,N21693,N21694);
and and12982(N21705,N21706,N21707);
and and12990(N21718,N21719,N21720);
and and12998(N21731,N21732,N21733);
and and13006(N21744,N21745,N21746);
and and13014(N21757,N21758,N21759);
and and13022(N21770,N21771,N21772);
and and13030(N21783,N21784,N21785);
and and13038(N21796,N21797,N21798);
and and13046(N21809,N21810,N21811);
and and13054(N21822,N21823,N21824);
and and13062(N21835,N21836,N21837);
and and13070(N21848,N21849,N21850);
and and13078(N21861,N21862,N21863);
and and13086(N21874,N21875,N21876);
and and13094(N21887,N21888,N21889);
and and13102(N21900,N21901,N21902);
and and13110(N21913,N21914,N21915);
and and13118(N21926,N21927,N21928);
and and13126(N21939,N21940,N21941);
and and13134(N21952,N21953,N21954);
and and13142(N21965,N21966,N21967);
and and13150(N21978,N21979,N21980);
and and13158(N21991,N21992,N21993);
and and13166(N22004,N22005,N22006);
and and13174(N22017,N22018,N22019);
and and13182(N22030,N22031,N22032);
and and13190(N22043,N22044,N22045);
and and13198(N22056,N22057,N22058);
and and13206(N22069,N22070,N22071);
and and13214(N22082,N22083,N22084);
and and13222(N22095,N22096,N22097);
and and13230(N22108,N22109,N22110);
and and13238(N22121,N22122,N22123);
and and13246(N22134,N22135,N22136);
and and13254(N22147,N22148,N22149);
and and13262(N22160,N22161,N22162);
and and13270(N22173,N22174,N22175);
and and13278(N22186,N22187,N22188);
and and13286(N22199,N22200,N22201);
and and13294(N22212,N22213,N22214);
and and13302(N22225,N22226,N22227);
and and13310(N22237,N22238,N22239);
and and13318(N22249,N22250,N22251);
and and13326(N22261,N22262,N22263);
and and13334(N22273,N22274,N22275);
and and13342(N22285,N22286,N22287);
and and13350(N22297,N22298,N22299);
and and13358(N22309,N22310,N22311);
and and13366(N22321,N22322,N22323);
and and13374(N22333,N22334,N22335);
and and13382(N22345,N22346,N22347);
and and13390(N22357,N22358,N22359);
and and13398(N22369,N22370,N22371);
and and13406(N22381,N22382,N22383);
and and13414(N22393,N22394,N22395);
and and13422(N22405,N22406,N22407);
and and13430(N22417,N22418,N22419);
and and13438(N22429,N22430,N22431);
and and13446(N22441,N22442,N22443);
and and13454(N22453,N22454,N22455);
and and13462(N22465,N22466,N22467);
and and13470(N22477,N22478,N22479);
and and13478(N22489,N22490,N22491);
and and13486(N22501,N22502,N22503);
and and13494(N22513,N22514,N22515);
and and13502(N22525,N22526,N22527);
and and13510(N22537,N22538,N22539);
and and13518(N22549,N22550,N22551);
and and13526(N22561,N22562,N22563);
and and13534(N22573,N22574,N22575);
and and13542(N22585,N22586,N22587);
and and13550(N22597,N22598,N22599);
and and13558(N22609,N22610,N22611);
and and13566(N22621,N22622,N22623);
and and13574(N22633,N22634,N22635);
and and13582(N22645,N22646,N22647);
and and13590(N22657,N22658,N22659);
and and13598(N22669,N22670,N22671);
and and13606(N22681,N22682,N22683);
and and13614(N22693,N22694,N22695);
and and13622(N22705,N22706,N22707);
and and13630(N22717,N22718,N22719);
and and13638(N22729,N22730,N22731);
and and13646(N22741,N22742,N22743);
and and13654(N22753,N22754,N22755);
and and13662(N22765,N22766,N22767);
and and13670(N22777,N22778,N22779);
and and13678(N22789,N22790,N22791);
and and13686(N22801,N22802,N22803);
and and13694(N22813,N22814,N22815);
and and13702(N22825,N22826,N22827);
and and13710(N22836,N22837,N22838);
and and13718(N22847,N22848,N22849);
and and13726(N22858,N22859,N22860);
and and13734(N22869,N22870,N22871);
and and13742(N22880,N22881,N22882);
and and13750(N22891,N22892,N22893);
and and13758(N22902,N22903,N22904);
and and13766(N22913,N22914,N22915);
and and13774(N22924,N22925,N22926);
and and13782(N22935,N22936,N22937);
and and13790(N22946,N22947,N22948);
and and13798(N22957,N22958,N22959);
and and13806(N22968,N22969,N22970);
and and13814(N22979,N22980,N22981);
and and13822(N22990,N22991,N22992);
and and13830(N23001,N23002,N23003);
and and13838(N23012,N23013,N23014);
and and13846(N23023,N23024,N23025);
and and13854(N23034,N23035,N23036);
and and13862(N23045,N23046,N23047);
and and13870(N23056,N23057,N23058);
and and13878(N23067,N23068,N23069);
and and13886(N23078,N23079,N23080);
and and13894(N23089,N23090,N23091);
and and13902(N23100,N23101,N23102);
and and13910(N23111,N23112,N23113);
and and13918(N23122,N23123,N23124);
and and13926(N23133,N23134,N23135);
and and13934(N23144,N23145,N23146);
and and13942(N23155,N23156,N23157);
and and13950(N23166,N23167,N23168);
and and13958(N23177,N23178,N23179);
and and13966(N23188,N23189,N23190);
and and13974(N23199,N23200,N23201);
and and13982(N23210,N23211,N23212);
and and13990(N23221,N23222,N23223);
and and13998(N23232,N23233,N23234);
and and14006(N23243,N23244,N23245);
and and14014(N23254,N23255,N23256);
and and14022(N23265,N23266,N23267);
and and14030(N23276,N23277,N23278);
and and14038(N23287,N23288,N23289);
and and14046(N23298,N23299,N23300);
and and14054(N23309,N23310,N23311);
and and14062(N23320,N23321,N23322);
and and14070(N23331,N23332,N23333);
and and14078(N23342,N23343,N23344);
and and14086(N23353,N23354,N23355);
and and14094(N23364,N23365,N23366);
and and14102(N23375,N23376,N23377);
and and14110(N23386,N23387,N23388);
and and14118(N23397,N23398,N23399);
and and14126(N23407,N23408,N23409);
and and14134(N23417,N23418,N23419);
and and14142(N23427,N23428,N23429);
and and14150(N23437,N23438,N23439);
and and14158(N23447,N23448,N23449);
and and14166(N23457,N23458,N23459);
and and14174(N23467,N23468,N23469);
and and14182(N23477,N23478,N23479);
and and14190(N23487,N23488,N23489);
and and14198(N23497,N23498,N23499);
and and14206(N23507,N23508,N23509);
and and14214(N23517,N23518,N23519);
and and14222(N23527,N23528,N23529);
and and14230(N23537,N23538,N23539);
and and14238(N23547,N23548,N23549);
and and14246(N23556,N23557,N23558);
and and14254(N23565,N23566,N23567);
and and14262(N23574,N23575,N23576);
and and14270(N23583,N23584,N23585);
and and14278(N23592,N23593,N23594);
and and14286(N23601,N23602,N23603);
and and14294(N23610,N23611,N23612);
and and14302(N23619,N23620,N23621);
and and14310(N23628,N23629,N23630);
and and14318(N23636,N23637,N23638);
and and14325(N23650,N23651,N23652);
and and14332(N23664,N23665,N23666);
and and14339(N23677,N23678,N23679);
and and14346(N23690,N23691,N23692);
and and14353(N23703,N23704,N23705);
and and14360(N23716,N23717,N23718);
and and14367(N23729,N23730,N23731);
and and14374(N23742,N23743,N23744);
and and14381(N23754,N23755,N23756);
and and14388(N23766,N23767,N23768);
and and14395(N23778,N23779,N23780);
and and14402(N23790,N23791,N23792);
and and14409(N23802,N23803,N23804);
and and14416(N23814,N23815,N23816);
and and14423(N23826,N23827,N23828);
and and14430(N23838,N23839,N23840);
and and14437(N23850,N23851,N23852);
and and14444(N23861,N23862,N23863);
and and14451(N23872,N23873,N23874);
and and14458(N23883,N23884,N23885);
and and14465(N23894,N23895,N23896);
and and14472(N23905,N23906,N23907);
and and14479(N23916,N23917,N23918);
and and14486(N23927,N23928,N23929);
and and14493(N23938,N23939,N23940);
and and14500(N23948,N23949,N23950);
and and14507(N23958,N23959,N23960);
and and14514(N23968,N23969,N23970);
and and14521(N23978,N23979,N23980);
and and14528(N23988,N23989,N23990);
and and14535(N23998,N23999,N24000);
and and14542(N24008,N24009,N24010);
and and14549(N24018,N24019,N24020);
and and14556(N24028,N24029,N24030);
and and14563(N24038,N24039,N24040);
and and14570(N24047,N24048,N24049);
and and10677(N18111,N18113,N18114);
and and10678(N18112,N18115,N18116);
and and10686(N18129,N18131,N18132);
and and10687(N18130,N18133,N18134);
and and10695(N18146,N18148,N18149);
and and10696(N18147,N18150,N18151);
and and10704(N18163,N18165,N18166);
and and10705(N18164,N18167,N18168);
and and10713(N18180,N18182,N18183);
and and10714(N18181,N18184,N18185);
and and10722(N18197,N18199,N18200);
and and10723(N18198,N18201,N18202);
and and10731(N18214,N18216,N18217);
and and10732(N18215,N18218,N18219);
and and10740(N18231,N18233,N18234);
and and10741(N18232,N18235,N18236);
and and10749(N18247,N18249,N18250);
and and10750(N18248,N18251,N18252);
and and10758(N18263,N18265,N18266);
and and10759(N18264,N18267,N18268);
and and10767(N18279,N18281,N18282);
and and10768(N18280,N18283,N18284);
and and10776(N18295,N18297,N18298);
and and10777(N18296,N18299,N18300);
and and10785(N18311,N18313,N18314);
and and10786(N18312,N18315,N18316);
and and10794(N18327,N18329,N18330);
and and10795(N18328,N18331,N18332);
and and10803(N18343,N18345,N18346);
and and10804(N18344,N18347,N18348);
and and10812(N18359,N18361,N18362);
and and10813(N18360,N18363,N18364);
and and10821(N18375,N18377,N18378);
and and10822(N18376,N18379,N18380);
and and10830(N18391,N18393,N18394);
and and10831(N18392,N18395,N18396);
and and10839(N18407,N18409,N18410);
and and10840(N18408,N18411,N18412);
and and10848(N18423,N18425,N18426);
and and10849(N18424,N18427,N18428);
and and10857(N18439,N18441,N18442);
and and10858(N18440,N18443,N18444);
and and10866(N18455,N18457,N18458);
and and10867(N18456,N18459,N18460);
and and10875(N18471,N18473,N18474);
and and10876(N18472,N18475,N18476);
and and10884(N18487,N18489,N18490);
and and10885(N18488,N18491,N18492);
and and10893(N18503,N18505,N18506);
and and10894(N18504,N18507,N18508);
and and10902(N18519,N18521,N18522);
and and10903(N18520,N18523,N18524);
and and10911(N18535,N18537,N18538);
and and10912(N18536,N18539,N18540);
and and10920(N18551,N18553,N18554);
and and10921(N18552,N18555,N18556);
and and10929(N18566,N18568,N18569);
and and10930(N18567,N18570,N18571);
and and10938(N18581,N18583,N18584);
and and10939(N18582,N18585,N18586);
and and10947(N18596,N18598,N18599);
and and10948(N18597,N18600,N18601);
and and10956(N18611,N18613,N18614);
and and10957(N18612,N18615,N18616);
and and10965(N18626,N18628,N18629);
and and10966(N18627,N18630,N18631);
and and10974(N18641,N18643,N18644);
and and10975(N18642,N18645,N18646);
and and10983(N18656,N18658,N18659);
and and10984(N18657,N18660,N18661);
and and10992(N18671,N18673,N18674);
and and10993(N18672,N18675,N18676);
and and11001(N18686,N18688,N18689);
and and11002(N18687,N18690,N18691);
and and11010(N18701,N18703,N18704);
and and11011(N18702,N18705,N18706);
and and11019(N18716,N18718,N18719);
and and11020(N18717,N18720,N18721);
and and11028(N18731,N18733,N18734);
and and11029(N18732,N18735,N18736);
and and11037(N18746,N18748,N18749);
and and11038(N18747,N18750,N18751);
and and11046(N18761,N18763,N18764);
and and11047(N18762,N18765,N18766);
and and11055(N18776,N18778,N18779);
and and11056(N18777,N18780,N18781);
and and11064(N18791,N18793,N18794);
and and11065(N18792,N18795,N18796);
and and11073(N18806,N18808,N18809);
and and11074(N18807,N18810,N18811);
and and11082(N18821,N18823,N18824);
and and11083(N18822,N18825,N18826);
and and11091(N18836,N18838,N18839);
and and11092(N18837,N18840,N18841);
and and11100(N18851,N18853,N18854);
and and11101(N18852,N18855,N18856);
and and11109(N18866,N18868,N18869);
and and11110(N18867,N18870,N18871);
and and11118(N18881,N18883,N18884);
and and11119(N18882,N18885,N18886);
and and11127(N18896,N18898,N18899);
and and11128(N18897,N18900,N18901);
and and11136(N18911,N18913,N18914);
and and11137(N18912,N18915,N18916);
and and11145(N18925,N18927,N18928);
and and11146(N18926,N18929,N18930);
and and11154(N18939,N18941,N18942);
and and11155(N18940,N18943,N18944);
and and11163(N18953,N18955,N18956);
and and11164(N18954,N18957,N18958);
and and11172(N18967,N18969,N18970);
and and11173(N18968,N18971,N18972);
and and11181(N18981,N18983,N18984);
and and11182(N18982,N18985,N18986);
and and11190(N18995,N18997,N18998);
and and11191(N18996,N18999,N19000);
and and11199(N19009,N19011,N19012);
and and11200(N19010,N19013,N19014);
and and11208(N19023,N19025,N19026);
and and11209(N19024,N19027,N19028);
and and11217(N19037,N19039,N19040);
and and11218(N19038,N19041,N19042);
and and11226(N19051,N19053,N19054);
and and11227(N19052,N19055,N19056);
and and11235(N19065,N19067,N19068);
and and11236(N19066,N19069,N19070);
and and11244(N19079,N19081,N19082);
and and11245(N19080,N19083,N19084);
and and11253(N19093,N19095,N19096);
and and11254(N19094,N19097,N19098);
and and11262(N19107,N19109,N19110);
and and11263(N19108,N19111,N19112);
and and11271(N19121,N19123,N19124);
and and11272(N19122,N19125,N19126);
and and11280(N19135,N19137,N19138);
and and11281(N19136,N19139,N19140);
and and11289(N19149,N19151,N19152);
and and11290(N19150,N19153,N19154);
and and11298(N19163,N19165,N19166);
and and11299(N19164,N19167,N19168);
and and11307(N19177,N19179,N19180);
and and11308(N19178,N19181,N19182);
and and11316(N19191,N19193,N19194);
and and11317(N19192,N19195,N19196);
and and11325(N19205,N19207,N19208);
and and11326(N19206,N19209,N19210);
and and11334(N19219,N19221,N19222);
and and11335(N19220,N19223,N19224);
and and11343(N19233,N19235,N19236);
and and11344(N19234,N19237,N19238);
and and11352(N19247,N19249,N19250);
and and11353(N19248,N19251,N19252);
and and11361(N19261,N19263,N19264);
and and11362(N19262,N19265,N19266);
and and11370(N19275,N19277,N19278);
and and11371(N19276,N19279,N19280);
and and11379(N19289,N19291,N19292);
and and11380(N19290,N19293,N19294);
and and11388(N19303,N19305,N19306);
and and11389(N19304,N19307,N19308);
and and11397(N19317,N19319,N19320);
and and11398(N19318,N19321,N19322);
and and11406(N19331,N19333,N19334);
and and11407(N19332,N19335,N19336);
and and11415(N19345,N19347,N19348);
and and11416(N19346,N19349,N19350);
and and11424(N19359,N19361,N19362);
and and11425(N19360,N19363,N19364);
and and11433(N19373,N19375,N19376);
and and11434(N19374,N19377,N19378);
and and11442(N19387,N19389,N19390);
and and11443(N19388,N19391,N19392);
and and11451(N19401,N19403,N19404);
and and11452(N19402,N19405,N19406);
and and11460(N19415,N19417,N19418);
and and11461(N19416,N19419,N19420);
and and11469(N19429,N19431,N19432);
and and11470(N19430,N19433,N19434);
and and11478(N19443,N19445,N19446);
and and11479(N19444,N19447,N19448);
and and11487(N19457,N19459,N19460);
and and11488(N19458,N19461,N19462);
and and11496(N19471,N19473,N19474);
and and11497(N19472,N19475,N19476);
and and11505(N19485,N19487,N19488);
and and11506(N19486,N19489,N19490);
and and11514(N19499,N19501,N19502);
and and11515(N19500,N19503,N19504);
and and11523(N19513,N19515,N19516);
and and11524(N19514,N19517,N19518);
and and11532(N19527,N19529,N19530);
and and11533(N19528,N19531,N19532);
and and11541(N19541,N19543,N19544);
and and11542(N19542,N19545,N19546);
and and11550(N19555,N19557,N19558);
and and11551(N19556,N19559,N19560);
and and11559(N19569,N19571,N19572);
and and11560(N19570,N19573,N19574);
and and11568(N19583,N19585,N19586);
and and11569(N19584,N19587,N19588);
and and11577(N19597,N19599,N19600);
and and11578(N19598,N19601,N19602);
and and11586(N19611,N19613,N19614);
and and11587(N19612,N19615,N19616);
and and11595(N19625,N19627,N19628);
and and11596(N19626,N19629,N19630);
and and11604(N19639,N19641,N19642);
and and11605(N19640,N19643,N19644);
and and11613(N19653,N19655,N19656);
and and11614(N19654,N19657,N19658);
and and11622(N19667,N19669,N19670);
and and11623(N19668,N19671,N19672);
and and11631(N19681,N19683,N19684);
and and11632(N19682,N19685,N19686);
and and11640(N19695,N19697,N19698);
and and11641(N19696,N19699,N19700);
and and11649(N19709,N19711,N19712);
and and11650(N19710,N19713,N19714);
and and11658(N19723,N19725,N19726);
and and11659(N19724,N19727,N19728);
and and11667(N19736,N19738,N19739);
and and11668(N19737,N19740,N19741);
and and11676(N19749,N19751,N19752);
and and11677(N19750,N19753,N19754);
and and11685(N19762,N19764,N19765);
and and11686(N19763,N19766,N19767);
and and11694(N19775,N19777,N19778);
and and11695(N19776,N19779,N19780);
and and11703(N19788,N19790,N19791);
and and11704(N19789,N19792,N19793);
and and11712(N19801,N19803,N19804);
and and11713(N19802,N19805,N19806);
and and11721(N19814,N19816,N19817);
and and11722(N19815,N19818,N19819);
and and11730(N19827,N19829,N19830);
and and11731(N19828,N19831,N19832);
and and11739(N19840,N19842,N19843);
and and11740(N19841,N19844,N19845);
and and11748(N19853,N19855,N19856);
and and11749(N19854,N19857,N19858);
and and11757(N19866,N19868,N19869);
and and11758(N19867,N19870,N19871);
and and11766(N19879,N19881,N19882);
and and11767(N19880,N19883,N19884);
and and11775(N19892,N19894,N19895);
and and11776(N19893,N19896,N19897);
and and11784(N19905,N19907,N19908);
and and11785(N19906,N19909,N19910);
and and11793(N19918,N19920,N19921);
and and11794(N19919,N19922,N19923);
and and11802(N19931,N19933,N19934);
and and11803(N19932,N19935,N19936);
and and11811(N19944,N19946,N19947);
and and11812(N19945,N19948,N19949);
and and11820(N19957,N19959,N19960);
and and11821(N19958,N19961,N19962);
and and11829(N19970,N19972,N19973);
and and11830(N19971,N19974,N19975);
and and11838(N19983,N19985,N19986);
and and11839(N19984,N19987,N19988);
and and11847(N19996,N19998,N19999);
and and11848(N19997,N20000,N20001);
and and11856(N20009,N20011,N20012);
and and11857(N20010,N20013,N20014);
and and11865(N20022,N20024,N20025);
and and11866(N20023,N20026,N20027);
and and11874(N20035,N20037,N20038);
and and11875(N20036,N20039,N20040);
and and11883(N20048,N20050,N20051);
and and11884(N20049,N20052,N20053);
and and11892(N20061,N20063,N20064);
and and11893(N20062,N20065,N20066);
and and11901(N20074,N20076,N20077);
and and11902(N20075,N20078,N20079);
and and11910(N20087,N20089,N20090);
and and11911(N20088,N20091,N20092);
and and11919(N20100,N20102,N20103);
and and11920(N20101,N20104,N20105);
and and11928(N20113,N20115,N20116);
and and11929(N20114,N20117,N20118);
and and11937(N20126,N20128,N20129);
and and11938(N20127,N20130,N20131);
and and11946(N20139,N20141,N20142);
and and11947(N20140,N20143,N20144);
and and11955(N20152,N20154,N20155);
and and11956(N20153,N20156,N20157);
and and11964(N20165,N20167,N20168);
and and11965(N20166,N20169,N20170);
and and11973(N20178,N20180,N20181);
and and11974(N20179,N20182,N20183);
and and11982(N20191,N20193,N20194);
and and11983(N20192,N20195,N20196);
and and11991(N20204,N20206,N20207);
and and11992(N20205,N20208,N20209);
and and12000(N20217,N20219,N20220);
and and12001(N20218,N20221,N20222);
and and12009(N20230,N20232,N20233);
and and12010(N20231,N20234,N20235);
and and12018(N20243,N20245,N20246);
and and12019(N20244,N20247,N20248);
and and12027(N20255,N20257,N20258);
and and12028(N20256,N20259,N20260);
and and12036(N20267,N20269,N20270);
and and12037(N20268,N20271,N20272);
and and12045(N20279,N20281,N20282);
and and12046(N20280,N20283,N20284);
and and12054(N20291,N20293,N20294);
and and12055(N20292,N20295,N20296);
and and12063(N20303,N20305,N20306);
and and12064(N20304,N20307,N20308);
and and12072(N20315,N20317,N20318);
and and12073(N20316,N20319,N20320);
and and12081(N20327,N20329,N20330);
and and12082(N20328,N20331,N20332);
and and12090(N20339,N20341,N20342);
and and12091(N20340,N20343,N20344);
and and12099(N20351,N20353,N20354);
and and12100(N20352,N20355,N20356);
and and12108(N20363,N20365,N20366);
and and12109(N20364,N20367,N20368);
and and12117(N20375,N20377,N20378);
and and12118(N20376,N20379,N20380);
and and12126(N20387,N20389,N20390);
and and12127(N20388,N20391,N20392);
and and12135(N20399,N20401,N20402);
and and12136(N20400,N20403,N20404);
and and12144(N20411,N20413,N20414);
and and12145(N20412,N20415,N20416);
and and12153(N20423,N20425,N20426);
and and12154(N20424,N20427,N20428);
and and12162(N20435,N20437,N20438);
and and12163(N20436,N20439,N20440);
and and12171(N20447,N20449,N20450);
and and12172(N20448,N20451,N20452);
and and12180(N20459,N20461,N20462);
and and12181(N20460,N20463,N20464);
and and12189(N20471,N20473,N20474);
and and12190(N20472,N20475,N20476);
and and12198(N20483,N20485,N20486);
and and12199(N20484,N20487,N20488);
and and12207(N20495,N20497,N20498);
and and12208(N20496,N20499,N20500);
and and12216(N20507,N20509,N20510);
and and12217(N20508,N20511,N20512);
and and12225(N20519,N20521,N20522);
and and12226(N20520,N20523,N20524);
and and12234(N20531,N20533,N20534);
and and12235(N20532,N20535,N20536);
and and12243(N20543,N20545,N20546);
and and12244(N20544,N20547,N20548);
and and12252(N20555,N20557,N20558);
and and12253(N20556,N20559,N20560);
and and12261(N20567,N20569,N20570);
and and12262(N20568,N20571,N20572);
and and12270(N20579,N20581,N20582);
and and12271(N20580,N20583,N20584);
and and12279(N20591,N20593,N20594);
and and12280(N20592,N20595,N20596);
and and12288(N20603,N20605,N20606);
and and12289(N20604,N20607,N20608);
and and12297(N20615,N20617,N20618);
and and12298(N20616,N20619,N20620);
and and12306(N20627,N20629,N20630);
and and12307(N20628,N20631,N20632);
and and12315(N20639,N20641,N20642);
and and12316(N20640,N20643,N20644);
and and12324(N20651,N20653,N20654);
and and12325(N20652,N20655,N20656);
and and12333(N20663,N20665,N20666);
and and12334(N20664,N20667,N20668);
and and12342(N20674,N20676,N20677);
and and12343(N20675,N20678,N20679);
and and12351(N20685,N20687,N20688);
and and12352(N20686,N20689,N20690);
and and12360(N20696,N20698,N20699);
and and12361(N20697,N20700,N20701);
and and12369(N20707,N20709,N20710);
and and12370(N20708,N20711,N20712);
and and12378(N20718,N20720,N20721);
and and12379(N20719,N20722,N20723);
and and12387(N20729,N20731,N20732);
and and12388(N20730,N20733,N20734);
and and12396(N20739,N20741,N20742);
and and12397(N20740,N20743,N20744);
and and12405(N20749,N20751,N20752);
and and12406(N20750,N20753,N20754);
and and12414(N20759,N20761,N20762);
and and12415(N20760,N20763,N20764);
and and12423(N20769,N20771,N20772);
and and12424(N20770,N20773,N20774);
and and12432(N20779,N20781,N20782);
and and12433(N20780,N20783,N20784);
and and12441(N20789,N20791,N20792);
and and12442(N20790,N20793,N20794);
and and12450(N20799,N20801,N20802);
and and12451(N20800,N20803,N20804);
and and12459(N20809,N20811,N20812);
and and12460(N20810,N20813,N20814);
and and12468(N20819,N20821,N20822);
and and12469(N20820,N20823,N20824);
and and12477(N20829,N20831,N20832);
and and12478(N20830,N20833,N20834);
and and12486(N20839,N20841,N20842);
and and12487(N20840,N20843,N20844);
and and12495(N20849,N20851,N20852);
and and12496(N20850,N20853,N20854);
and and12503(N20865,N20867,N20868);
and and12504(N20866,N20869,N20870);
and and12511(N20881,N20883,N20884);
and and12512(N20882,N20885,N20886);
and and12519(N20896,N20898,N20899);
and and12520(N20897,N20900,N20901);
and and12527(N20911,N20913,N20914);
and and12528(N20912,N20915,N20916);
and and12535(N20926,N20928,N20929);
and and12536(N20927,N20930,N20931);
and and12543(N20941,N20943,N20944);
and and12544(N20942,N20945,N20946);
and and12551(N20956,N20958,N20959);
and and12552(N20957,N20960,N20961);
and and12559(N20971,N20973,N20974);
and and12560(N20972,N20975,N20976);
and and12567(N20986,N20988,N20989);
and and12568(N20987,N20990,N20991);
and and12575(N21001,N21003,N21004);
and and12576(N21002,N21005,N21006);
and and12583(N21016,N21018,N21019);
and and12584(N21017,N21020,N21021);
and and12591(N21031,N21033,N21034);
and and12592(N21032,N21035,N21036);
and and12599(N21046,N21048,N21049);
and and12600(N21047,N21050,N21051);
and and12607(N21061,N21063,N21064);
and and12608(N21062,N21065,N21066);
and and12615(N21076,N21078,N21079);
and and12616(N21077,N21080,N21081);
and and12623(N21090,N21092,N21093);
and and12624(N21091,N21094,N21095);
and and12631(N21104,N21106,N21107);
and and12632(N21105,N21108,N21109);
and and12639(N21118,N21120,N21121);
and and12640(N21119,N21122,N21123);
and and12647(N21132,N21134,N21135);
and and12648(N21133,N21136,N21137);
and and12655(N21146,N21148,N21149);
and and12656(N21147,N21150,N21151);
and and12663(N21160,N21162,N21163);
and and12664(N21161,N21164,N21165);
and and12671(N21174,N21176,N21177);
and and12672(N21175,N21178,N21179);
and and12679(N21188,N21190,N21191);
and and12680(N21189,N21192,N21193);
and and12687(N21202,N21204,N21205);
and and12688(N21203,N21206,N21207);
and and12695(N21216,N21218,N21219);
and and12696(N21217,N21220,N21221);
and and12703(N21230,N21232,N21233);
and and12704(N21231,N21234,N21235);
and and12711(N21244,N21246,N21247);
and and12712(N21245,N21248,N21249);
and and12719(N21258,N21260,N21261);
and and12720(N21259,N21262,N21263);
and and12727(N21272,N21274,N21275);
and and12728(N21273,N21276,N21277);
and and12735(N21286,N21288,N21289);
and and12736(N21287,N21290,N21291);
and and12743(N21300,N21302,N21303);
and and12744(N21301,N21304,N21305);
and and12751(N21314,N21316,N21317);
and and12752(N21315,N21318,N21319);
and and12759(N21328,N21330,N21331);
and and12760(N21329,N21332,N21333);
and and12767(N21342,N21344,N21345);
and and12768(N21343,N21346,N21347);
and and12775(N21356,N21358,N21359);
and and12776(N21357,N21360,N21361);
and and12783(N21370,N21372,N21373);
and and12784(N21371,N21374,N21375);
and and12791(N21384,N21386,N21387);
and and12792(N21385,N21388,N21389);
and and12799(N21398,N21400,N21401);
and and12800(N21399,N21402,N21403);
and and12807(N21412,N21414,N21415);
and and12808(N21413,N21416,N21417);
and and12815(N21426,N21428,N21429);
and and12816(N21427,N21430,N21431);
and and12823(N21440,N21442,N21443);
and and12824(N21441,N21444,N21445);
and and12831(N21454,N21456,N21457);
and and12832(N21455,N21458,N21459);
and and12839(N21468,N21470,N21471);
and and12840(N21469,N21472,N21473);
and and12847(N21482,N21484,N21485);
and and12848(N21483,N21486,N21487);
and and12855(N21496,N21498,N21499);
and and12856(N21497,N21500,N21501);
and and12863(N21510,N21512,N21513);
and and12864(N21511,N21514,N21515);
and and12871(N21524,N21526,N21527);
and and12872(N21525,N21528,N21529);
and and12879(N21537,N21539,N21540);
and and12880(N21538,N21541,N21542);
and and12887(N21550,N21552,N21553);
and and12888(N21551,N21554,N21555);
and and12895(N21563,N21565,N21566);
and and12896(N21564,N21567,N21568);
and and12903(N21576,N21578,N21579);
and and12904(N21577,N21580,N21581);
and and12911(N21589,N21591,N21592);
and and12912(N21590,N21593,N21594);
and and12919(N21602,N21604,N21605);
and and12920(N21603,N21606,N21607);
and and12927(N21615,N21617,N21618);
and and12928(N21616,N21619,N21620);
and and12935(N21628,N21630,N21631);
and and12936(N21629,N21632,N21633);
and and12943(N21641,N21643,N21644);
and and12944(N21642,N21645,N21646);
and and12951(N21654,N21656,N21657);
and and12952(N21655,N21658,N21659);
and and12959(N21667,N21669,N21670);
and and12960(N21668,N21671,N21672);
and and12967(N21680,N21682,N21683);
and and12968(N21681,N21684,N21685);
and and12975(N21693,N21695,N21696);
and and12976(N21694,N21697,N21698);
and and12983(N21706,N21708,N21709);
and and12984(N21707,N21710,N21711);
and and12991(N21719,N21721,N21722);
and and12992(N21720,N21723,N21724);
and and12999(N21732,N21734,N21735);
and and13000(N21733,N21736,N21737);
and and13007(N21745,N21747,N21748);
and and13008(N21746,N21749,N21750);
and and13015(N21758,N21760,N21761);
and and13016(N21759,N21762,N21763);
and and13023(N21771,N21773,N21774);
and and13024(N21772,N21775,N21776);
and and13031(N21784,N21786,N21787);
and and13032(N21785,N21788,N21789);
and and13039(N21797,N21799,N21800);
and and13040(N21798,N21801,N21802);
and and13047(N21810,N21812,N21813);
and and13048(N21811,N21814,N21815);
and and13055(N21823,N21825,N21826);
and and13056(N21824,N21827,N21828);
and and13063(N21836,N21838,N21839);
and and13064(N21837,N21840,N21841);
and and13071(N21849,N21851,N21852);
and and13072(N21850,N21853,N21854);
and and13079(N21862,N21864,N21865);
and and13080(N21863,N21866,N21867);
and and13087(N21875,N21877,N21878);
and and13088(N21876,N21879,N21880);
and and13095(N21888,N21890,N21891);
and and13096(N21889,N21892,N21893);
and and13103(N21901,N21903,N21904);
and and13104(N21902,N21905,N21906);
and and13111(N21914,N21916,N21917);
and and13112(N21915,N21918,N21919);
and and13119(N21927,N21929,N21930);
and and13120(N21928,N21931,N21932);
and and13127(N21940,N21942,N21943);
and and13128(N21941,N21944,N21945);
and and13135(N21953,N21955,N21956);
and and13136(N21954,N21957,N21958);
and and13143(N21966,N21968,N21969);
and and13144(N21967,N21970,N21971);
and and13151(N21979,N21981,N21982);
and and13152(N21980,N21983,N21984);
and and13159(N21992,N21994,N21995);
and and13160(N21993,N21996,N21997);
and and13167(N22005,N22007,N22008);
and and13168(N22006,N22009,N22010);
and and13175(N22018,N22020,N22021);
and and13176(N22019,N22022,N22023);
and and13183(N22031,N22033,N22034);
and and13184(N22032,N22035,N22036);
and and13191(N22044,N22046,N22047);
and and13192(N22045,N22048,N22049);
and and13199(N22057,N22059,N22060);
and and13200(N22058,N22061,N22062);
and and13207(N22070,N22072,N22073);
and and13208(N22071,N22074,N22075);
and and13215(N22083,N22085,N22086);
and and13216(N22084,N22087,N22088);
and and13223(N22096,N22098,N22099);
and and13224(N22097,N22100,N22101);
and and13231(N22109,N22111,N22112);
and and13232(N22110,N22113,N22114);
and and13239(N22122,N22124,N22125);
and and13240(N22123,N22126,N22127);
and and13247(N22135,N22137,N22138);
and and13248(N22136,N22139,N22140);
and and13255(N22148,N22150,N22151);
and and13256(N22149,N22152,N22153);
and and13263(N22161,N22163,N22164);
and and13264(N22162,N22165,N22166);
and and13271(N22174,N22176,N22177);
and and13272(N22175,N22178,N22179);
and and13279(N22187,N22189,N22190);
and and13280(N22188,N22191,N22192);
and and13287(N22200,N22202,N22203);
and and13288(N22201,N22204,N22205);
and and13295(N22213,N22215,N22216);
and and13296(N22214,N22217,N22218);
and and13303(N22226,N22228,N22229);
and and13304(N22227,N22230,N22231);
and and13311(N22238,N22240,N22241);
and and13312(N22239,N22242,N22243);
and and13319(N22250,N22252,N22253);
and and13320(N22251,N22254,N22255);
and and13327(N22262,N22264,N22265);
and and13328(N22263,N22266,N22267);
and and13335(N22274,N22276,N22277);
and and13336(N22275,N22278,N22279);
and and13343(N22286,N22288,N22289);
and and13344(N22287,N22290,N22291);
and and13351(N22298,N22300,N22301);
and and13352(N22299,N22302,N22303);
and and13359(N22310,N22312,N22313);
and and13360(N22311,N22314,N22315);
and and13367(N22322,N22324,N22325);
and and13368(N22323,N22326,N22327);
and and13375(N22334,N22336,N22337);
and and13376(N22335,N22338,N22339);
and and13383(N22346,N22348,N22349);
and and13384(N22347,N22350,N22351);
and and13391(N22358,N22360,N22361);
and and13392(N22359,N22362,N22363);
and and13399(N22370,N22372,N22373);
and and13400(N22371,N22374,N22375);
and and13407(N22382,N22384,N22385);
and and13408(N22383,N22386,N22387);
and and13415(N22394,N22396,N22397);
and and13416(N22395,N22398,N22399);
and and13423(N22406,N22408,N22409);
and and13424(N22407,N22410,N22411);
and and13431(N22418,N22420,N22421);
and and13432(N22419,N22422,N22423);
and and13439(N22430,N22432,N22433);
and and13440(N22431,N22434,N22435);
and and13447(N22442,N22444,N22445);
and and13448(N22443,N22446,N22447);
and and13455(N22454,N22456,N22457);
and and13456(N22455,N22458,N22459);
and and13463(N22466,N22468,N22469);
and and13464(N22467,N22470,N22471);
and and13471(N22478,N22480,N22481);
and and13472(N22479,N22482,N22483);
and and13479(N22490,N22492,N22493);
and and13480(N22491,N22494,N22495);
and and13487(N22502,N22504,N22505);
and and13488(N22503,N22506,N22507);
and and13495(N22514,N22516,N22517);
and and13496(N22515,N22518,N22519);
and and13503(N22526,N22528,N22529);
and and13504(N22527,N22530,N22531);
and and13511(N22538,N22540,N22541);
and and13512(N22539,N22542,N22543);
and and13519(N22550,N22552,N22553);
and and13520(N22551,N22554,N22555);
and and13527(N22562,N22564,N22565);
and and13528(N22563,N22566,N22567);
and and13535(N22574,N22576,N22577);
and and13536(N22575,N22578,N22579);
and and13543(N22586,N22588,N22589);
and and13544(N22587,N22590,N22591);
and and13551(N22598,N22600,N22601);
and and13552(N22599,N22602,N22603);
and and13559(N22610,N22612,N22613);
and and13560(N22611,N22614,N22615);
and and13567(N22622,N22624,N22625);
and and13568(N22623,N22626,N22627);
and and13575(N22634,N22636,N22637);
and and13576(N22635,N22638,N22639);
and and13583(N22646,N22648,N22649);
and and13584(N22647,N22650,N22651);
and and13591(N22658,N22660,N22661);
and and13592(N22659,N22662,N22663);
and and13599(N22670,N22672,N22673);
and and13600(N22671,N22674,N22675);
and and13607(N22682,N22684,N22685);
and and13608(N22683,N22686,N22687);
and and13615(N22694,N22696,N22697);
and and13616(N22695,N22698,N22699);
and and13623(N22706,N22708,N22709);
and and13624(N22707,N22710,N22711);
and and13631(N22718,N22720,N22721);
and and13632(N22719,N22722,N22723);
and and13639(N22730,N22732,N22733);
and and13640(N22731,N22734,N22735);
and and13647(N22742,N22744,N22745);
and and13648(N22743,N22746,N22747);
and and13655(N22754,N22756,N22757);
and and13656(N22755,N22758,N22759);
and and13663(N22766,N22768,N22769);
and and13664(N22767,N22770,N22771);
and and13671(N22778,N22780,N22781);
and and13672(N22779,N22782,N22783);
and and13679(N22790,N22792,N22793);
and and13680(N22791,N22794,N22795);
and and13687(N22802,N22804,N22805);
and and13688(N22803,N22806,N22807);
and and13695(N22814,N22816,N22817);
and and13696(N22815,N22818,N22819);
and and13703(N22826,N22828,N22829);
and and13704(N22827,N22830,N22831);
and and13711(N22837,N22839,N22840);
and and13712(N22838,N22841,N22842);
and and13719(N22848,N22850,N22851);
and and13720(N22849,N22852,N22853);
and and13727(N22859,N22861,N22862);
and and13728(N22860,N22863,N22864);
and and13735(N22870,N22872,N22873);
and and13736(N22871,N22874,N22875);
and and13743(N22881,N22883,N22884);
and and13744(N22882,N22885,N22886);
and and13751(N22892,N22894,N22895);
and and13752(N22893,N22896,N22897);
and and13759(N22903,N22905,N22906);
and and13760(N22904,N22907,N22908);
and and13767(N22914,N22916,N22917);
and and13768(N22915,N22918,N22919);
and and13775(N22925,N22927,N22928);
and and13776(N22926,N22929,N22930);
and and13783(N22936,N22938,N22939);
and and13784(N22937,N22940,N22941);
and and13791(N22947,N22949,N22950);
and and13792(N22948,N22951,N22952);
and and13799(N22958,N22960,N22961);
and and13800(N22959,N22962,N22963);
and and13807(N22969,N22971,N22972);
and and13808(N22970,N22973,N22974);
and and13815(N22980,N22982,N22983);
and and13816(N22981,N22984,N22985);
and and13823(N22991,N22993,N22994);
and and13824(N22992,N22995,N22996);
and and13831(N23002,N23004,N23005);
and and13832(N23003,N23006,N23007);
and and13839(N23013,N23015,N23016);
and and13840(N23014,N23017,N23018);
and and13847(N23024,N23026,N23027);
and and13848(N23025,N23028,N23029);
and and13855(N23035,N23037,N23038);
and and13856(N23036,N23039,N23040);
and and13863(N23046,N23048,N23049);
and and13864(N23047,N23050,N23051);
and and13871(N23057,N23059,N23060);
and and13872(N23058,N23061,N23062);
and and13879(N23068,N23070,N23071);
and and13880(N23069,N23072,N23073);
and and13887(N23079,N23081,N23082);
and and13888(N23080,N23083,N23084);
and and13895(N23090,N23092,N23093);
and and13896(N23091,N23094,N23095);
and and13903(N23101,N23103,N23104);
and and13904(N23102,N23105,N23106);
and and13911(N23112,N23114,N23115);
and and13912(N23113,N23116,N23117);
and and13919(N23123,N23125,N23126);
and and13920(N23124,N23127,N23128);
and and13927(N23134,N23136,N23137);
and and13928(N23135,N23138,N23139);
and and13935(N23145,N23147,N23148);
and and13936(N23146,N23149,N23150);
and and13943(N23156,N23158,N23159);
and and13944(N23157,N23160,N23161);
and and13951(N23167,N23169,N23170);
and and13952(N23168,N23171,N23172);
and and13959(N23178,N23180,N23181);
and and13960(N23179,N23182,N23183);
and and13967(N23189,N23191,N23192);
and and13968(N23190,N23193,N23194);
and and13975(N23200,N23202,N23203);
and and13976(N23201,N23204,N23205);
and and13983(N23211,N23213,N23214);
and and13984(N23212,N23215,N23216);
and and13991(N23222,N23224,N23225);
and and13992(N23223,N23226,N23227);
and and13999(N23233,N23235,N23236);
and and14000(N23234,N23237,N23238);
and and14007(N23244,N23246,N23247);
and and14008(N23245,N23248,N23249);
and and14015(N23255,N23257,N23258);
and and14016(N23256,N23259,N23260);
and and14023(N23266,N23268,N23269);
and and14024(N23267,N23270,N23271);
and and14031(N23277,N23279,N23280);
and and14032(N23278,N23281,N23282);
and and14039(N23288,N23290,N23291);
and and14040(N23289,N23292,N23293);
and and14047(N23299,N23301,N23302);
and and14048(N23300,N23303,N23304);
and and14055(N23310,N23312,N23313);
and and14056(N23311,N23314,N23315);
and and14063(N23321,N23323,N23324);
and and14064(N23322,N23325,N23326);
and and14071(N23332,N23334,N23335);
and and14072(N23333,N23336,N23337);
and and14079(N23343,N23345,N23346);
and and14080(N23344,N23347,N23348);
and and14087(N23354,N23356,N23357);
and and14088(N23355,N23358,N23359);
and and14095(N23365,N23367,N23368);
and and14096(N23366,N23369,N23370);
and and14103(N23376,N23378,N23379);
and and14104(N23377,N23380,N23381);
and and14111(N23387,N23389,N23390);
and and14112(N23388,N23391,N23392);
and and14119(N23398,N23400,N23401);
and and14120(N23399,N23402,N23403);
and and14127(N23408,N23410,N23411);
and and14128(N23409,N23412,N23413);
and and14135(N23418,N23420,N23421);
and and14136(N23419,N23422,N23423);
and and14143(N23428,N23430,N23431);
and and14144(N23429,N23432,N23433);
and and14151(N23438,N23440,N23441);
and and14152(N23439,N23442,N23443);
and and14159(N23448,N23450,N23451);
and and14160(N23449,N23452,N23453);
and and14167(N23458,N23460,N23461);
and and14168(N23459,N23462,N23463);
and and14175(N23468,N23470,N23471);
and and14176(N23469,N23472,N23473);
and and14183(N23478,N23480,N23481);
and and14184(N23479,N23482,N23483);
and and14191(N23488,N23490,N23491);
and and14192(N23489,N23492,N23493);
and and14199(N23498,N23500,N23501);
and and14200(N23499,N23502,N23503);
and and14207(N23508,N23510,N23511);
and and14208(N23509,N23512,N23513);
and and14215(N23518,N23520,N23521);
and and14216(N23519,N23522,N23523);
and and14223(N23528,N23530,N23531);
and and14224(N23529,N23532,N23533);
and and14231(N23538,N23540,N23541);
and and14232(N23539,N23542,N23543);
and and14239(N23548,N23550,N23551);
and and14240(N23549,N23552,N23553);
and and14247(N23557,N23559,N23560);
and and14248(N23558,N23561,N23562);
and and14255(N23566,N23568,N23569);
and and14256(N23567,N23570,N23571);
and and14263(N23575,N23577,N23578);
and and14264(N23576,N23579,N23580);
and and14271(N23584,N23586,N23587);
and and14272(N23585,N23588,N23589);
and and14279(N23593,N23595,N23596);
and and14280(N23594,N23597,N23598);
and and14287(N23602,N23604,N23605);
and and14288(N23603,N23606,N23607);
and and14295(N23611,N23613,N23614);
and and14296(N23612,N23615,N23616);
and and14303(N23620,N23622,N23623);
and and14304(N23621,N23624,N23625);
and and14311(N23629,N23631,N23632);
and and14312(N23630,N23633,N23634);
and and14319(N23637,N23639,N23640);
and and14320(N23638,N23641,N23642);
and and14326(N23651,N23653,N23654);
and and14327(N23652,N23655,N23656);
and and14333(N23665,N23667,N23668);
and and14334(N23666,N23669,N23670);
and and14340(N23678,N23680,N23681);
and and14341(N23679,N23682,N23683);
and and14347(N23691,N23693,N23694);
and and14348(N23692,N23695,N23696);
and and14354(N23704,N23706,N23707);
and and14355(N23705,N23708,N23709);
and and14361(N23717,N23719,N23720);
and and14362(N23718,N23721,N23722);
and and14368(N23730,N23732,N23733);
and and14369(N23731,N23734,N23735);
and and14375(N23743,N23745,N23746);
and and14376(N23744,N23747,N23748);
and and14382(N23755,N23757,N23758);
and and14383(N23756,N23759,N23760);
and and14389(N23767,N23769,N23770);
and and14390(N23768,N23771,N23772);
and and14396(N23779,N23781,N23782);
and and14397(N23780,N23783,N23784);
and and14403(N23791,N23793,N23794);
and and14404(N23792,N23795,N23796);
and and14410(N23803,N23805,N23806);
and and14411(N23804,N23807,N23808);
and and14417(N23815,N23817,N23818);
and and14418(N23816,N23819,N23820);
and and14424(N23827,N23829,N23830);
and and14425(N23828,N23831,N23832);
and and14431(N23839,N23841,N23842);
and and14432(N23840,N23843,N23844);
and and14438(N23851,N23853,N23854);
and and14439(N23852,N23855,N23856);
and and14445(N23862,N23864,N23865);
and and14446(N23863,N23866,N23867);
and and14452(N23873,N23875,N23876);
and and14453(N23874,N23877,N23878);
and and14459(N23884,N23886,N23887);
and and14460(N23885,N23888,N23889);
and and14466(N23895,N23897,N23898);
and and14467(N23896,N23899,N23900);
and and14473(N23906,N23908,N23909);
and and14474(N23907,N23910,N23911);
and and14480(N23917,N23919,N23920);
and and14481(N23918,N23921,N23922);
and and14487(N23928,N23930,N23931);
and and14488(N23929,N23932,N23933);
and and14494(N23939,N23941,N23942);
and and14495(N23940,N23943,N23944);
and and14501(N23949,N23951,N23952);
and and14502(N23950,N23953,N23954);
and and14508(N23959,N23961,N23962);
and and14509(N23960,N23963,N23964);
and and14515(N23969,N23971,N23972);
and and14516(N23970,N23973,N23974);
and and14522(N23979,N23981,N23982);
and and14523(N23980,N23983,N23984);
and and14529(N23989,N23991,N23992);
and and14530(N23990,N23993,N23994);
and and14536(N23999,N24001,N24002);
and and14537(N24000,N24003,N24004);
and and14543(N24009,N24011,N24012);
and and14544(N24010,N24013,N24014);
and and14550(N24019,N24021,N24022);
and and14551(N24020,N24023,N24024);
and and14557(N24029,N24031,N24032);
and and14558(N24030,N24033,N24034);
and and14564(N24039,N24041,N24042);
and and14565(N24040,N24043,N24044);
and and14571(N24048,N24050,N24051);
and and14572(N24049,N24052,N24053);
and and10679(N18113,N18117,N18118);
and and10680(N18114,N18119,N18120);
and and10681(N18115,N18121,R1);
and and10682(N18116,N18122,N18123);
and and10688(N18131,N18135,N18136);
and and10689(N18132,N18137,N18138);
and and10690(N18133,R0,N18139);
and and10691(N18134,N18140,N18141);
and and10697(N18148,N18152,N18153);
and and10698(N18149,N18154,in2);
and and10699(N18150,N18155,N18156);
and and10700(N18151,N18157,N18158);
and and10706(N18165,N18169,N18170);
and and10707(N18166,N18171,N18172);
and and10708(N18167,N18173,N18174);
and and10709(N18168,R2,N18175);
and and10715(N18182,N18186,N18187);
and and10716(N18183,N18188,in2);
and and10717(N18184,N18189,N18190);
and and10718(N18185,N18191,N18192);
and and10724(N18199,N18203,N18204);
and and10725(N18200,N18205,N18206);
and and10726(N18201,N18207,N18208);
and and10727(N18202,N18209,N18210);
and and10733(N18216,N18220,N18221);
and and10734(N18217,N18222,N18223);
and and10735(N18218,N18224,R0);
and and10736(N18219,N18225,N18226);
and and10742(N18233,N18237,N18238);
and and10743(N18234,N18239,in2);
and and10744(N18235,N18240,R1);
and and10745(N18236,N18241,R3);
and and10751(N18249,N18253,N18254);
and and10752(N18250,N18255,in2);
and and10753(N18251,N18256,N18257);
and and10754(N18252,N18258,N18259);
and and10760(N18265,N18269,N18270);
and and10761(N18266,N18271,in2);
and and10762(N18267,N18272,N18273);
and and10763(N18268,N18274,R3);
and and10769(N18281,N18285,N18286);
and and10770(N18282,in1,N18287);
and and10771(N18283,N18288,N18289);
and and10772(N18284,R2,N18290);
and and10778(N18297,N18301,N18302);
and and10779(N18298,N18303,in2);
and and10780(N18299,N18304,N18305);
and and10781(N18300,R2,N18306);
and and10787(N18313,N18317,N18318);
and and10788(N18314,N18319,N18320);
and and10789(N18315,N18321,R1);
and and10790(N18316,N18322,R3);
and and10796(N18329,N18333,N18334);
and and10797(N18330,N18335,N18336);
and and10798(N18331,N18337,R0);
and and10799(N18332,R1,N18338);
and and10805(N18345,N18349,N18350);
and and10806(N18346,N18351,N18352);
and and10807(N18347,N18353,N18354);
and and10808(N18348,R1,R2);
and and10814(N18361,N18365,N18366);
and and10815(N18362,N18367,N18368);
and and10816(N18363,N18369,N18370);
and and10817(N18364,R1,N18371);
and and10823(N18377,N18381,N18382);
and and10824(N18378,N18383,in1);
and and10825(N18379,N18384,R1);
and and10826(N18380,N18385,N18386);
and and10832(N18393,N18397,N18398);
and and10833(N18394,N18399,N18400);
and and10834(N18395,in2,R0);
and and10835(N18396,N18401,R2);
and and10841(N18409,N18413,N18414);
and and10842(N18410,N18415,in1);
and and10843(N18411,R0,N18416);
and and10844(N18412,R2,N18417);
and and10850(N18425,N18429,N18430);
and and10851(N18426,N18431,N18432);
and and10852(N18427,N18433,R0);
and and10853(N18428,N18434,R2);
and and10859(N18441,N18445,N18446);
and and10860(N18442,N18447,in1);
and and10861(N18443,N18448,R1);
and and10862(N18444,N18449,N18450);
and and10868(N18457,N18461,N18462);
and and10869(N18458,N18463,in2);
and and10870(N18459,N18464,N18465);
and and10871(N18460,N18466,R3);
and and10877(N18473,N18477,N18478);
and and10878(N18474,N18479,N18480);
and and10879(N18475,in2,R0);
and and10880(N18476,N18481,N18482);
and and10886(N18489,N18493,N18494);
and and10887(N18490,N18495,in1);
and and10888(N18491,N18496,R0);
and and10889(N18492,N18497,N18498);
and and10895(N18505,N18509,N18510);
and and10896(N18506,in0,N18511);
and and10897(N18507,N18512,N18513);
and and10898(N18508,R1,N18514);
and and10904(N18521,N18525,N18526);
and and10905(N18522,N18527,N18528);
and and10906(N18523,in2,N18529);
and and10907(N18524,R1,N18530);
and and10913(N18537,N18541,N18542);
and and10914(N18538,N18543,N18544);
and and10915(N18539,N18545,N18546);
and and10916(N18540,R2,N18547);
and and10922(N18553,N18557,N18558);
and and10923(N18554,N18559,N18560);
and and10924(N18555,R0,R1);
and and10925(N18556,N18561,N18562);
and and10931(N18568,N18572,N18573);
and and10932(N18569,N18574,N18575);
and and10933(N18570,in2,R0);
and and10934(N18571,R1,R3);
and and10940(N18583,N18587,N18588);
and and10941(N18584,N18589,N18590);
and and10942(N18585,R0,N18591);
and and10943(N18586,R2,R3);
and and10949(N18598,N18602,N18603);
and and10950(N18599,N18604,in2);
and and10951(N18600,R0,R1);
and and10952(N18601,R2,N18605);
and and10958(N18613,N18617,N18618);
and and10959(N18614,N18619,N18620);
and and10960(N18615,N18621,R1);
and and10961(N18616,N18622,R3);
and and10967(N18628,N18632,N18633);
and and10968(N18629,in0,N18634);
and and10969(N18630,N18635,N18636);
and and10970(N18631,R2,R3);
and and10976(N18643,N18647,N18648);
and and10977(N18644,N18649,in2);
and and10978(N18645,R0,R1);
and and10979(N18646,N18650,N18651);
and and10985(N18658,N18662,N18663);
and and10986(N18659,in0,N18664);
and and10987(N18660,R0,R1);
and and10988(N18661,N18665,N18666);
and and10994(N18673,N18677,N18678);
and and10995(N18674,N18679,N18680);
and and10996(N18675,N18681,N18682);
and and10997(N18676,R2,R3);
and and11003(N18688,N18692,N18693);
and and11004(N18689,N18694,N18695);
and and11005(N18690,in2,N18696);
and and11006(N18691,R1,R2);
and and11012(N18703,N18707,N18708);
and and11013(N18704,N18709,N18710);
and and11014(N18705,N18711,R1);
and and11015(N18706,R2,N18712);
and and11021(N18718,N18722,N18723);
and and11022(N18719,in0,N18724);
and and11023(N18720,N18725,N18726);
and and11024(N18721,N18727,R3);
and and11030(N18733,N18737,N18738);
and and11031(N18734,N18739,in1);
and and11032(N18735,in2,R0);
and and11033(N18736,R1,N18740);
and and11039(N18748,N18752,N18753);
and and11040(N18749,in0,in1);
and and11041(N18750,N18754,R0);
and and11042(N18751,R1,N18755);
and and11048(N18763,N18767,N18768);
and and11049(N18764,in0,in1);
and and11050(N18765,N18769,R0);
and and11051(N18766,N18770,R2);
and and11057(N18778,N18782,N18783);
and and11058(N18779,N18784,in2);
and and11059(N18780,N18785,N18786);
and and11060(N18781,N18787,R3);
and and11066(N18793,N18797,N18798);
and and11067(N18794,in0,N18799);
and and11068(N18795,N18800,N18801);
and and11069(N18796,N18802,R3);
and and11075(N18808,N18812,N18813);
and and11076(N18809,N18814,in2);
and and11077(N18810,N18815,R1);
and and11078(N18811,N18816,N18817);
and and11084(N18823,N18827,N18828);
and and11085(N18824,in1,in2);
and and11086(N18825,N18829,R1);
and and11087(N18826,N18830,N18831);
and and11093(N18838,N18842,N18843);
and and11094(N18839,N18844,N18845);
and and11095(N18840,R0,N18846);
and and11096(N18841,R2,R3);
and and11102(N18853,N18857,N18858);
and and11103(N18854,N18859,N18860);
and and11104(N18855,N18861,R0);
and and11105(N18856,R1,N18862);
and and11111(N18868,N18872,N18873);
and and11112(N18869,N18874,in2);
and and11113(N18870,R0,R1);
and and11114(N18871,N18875,N18876);
and and11120(N18883,N18887,N18888);
and and11121(N18884,N18889,N18890);
and and11122(N18885,N18891,R0);
and and11123(N18886,R1,R2);
and and11129(N18898,N18902,N18903);
and and11130(N18899,N18904,N18905);
and and11131(N18900,R0,R1);
and and11132(N18901,N18906,N18907);
and and11138(N18913,N18917,N18918);
and and11139(N18914,in0,N18919);
and and11140(N18915,in2,N18920);
and and11141(N18916,R2,R3);
and and11147(N18927,N18931,N18932);
and and11148(N18928,in1,N18933);
and and11149(N18929,R0,R1);
and and11150(N18930,R2,N18934);
and and11156(N18941,N18945,N18946);
and and11157(N18942,in1,in2);
and and11158(N18943,R0,N18947);
and and11159(N18944,R2,N18948);
and and11165(N18955,N18959,N18960);
and and11166(N18956,in0,in2);
and and11167(N18957,R0,N18961);
and and11168(N18958,N18962,R3);
and and11174(N18969,N18973,N18974);
and and11175(N18970,N18975,N18976);
and and11176(N18971,in2,R0);
and and11177(N18972,R2,R3);
and and11183(N18983,N18987,N18988);
and and11184(N18984,in1,N18989);
and and11185(N18985,N18990,R1);
and and11186(N18986,N18991,R3);
and and11192(N18997,N19001,N19002);
and and11193(N18998,N19003,in2);
and and11194(N18999,N19004,R1);
and and11195(N19000,N19005,R3);
and and11201(N19011,N19015,N19016);
and and11202(N19012,in0,in2);
and and11203(N19013,N19017,R1);
and and11204(N19014,N19018,R3);
and and11210(N19025,N19029,N19030);
and and11211(N19026,in0,in1);
and and11212(N19027,N19031,N19032);
and and11213(N19028,R1,N19033);
and and11219(N19039,N19043,N19044);
and and11220(N19040,N19045,in1);
and and11221(N19041,R0,R1);
and and11222(N19042,N19046,N19047);
and and11228(N19053,N19057,N19058);
and and11229(N19054,in0,N19059);
and and11230(N19055,R0,R1);
and and11231(N19056,N19060,N19061);
and and11237(N19067,N19071,N19072);
and and11238(N19068,in1,N19073);
and and11239(N19069,N19074,R1);
and and11240(N19070,R2,N19075);
and and11246(N19081,N19085,N19086);
and and11247(N19082,N19087,in1);
and and11248(N19083,in2,N19088);
and and11249(N19084,N19089,R3);
and and11255(N19095,N19099,N19100);
and and11256(N19096,N19101,N19102);
and and11257(N19097,N19103,R0);
and and11258(N19098,R1,N19104);
and and11264(N19109,N19113,N19114);
and and11265(N19110,N19115,N19116);
and and11266(N19111,in2,R0);
and and11267(N19112,N19117,R3);
and and11273(N19123,N19127,N19128);
and and11274(N19124,in0,in1);
and and11275(N19125,N19129,N19130);
and and11276(N19126,R2,N19131);
and and11282(N19137,N19141,N19142);
and and11283(N19138,in1,N19143);
and and11284(N19139,N19144,R1);
and and11285(N19140,R2,N19145);
and and11291(N19151,N19155,N19156);
and and11292(N19152,N19157,N19158);
and and11293(N19153,R0,N19159);
and and11294(N19154,R2,N19160);
and and11300(N19165,N19169,N19170);
and and11301(N19166,in0,in2);
and and11302(N19167,N19171,N19172);
and and11303(N19168,R2,R3);
and and11309(N19179,N19183,N19184);
and and11310(N19180,N19185,in1);
and and11311(N19181,in2,N19186);
and and11312(N19182,R2,R3);
and and11318(N19193,N19197,N19198);
and and11319(N19194,in0,N19199);
and and11320(N19195,in2,R1);
and and11321(N19196,R2,N19200);
and and11327(N19207,N19211,N19212);
and and11328(N19208,in0,N19213);
and and11329(N19209,N19214,R1);
and and11330(N19210,N19215,N19216);
and and11336(N19221,N19225,N19226);
and and11337(N19222,in0,in2);
and and11338(N19223,N19227,N19228);
and and11339(N19224,N19229,R3);
and and11345(N19235,N19239,N19240);
and and11346(N19236,in0,in1);
and and11347(N19237,N19241,N19242);
and and11348(N19238,N19243,R3);
and and11354(N19249,N19253,N19254);
and and11355(N19250,N19255,in1);
and and11356(N19251,N19256,R0);
and and11357(N19252,N19257,R2);
and and11363(N19263,N19267,N19268);
and and11364(N19264,N19269,in2);
and and11365(N19265,N19270,R1);
and and11366(N19266,N19271,R3);
and and11372(N19277,N19281,N19282);
and and11373(N19278,in0,N19283);
and and11374(N19279,N19284,N19285);
and and11375(N19280,R1,R3);
and and11381(N19291,N19295,N19296);
and and11382(N19292,in1,N19297);
and and11383(N19293,N19298,R1);
and and11384(N19294,N19299,R3);
and and11390(N19305,N19309,N19310);
and and11391(N19306,in1,N19311);
and and11392(N19307,N19312,N19313);
and and11393(N19308,R2,N19314);
and and11399(N19319,N19323,N19324);
and and11400(N19320,in0,in1);
and and11401(N19321,N19325,N19326);
and and11402(N19322,N19327,R2);
and and11408(N19333,N19337,N19338);
and and11409(N19334,in0,in2);
and and11410(N19335,R0,N19339);
and and11411(N19336,N19340,N19341);
and and11417(N19347,N19351,N19352);
and and11418(N19348,in0,N19353);
and and11419(N19349,in2,R0);
and and11420(N19350,N19354,N19355);
and and11426(N19361,N19365,N19366);
and and11427(N19362,N19367,in1);
and and11428(N19363,in2,R0);
and and11429(N19364,R2,N19368);
and and11435(N19375,N19379,N19380);
and and11436(N19376,in0,in1);
and and11437(N19377,in2,N19381);
and and11438(N19378,N19382,N19383);
and and11444(N19389,N19393,N19394);
and and11445(N19390,N19395,N19396);
and and11446(N19391,N19397,R0);
and and11447(N19392,R2,R3);
and and11453(N19403,N19407,N19408);
and and11454(N19404,N19409,N19410);
and and11455(N19405,N19411,R0);
and and11456(N19406,R2,N19412);
and and11462(N19417,N19421,N19422);
and and11463(N19418,in0,N19423);
and and11464(N19419,N19424,N19425);
and and11465(N19420,R2,N19426);
and and11471(N19431,N19435,N19436);
and and11472(N19432,N19437,in1);
and and11473(N19433,N19438,N19439);
and and11474(N19434,N19440,R2);
and and11480(N19445,N19449,N19450);
and and11481(N19446,N19451,in1);
and and11482(N19447,in2,N19452);
and and11483(N19448,R1,R2);
and and11489(N19459,N19463,N19464);
and and11490(N19460,N19465,in1);
and and11491(N19461,in2,N19466);
and and11492(N19462,R2,R3);
and and11498(N19473,N19477,N19478);
and and11499(N19474,in0,N19479);
and and11500(N19475,N19480,R0);
and and11501(N19476,R1,N19481);
and and11507(N19487,N19491,N19492);
and and11508(N19488,in1,N19493);
and and11509(N19489,R0,R1);
and and11510(N19490,N19494,R3);
and and11516(N19501,N19505,N19506);
and and11517(N19502,N19507,in1);
and and11518(N19503,N19508,R0);
and and11519(N19504,N19509,R2);
and and11525(N19515,N19519,N19520);
and and11526(N19516,in0,N19521);
and and11527(N19517,N19522,R0);
and and11528(N19518,N19523,R2);
and and11534(N19529,N19533,N19534);
and and11535(N19530,N19535,N19536);
and and11536(N19531,in2,R0);
and and11537(N19532,N19537,R2);
and and11543(N19543,N19547,N19548);
and and11544(N19544,N19549,N19550);
and and11545(N19545,in2,N19551);
and and11546(N19546,R2,R3);
and and11552(N19557,N19561,N19562);
and and11553(N19558,N19563,in1);
and and11554(N19559,N19564,R0);
and and11555(N19560,N19565,N19566);
and and11561(N19571,N19575,N19576);
and and11562(N19572,N19577,N19578);
and and11563(N19573,in2,R0);
and and11564(N19574,N19579,R3);
and and11570(N19585,N19589,N19590);
and and11571(N19586,N19591,N19592);
and and11572(N19587,in2,R0);
and and11573(N19588,R1,R2);
and and11579(N19599,N19603,N19604);
and and11580(N19600,N19605,N19606);
and and11581(N19601,R0,R1);
and and11582(N19602,N19607,R3);
and and11588(N19613,N19617,N19618);
and and11589(N19614,N19619,N19620);
and and11590(N19615,N19621,N19622);
and and11591(N19616,R1,R2);
and and11597(N19627,N19631,N19632);
and and11598(N19628,in0,in1);
and and11599(N19629,N19633,N19634);
and and11600(N19630,N19635,R2);
and and11606(N19641,N19645,N19646);
and and11607(N19642,N19647,in1);
and and11608(N19643,in2,N19648);
and and11609(N19644,R1,R2);
and and11615(N19655,N19659,N19660);
and and11616(N19656,in0,in1);
and and11617(N19657,N19661,R1);
and and11618(N19658,R2,N19662);
and and11624(N19669,N19673,N19674);
and and11625(N19670,in0,N19675);
and and11626(N19671,N19676,R0);
and and11627(N19672,N19677,N19678);
and and11633(N19683,N19687,N19688);
and and11634(N19684,in0,N19689);
and and11635(N19685,N19690,N19691);
and and11636(N19686,R2,R3);
and and11642(N19697,N19701,N19702);
and and11643(N19698,N19703,N19704);
and and11644(N19699,in2,N19705);
and and11645(N19700,R2,R3);
and and11651(N19711,N19715,N19716);
and and11652(N19712,in1,N19717);
and and11653(N19713,N19718,N19719);
and and11654(N19714,R2,R3);
and and11660(N19725,N19729,N19730);
and and11661(N19726,in1,in2);
and and11662(N19727,N19731,R1);
and and11663(N19728,N19732,R3);
and and11669(N19738,N19742,N19743);
and and11670(N19739,in0,in1);
and and11671(N19740,R0,R1);
and and11672(N19741,N19744,R3);
and and11678(N19751,N19755,N19756);
and and11679(N19752,N19757,in1);
and and11680(N19753,in2,R0);
and and11681(N19754,R1,N19758);
and and11687(N19764,N19768,N19769);
and and11688(N19765,N19770,N19771);
and and11689(N19766,N19772,R1);
and and11690(N19767,R2,N19773);
and and11696(N19777,N19781,N19782);
and and11697(N19778,in1,in2);
and and11698(N19779,R0,N19783);
and and11699(N19780,N19784,R3);
and and11705(N19790,N19794,N19795);
and and11706(N19791,N19796,in1);
and and11707(N19792,in2,R0);
and and11708(N19793,N19797,R2);
and and11714(N19803,N19807,N19808);
and and11715(N19804,in0,in2);
and and11716(N19805,R0,N19809);
and and11717(N19806,R2,R3);
and and11723(N19816,N19820,N19821);
and and11724(N19817,in0,in1);
and and11725(N19818,N19822,R0);
and and11726(N19819,N19823,R2);
and and11732(N19829,N19833,N19834);
and and11733(N19830,N19835,in1);
and and11734(N19831,in2,R0);
and and11735(N19832,N19836,R2);
and and11741(N19842,N19846,N19847);
and and11742(N19843,N19848,in1);
and and11743(N19844,N19849,R0);
and and11744(N19845,N19850,R2);
and and11750(N19855,N19859,N19860);
and and11751(N19856,in0,in1);
and and11752(N19857,in2,N19861);
and and11753(N19858,R2,R3);
and and11759(N19868,N19872,N19873);
and and11760(N19869,in0,N19874);
and and11761(N19870,R0,N19875);
and and11762(N19871,N19876,R3);
and and11768(N19881,N19885,N19886);
and and11769(N19882,N19887,N19888);
and and11770(N19883,in2,R0);
and and11771(N19884,R1,N19889);
and and11777(N19894,N19898,N19899);
and and11778(N19895,N19900,in1);
and and11779(N19896,R0,N19901);
and and11780(N19897,N19902,R3);
and and11786(N19907,N19911,N19912);
and and11787(N19908,in0,N19913);
and and11788(N19909,N19914,R1);
and and11789(N19910,R2,R3);
and and11795(N19920,N19924,N19925);
and and11796(N19921,N19926,in2);
and and11797(N19922,N19927,R1);
and and11798(N19923,R2,R3);
and and11804(N19933,N19937,N19938);
and and11805(N19934,in0,in2);
and and11806(N19935,N19939,R1);
and and11807(N19936,R2,N19940);
and and11813(N19946,N19950,N19951);
and and11814(N19947,N19952,N19953);
and and11815(N19948,in2,R0);
and and11816(N19949,R1,N19954);
and and11822(N19959,N19963,N19964);
and and11823(N19960,N19965,in2);
and and11824(N19961,N19966,R1);
and and11825(N19962,N19967,R3);
and and11831(N19972,N19976,N19977);
and and11832(N19973,N19978,N19979);
and and11833(N19974,in2,R1);
and and11834(N19975,R2,N19980);
and and11840(N19985,N19989,N19990);
and and11841(N19986,N19991,N19992);
and and11842(N19987,in2,R0);
and and11843(N19988,R1,R2);
and and11849(N19998,N20002,N20003);
and and11850(N19999,in0,in1);
and and11851(N20000,in2,N20004);
and and11852(N20001,N20005,N20006);
and and11858(N20011,N20015,N20016);
and and11859(N20012,N20017,in1);
and and11860(N20013,in2,N20018);
and and11861(N20014,N20019,R3);
and and11867(N20024,N20028,N20029);
and and11868(N20025,in0,in1);
and and11869(N20026,in2,R0);
and and11870(N20027,N20030,N20031);
and and11876(N20037,N20041,N20042);
and and11877(N20038,N20043,in1);
and and11878(N20039,N20044,R1);
and and11879(N20040,R2,R3);
and and11885(N20050,N20054,N20055);
and and11886(N20051,in0,N20056);
and and11887(N20052,N20057,R1);
and and11888(N20053,R2,R3);
and and11894(N20063,N20067,N20068);
and and11895(N20064,in1,N20069);
and and11896(N20065,R0,R1);
and and11897(N20066,N20070,R3);
and and11903(N20076,N20080,N20081);
and and11904(N20077,N20082,in2);
and and11905(N20078,R0,R1);
and and11906(N20079,N20083,R3);
and and11912(N20089,N20093,N20094);
and and11913(N20090,N20095,N20096);
and and11914(N20091,N20097,R0);
and and11915(N20092,R1,R2);
and and11921(N20102,N20106,N20107);
and and11922(N20103,N20108,in1);
and and11923(N20104,in2,R0);
and and11924(N20105,R1,N20109);
and and11930(N20115,N20119,N20120);
and and11931(N20116,N20121,in1);
and and11932(N20117,N20122,N20123);
and and11933(N20118,R1,R3);
and and11939(N20128,N20132,N20133);
and and11940(N20129,N20134,in2);
and and11941(N20130,N20135,R1);
and and11942(N20131,R2,N20136);
and and11948(N20141,N20145,N20146);
and and11949(N20142,in0,N20147);
and and11950(N20143,in2,R0);
and and11951(N20144,R1,N20148);
and and11957(N20154,N20158,N20159);
and and11958(N20155,N20160,N20161);
and and11959(N20156,N20162,R1);
and and11960(N20157,R2,R3);
and and11966(N20167,N20171,N20172);
and and11967(N20168,N20173,in1);
and and11968(N20169,in2,N20174);
and and11969(N20170,N20175,R2);
and and11975(N20180,N20184,N20185);
and and11976(N20181,N20186,in1);
and and11977(N20182,N20187,R0);
and and11978(N20183,R1,R2);
and and11984(N20193,N20197,N20198);
and and11985(N20194,in0,N20199);
and and11986(N20195,in2,R0);
and and11987(N20196,R1,N20200);
and and11993(N20206,N20210,N20211);
and and11994(N20207,in0,in1);
and and11995(N20208,N20212,R0);
and and11996(N20209,R1,N20213);
and and12002(N20219,N20223,N20224);
and and12003(N20220,N20225,N20226);
and and12004(N20221,N20227,R0);
and and12005(N20222,R1,R2);
and and12011(N20232,N20236,N20237);
and and12012(N20233,in1,in2);
and and12013(N20234,R0,N20238);
and and12014(N20235,N20239,R3);
and and12020(N20245,N20249,N20250);
and and12021(N20246,in0,in1);
and and12022(N20247,R0,R1);
and and12023(N20248,N20251,R3);
and and12029(N20257,N20261,N20262);
and and12030(N20258,in0,in1);
and and12031(N20259,in2,R1);
and and12032(N20260,N20263,R3);
and and12038(N20269,N20273,N20274);
and and12039(N20270,in0,in1);
and and12040(N20271,N20275,N20276);
and and12041(N20272,R1,R2);
and and12047(N20281,N20285,N20286);
and and12048(N20282,N20287,in1);
and and12049(N20283,in2,N20288);
and and12050(N20284,R1,R2);
and and12056(N20293,N20297,N20298);
and and12057(N20294,in0,in1);
and and12058(N20295,in2,R0);
and and12059(N20296,R1,N20299);
and and12065(N20305,N20309,N20310);
and and12066(N20306,in0,in2);
and and12067(N20307,N20311,R1);
and and12068(N20308,N20312,R3);
and and12074(N20317,N20321,N20322);
and and12075(N20318,in0,in1);
and and12076(N20319,in2,R0);
and and12077(N20320,R2,N20323);
and and12083(N20329,N20333,N20334);
and and12084(N20330,N20335,in1);
and and12085(N20331,in2,R0);
and and12086(N20332,R2,R3);
and and12092(N20341,N20345,N20346);
and and12093(N20342,in0,in1);
and and12094(N20343,N20347,R0);
and and12095(N20344,N20348,R3);
and and12101(N20353,N20357,N20358);
and and12102(N20354,in0,in1);
and and12103(N20355,R0,N20359);
and and12104(N20356,R2,R3);
and and12110(N20365,N20369,N20370);
and and12111(N20366,N20371,in1);
and and12112(N20367,in2,R0);
and and12113(N20368,R2,N20372);
and and12119(N20377,N20381,N20382);
and and12120(N20378,in0,in1);
and and12121(N20379,N20383,R1);
and and12122(N20380,R2,R3);
and and12128(N20389,N20393,N20394);
and and12129(N20390,in1,in2);
and and12130(N20391,R0,R1);
and and12131(N20392,R2,R3);
and and12137(N20401,N20405,N20406);
and and12138(N20402,in1,N20407);
and and12139(N20403,R0,R1);
and and12140(N20404,R2,R3);
and and12146(N20413,N20417,N20418);
and and12147(N20414,in0,in1);
and and12148(N20415,in2,N20419);
and and12149(N20416,R1,N20420);
and and12155(N20425,N20429,N20430);
and and12156(N20426,in0,in1);
and and12157(N20427,N20431,R1);
and and12158(N20428,N20432,R3);
and and12164(N20437,N20441,N20442);
and and12165(N20438,N20443,in2);
and and12166(N20439,R0,R1);
and and12167(N20440,R2,R3);
and and12173(N20449,N20453,N20454);
and and12174(N20450,in0,in1);
and and12175(N20451,R0,R1);
and and12176(N20452,R2,R3);
and and12182(N20461,N20465,N20466);
and and12183(N20462,N20467,in1);
and and12184(N20463,in2,R0);
and and12185(N20464,R1,R2);
and and12191(N20473,N20477,N20478);
and and12192(N20474,N20479,in2);
and and12193(N20475,R0,N20480);
and and12194(N20476,R2,R3);
and and12200(N20485,N20489,N20490);
and and12201(N20486,N20491,N20492);
and and12202(N20487,in2,R0);
and and12203(N20488,R1,N20493);
and and12209(N20497,N20501,N20502);
and and12210(N20498,in0,N20503);
and and12211(N20499,R0,R1);
and and12212(N20500,R2,R3);
and and12218(N20509,N20513,N20514);
and and12219(N20510,in1,in2);
and and12220(N20511,R0,R1);
and and12221(N20512,R2,N20515);
and and12227(N20521,N20525,N20526);
and and12228(N20522,N20527,in2);
and and12229(N20523,N20528,R1);
and and12230(N20524,N20529,R3);
and and12236(N20533,N20537,N20538);
and and12237(N20534,N20539,in2);
and and12238(N20535,R0,N20540);
and and12239(N20536,R2,R3);
and and12245(N20545,N20549,N20550);
and and12246(N20546,in0,N20551);
and and12247(N20547,R0,N20552);
and and12248(N20548,R2,R3);
and and12254(N20557,N20561,N20562);
and and12255(N20558,in0,in1);
and and12256(N20559,N20563,R1);
and and12257(N20560,N20564,R3);
and and12263(N20569,N20573,N20574);
and and12264(N20570,N20575,in1);
and and12265(N20571,in2,N20576);
and and12266(N20572,R1,N20577);
and and12272(N20581,N20585,N20586);
and and12273(N20582,in0,in1);
and and12274(N20583,N20587,R1);
and and12275(N20584,N20588,R3);
and and12281(N20593,N20597,N20598);
and and12282(N20594,N20599,N20600);
and and12283(N20595,in2,R0);
and and12284(N20596,R2,R3);
and and12290(N20605,N20609,N20610);
and and12291(N20606,in0,in1);
and and12292(N20607,in2,N20611);
and and12293(N20608,N20612,R2);
and and12299(N20617,N20621,N20622);
and and12300(N20618,in1,in2);
and and12301(N20619,R0,R1);
and and12302(N20620,R2,N20623);
and and12308(N20629,N20633,N20634);
and and12309(N20630,in0,in1);
and and12310(N20631,N20635,R0);
and and12311(N20632,R1,R3);
and and12317(N20641,N20645,N20646);
and and12318(N20642,in1,in2);
and and12319(N20643,R0,N20647);
and and12320(N20644,R2,R3);
and and12326(N20653,N20657,N20658);
and and12327(N20654,in0,in1);
and and12328(N20655,in2,N20659);
and and12329(N20656,R2,R3);
and and12335(N20665,N20669,N20670);
and and12336(N20666,in0,in1);
and and12337(N20667,in2,R1);
and and12338(N20668,R2,R3);
and and12344(N20676,N20680,N20681);
and and12345(N20677,in0,in1);
and and12346(N20678,in2,R0);
and and12347(N20679,N20682,R3);
and and12353(N20687,N20691,N20692);
and and12354(N20688,in0,in1);
and and12355(N20689,in2,R0);
and and12356(N20690,R1,N20693);
and and12362(N20698,N20702,N20703);
and and12363(N20699,in0,in1);
and and12364(N20700,N20704,R1);
and and12365(N20701,R2,R3);
and and12371(N20709,N20713,N20714);
and and12372(N20710,N20715,in1);
and and12373(N20711,in2,N20716);
and and12374(N20712,R1,R2);
and and12380(N20720,N20724,N20725);
and and12381(N20721,N20726,in1);
and and12382(N20722,in2,R0);
and and12383(N20723,R1,R2);
and and12389(N20731,N20735,N20736);
and and12390(N20732,in0,in1);
and and12391(N20733,in2,R0);
and and12392(N20734,R1,R2);
and and12398(N20741,N20745,N20746);
and and12399(N20742,in0,in2);
and and12400(N20743,R0,R1);
and and12401(N20744,N20747,R3);
and and12407(N20751,N20755,N20756);
and and12408(N20752,in0,in1);
and and12409(N20753,in2,N20757);
and and12410(N20754,R1,R2);
and and12416(N20761,N20765,N20766);
and and12417(N20762,in0,in1);
and and12418(N20763,in2,R0);
and and12419(N20764,R1,R2);
and and12425(N20771,N20775,N20776);
and and12426(N20772,in1,in2);
and and12427(N20773,R0,N20777);
and and12428(N20774,R2,R3);
and and12434(N20781,N20785,N20786);
and and12435(N20782,in0,in1);
and and12436(N20783,in2,R0);
and and12437(N20784,R1,R2);
and and12443(N20791,N20795,N20796);
and and12444(N20792,in0,in1);
and and12445(N20793,in2,R0);
and and12446(N20794,R1,R2);
and and12452(N20801,N20805,N20806);
and and12453(N20802,in1,in2);
and and12454(N20803,R0,R1);
and and12455(N20804,R2,R3);
and and12461(N20811,N20815,N20816);
and and12462(N20812,in1,in2);
and and12463(N20813,R0,R1);
and and12464(N20814,R2,R3);
and and12470(N20821,N20825,N20826);
and and12471(N20822,in0,in1);
and and12472(N20823,in2,R1);
and and12473(N20824,N20827,R3);
and and12479(N20831,N20835,N20836);
and and12480(N20832,in0,in1);
and and12481(N20833,in2,R0);
and and12482(N20834,R2,R3);
and and12488(N20841,N20845,N20846);
and and12489(N20842,in0,in1);
and and12490(N20843,in2,R0);
and and12491(N20844,N20847,R2);
and and12497(N20851,N20855,N20856);
and and12498(N20852,in2,N20857);
and and12499(N20853,N20858,N20859);
and and12500(N20854,N20860,N20861);
and and12505(N20867,N20871,N20872);
and and12506(N20868,N20873,N20874);
and and12507(N20869,N20875,N20876);
and and12508(N20870,N20877,R4);
and and12513(N20883,N20887,N20888);
and and12514(N20884,N20889,N20890);
and and12515(N20885,N20891,N20892);
and and12516(N20886,R4,R5);
and and12521(N20898,N20902,N20903);
and and12522(N20899,N20904,N20905);
and and12523(N20900,N20906,N20907);
and and12524(N20901,R3,N20908);
and and12529(N20913,N20917,N20918);
and and12530(N20914,N20919,R0);
and and12531(N20915,N20920,N20921);
and and12532(N20916,R3,N20922);
and and12537(N20928,N20932,N20933);
and and12538(N20929,N20934,R0);
and and12539(N20930,N20935,N20936);
and and12540(N20931,N20937,N20938);
and and12545(N20943,N20947,N20948);
and and12546(N20944,N20949,N20950);
and and12547(N20945,N20951,N20952);
and and12548(N20946,R4,N20953);
and and12553(N20958,N20962,N20963);
and and12554(N20959,N20964,R0);
and and12555(N20960,R2,N20965);
and and12556(N20961,N20966,N20967);
and and12561(N20973,N20977,in0);
and and12562(N20974,N20978,N20979);
and and12563(N20975,N20980,N20981);
and and12564(N20976,N20982,R4);
and and12569(N20988,N20992,N20993);
and and12570(N20989,in1,N20994);
and and12571(N20990,N20995,N20996);
and and12572(N20991,R3,N20997);
and and12577(N21003,N21007,in0);
and and12578(N21004,N21008,N21009);
and and12579(N21005,R0,N21010);
and and12580(N21006,N21011,N21012);
and and12585(N21018,N21022,N21023);
and and12586(N21019,in2,R0);
and and12587(N21020,N21024,N21025);
and and12588(N21021,N21026,N21027);
and and12593(N21033,N21037,in1);
and and12594(N21034,N21038,R0);
and and12595(N21035,N21039,N21040);
and and12596(N21036,N21041,N21042);
and and12601(N21048,N21052,N21053);
and and12602(N21049,N21054,N21055);
and and12603(N21050,N21056,N21057);
and and12604(N21051,R4,N21058);
and and12609(N21063,N21067,N21068);
and and12610(N21064,in1,N21069);
and and12611(N21065,N21070,N21071);
and and12612(N21066,N21072,R4);
and and12617(N21078,N21082,in0);
and and12618(N21079,N21083,N21084);
and and12619(N21080,N21085,R2);
and and12620(N21081,R4,N21086);
and and12625(N21092,N21096,in1);
and and12626(N21093,N21097,N21098);
and and12627(N21094,R1,R2);
and and12628(N21095,N21099,N21100);
and and12633(N21106,N21110,in0);
and and12634(N21107,N21111,N21112);
and and12635(N21108,R1,R2);
and and12636(N21109,N21113,N21114);
and and12641(N21120,N21124,N21125);
and and12642(N21121,N21126,N21127);
and and12643(N21122,R2,N21128);
and and12644(N21123,R4,R5);
and and12649(N21134,N21138,in1);
and and12650(N21135,N21139,N21140);
and and12651(N21136,R2,N21141);
and and12652(N21137,N21142,N21143);
and and12657(N21148,N21152,in0);
and and12658(N21149,N21153,N21154);
and and12659(N21150,R2,N21155);
and and12660(N21151,N21156,N21157);
and and12665(N21162,N21166,N21167);
and and12666(N21163,in1,N21168);
and and12667(N21164,N21169,R2);
and and12668(N21165,R3,N21170);
and and12673(N21176,N21180,N21181);
and and12674(N21177,N21182,N21183);
and and12675(N21178,R2,R3);
and and12676(N21179,N21184,R5);
and and12681(N21190,N21194,N21195);
and and12682(N21191,in2,N21196);
and and12683(N21192,R1,N21197);
and and12684(N21193,N21198,N21199);
and and12689(N21204,N21208,in0);
and and12690(N21205,N21209,R0);
and and12691(N21206,N21210,N21211);
and and12692(N21207,N21212,N21213);
and and12697(N21218,N21222,N21223);
and and12698(N21219,N21224,N21225);
and and12699(N21220,N21226,R3);
and and12700(N21221,N21227,R5);
and and12705(N21232,N21236,N21237);
and and12706(N21233,N21238,N21239);
and and12707(N21234,N21240,R2);
and and12708(N21235,N21241,R5);
and and12713(N21246,N21250,in0);
and and12714(N21247,N21251,N21252);
and and12715(N21248,N21253,N21254);
and and12716(N21249,R4,N21255);
and and12721(N21260,N21264,in0);
and and12722(N21261,N21265,N21266);
and and12723(N21262,N21267,R1);
and and12724(N21263,N21268,R5);
and and12729(N21274,N21278,in1);
and and12730(N21275,N21279,R1);
and and12731(N21276,N21280,N21281);
and and12732(N21277,R4,N21282);
and and12737(N21288,N21292,in0);
and and12738(N21289,N21293,R1);
and and12739(N21290,N21294,N21295);
and and12740(N21291,R4,N21296);
and and12745(N21302,N21306,N21307);
and and12746(N21303,R0,N21308);
and and12747(N21304,N21309,R3);
and and12748(N21305,R4,N21310);
and and12753(N21316,N21320,N21321);
and and12754(N21317,N21322,N21323);
and and12755(N21318,R1,N21324);
and and12756(N21319,N21325,R4);
and and12761(N21330,N21334,N21335);
and and12762(N21331,N21336,N21337);
and and12763(N21332,R1,N21338);
and and12764(N21333,R4,N21339);
and and12769(N21344,N21348,N21349);
and and12770(N21345,N21350,in2);
and and12771(N21346,R0,N21351);
and and12772(N21347,N21352,R4);
and and12777(N21358,N21362,in0);
and and12778(N21359,N21363,R0);
and and12779(N21360,N21364,N21365);
and and12780(N21361,N21366,R4);
and and12785(N21372,N21376,in0);
and and12786(N21373,N21377,in2);
and and12787(N21374,N21378,R3);
and and12788(N21375,N21379,N21380);
and and12793(N21386,N21390,N21391);
and and12794(N21387,N21392,R0);
and and12795(N21388,N21393,R2);
and and12796(N21389,N21394,N21395);
and and12801(N21400,N21404,N21405);
and and12802(N21401,N21406,N21407);
and and12803(N21402,R1,R2);
and and12804(N21403,R3,N21408);
and and12809(N21414,N21418,in1);
and and12810(N21415,N21419,R0);
and and12811(N21416,N21420,N21421);
and and12812(N21417,N21422,N21423);
and and12817(N21428,N21432,N21433);
and and12818(N21429,N21434,N21435);
and and12819(N21430,N21436,R3);
and and12820(N21431,N21437,R5);
and and12825(N21442,N21446,in0);
and and12826(N21443,N21447,N21448);
and and12827(N21444,R0,N21449);
and and12828(N21445,N21450,N21451);
and and12833(N21456,N21460,in0);
and and12834(N21457,N21461,N21462);
and and12835(N21458,R0,R2);
and and12836(N21459,N21463,N21464);
and and12841(N21470,N21474,in0);
and and12842(N21471,N21475,N21476);
and and12843(N21472,R1,N21477);
and and12844(N21473,N21478,R5);
and and12849(N21484,N21488,in0);
and and12850(N21485,N21489,N21490);
and and12851(N21486,R1,N21491);
and and12852(N21487,N21492,R5);
and and12857(N21498,N21502,N21503);
and and12858(N21499,N21504,N21505);
and and12859(N21500,N21506,R1);
and and12860(N21501,R4,N21507);
and and12865(N21512,N21516,in0);
and and12866(N21513,in2,R0);
and and12867(N21514,N21517,N21518);
and and12868(N21515,N21519,N21520);
and and12873(N21526,N21530,N21531);
and and12874(N21527,N21532,R0);
and and12875(N21528,R1,R2);
and and12876(N21529,R3,N21533);
and and12881(N21539,N21543,in1);
and and12882(N21540,N21544,R0);
and and12883(N21541,R1,N21545);
and and12884(N21542,N21546,N21547);
and and12889(N21552,N21556,in0);
and and12890(N21553,N21557,N21558);
and and12891(N21554,R0,R1);
and and12892(N21555,R3,N21559);
and and12897(N21565,N21569,in0);
and and12898(N21566,N21570,R0);
and and12899(N21567,N21571,N21572);
and and12900(N21568,R3,N21573);
and and12905(N21578,N21582,in0);
and and12906(N21579,N21583,N21584);
and and12907(N21580,N21585,R3);
and and12908(N21581,R4,R5);
and and12913(N21591,N21595,N21596);
and and12914(N21592,N21597,N21598);
and and12915(N21593,R0,R1);
and and12916(N21594,N21599,R3);
and and12921(N21604,N21608,N21609);
and and12922(N21605,in1,in2);
and and12923(N21606,N21610,N21611);
and and12924(N21607,R3,N21612);
and and12929(N21617,N21621,in0);
and and12930(N21618,N21622,in2);
and and12931(N21619,N21623,N21624);
and and12932(N21620,R3,N21625);
and and12937(N21630,N21634,N21635);
and and12938(N21631,in2,N21636);
and and12939(N21632,N21637,R2);
and and12940(N21633,R3,N21638);
and and12945(N21643,N21647,N21648);
and and12946(N21644,N21649,in2);
and and12947(N21645,R0,N21650);
and and12948(N21646,R3,N21651);
and and12953(N21656,N21660,N21661);
and and12954(N21657,in1,N21662);
and and12955(N21658,N21663,R1);
and and12956(N21659,R2,R4);
and and12961(N21669,N21673,in0);
and and12962(N21670,in1,R0);
and and12963(N21671,N21674,R3);
and and12964(N21672,N21675,N21676);
and and12969(N21682,N21686,N21687);
and and12970(N21683,N21688,in2);
and and12971(N21684,N21689,N21690);
and and12972(N21685,R3,N21691);
and and12977(N21695,N21699,N21700);
and and12978(N21696,N21701,R0);
and and12979(N21697,R2,N21702);
and and12980(N21698,N21703,N21704);
and and12985(N21708,N21712,N21713);
and and12986(N21709,N21714,R0);
and and12987(N21710,N21715,R3);
and and12988(N21711,N21716,N21717);
and and12993(N21721,N21725,in0);
and and12994(N21722,N21726,N21727);
and and12995(N21723,R2,N21728);
and and12996(N21724,N21729,R5);
and and13001(N21734,N21738,N21739);
and and13002(N21735,N21740,in2);
and and13003(N21736,R2,N21741);
and and13004(N21737,N21742,R5);
and and13009(N21747,N21751,N21752);
and and13010(N21748,in1,in2);
and and13011(N21749,N21753,N21754);
and and13012(N21750,R4,N21755);
and and13017(N21760,N21764,in0);
and and13018(N21761,N21765,N21766);
and and13019(N21762,N21767,R3);
and and13020(N21763,R4,N21768);
and and13025(N21773,N21777,in1);
and and13026(N21774,N21778,N21779);
and and13027(N21775,N21780,R3);
and and13028(N21776,R4,N21781);
and and13033(N21786,N21790,N21791);
and and13034(N21787,in2,N21792);
and and13035(N21788,N21793,R3);
and and13036(N21789,R4,N21794);
and and13041(N21799,N21803,in0);
and and13042(N21800,in2,R0);
and and13043(N21801,N21804,R2);
and and13044(N21802,N21805,N21806);
and and13049(N21812,N21816,in1);
and and13050(N21813,N21817,N21818);
and and13051(N21814,R1,N21819);
and and13052(N21815,N21820,R5);
and and13057(N21825,N21829,in0);
and and13058(N21826,N21830,N21831);
and and13059(N21827,R1,N21832);
and and13060(N21828,N21833,R5);
and and13065(N21838,N21842,N21843);
and and13066(N21839,N21844,N21845);
and and13067(N21840,N21846,R3);
and and13068(N21841,R4,N21847);
and and13073(N21851,N21855,N21856);
and and13074(N21852,N21857,R0);
and and13075(N21853,R1,N21858);
and and13076(N21854,N21859,R4);
and and13081(N21864,N21868,in0);
and and13082(N21865,in1,in2);
and and13083(N21866,N21869,N21870);
and and13084(N21867,N21871,R4);
and and13089(N21877,N21881,in0);
and and13090(N21878,N21882,N21883);
and and13091(N21879,R1,N21884);
and and13092(N21880,R4,N21885);
and and13097(N21890,N21894,in0);
and and13098(N21891,in2,R0);
and and13099(N21892,N21895,N21896);
and and13100(N21893,N21897,N21898);
and and13105(N21903,N21907,in0);
and and13106(N21904,in1,R0);
and and13107(N21905,N21908,N21909);
and and13108(N21906,N21910,N21911);
and and13113(N21916,N21920,in1);
and and13114(N21917,in2,R0);
and and13115(N21918,N21921,N21922);
and and13116(N21919,N21923,N21924);
and and13121(N21929,N21933,N21934);
and and13122(N21930,N21935,R0);
and and13123(N21931,R1,N21936);
and and13124(N21932,N21937,N21938);
and and13129(N21942,N21946,N21947);
and and13130(N21943,N21948,N21949);
and and13131(N21944,R2,R3);
and and13132(N21945,N21950,N21951);
and and13137(N21955,N21959,in0);
and and13138(N21956,N21960,N21961);
and and13139(N21957,R1,N21962);
and and13140(N21958,N21963,R4);
and and13145(N21968,N21972,in1);
and and13146(N21969,N21973,N21974);
and and13147(N21970,R1,N21975);
and and13148(N21971,N21976,R4);
and and13153(N21981,N21985,in0);
and and13154(N21982,N21986,in2);
and and13155(N21983,N21987,R1);
and and13156(N21984,N21988,N21989);
and and13161(N21994,N21998,in0);
and and13162(N21995,in1,N21999);
and and13163(N21996,N22000,R1);
and and13164(N21997,N22001,N22002);
and and13169(N22007,N22011,in1);
and and13170(N22008,in2,N22012);
and and13171(N22009,R1,N22013);
and and13172(N22010,N22014,N22015);
and and13177(N22020,N22024,in1);
and and13178(N22021,N22025,N22026);
and and13179(N22022,N22027,R2);
and and13180(N22023,R3,N22028);
and and13185(N22033,N22037,N22038);
and and13186(N22034,in2,N22039);
and and13187(N22035,N22040,R2);
and and13188(N22036,R3,N22041);
and and13193(N22046,N22050,in0);
and and13194(N22047,N22051,N22052);
and and13195(N22048,N22053,R2);
and and13196(N22049,R3,N22054);
and and13201(N22059,N22063,N22064);
and and13202(N22060,in1,R0);
and and13203(N22061,N22065,R2);
and and13204(N22062,N22066,R5);
and and13209(N22072,N22076,N22077);
and and13210(N22073,in2,N22078);
and and13211(N22074,N22079,R2);
and and13212(N22075,N22080,R4);
and and13217(N22085,N22089,in0);
and and13218(N22086,N22090,N22091);
and and13219(N22087,N22092,R2);
and and13220(N22088,N22093,R4);
and and13225(N22098,N22102,in0);
and and13226(N22099,N22103,N22104);
and and13227(N22100,R2,N22105);
and and13228(N22101,R4,R5);
and and13233(N22111,N22115,in0);
and and13234(N22112,in2,N22116);
and and13235(N22113,R2,N22117);
and and13236(N22114,N22118,N22119);
and and13241(N22124,N22128,in1);
and and13242(N22125,N22129,N22130);
and and13243(N22126,R2,R3);
and and13244(N22127,N22131,R5);
and and13249(N22137,N22141,N22142);
and and13250(N22138,in1,N22143);
and and13251(N22139,R1,R2);
and and13252(N22140,N22144,N22145);
and and13257(N22150,N22154,in0);
and and13258(N22151,N22155,N22156);
and and13259(N22152,N22157,R3);
and and13260(N22153,N22158,R5);
and and13265(N22163,N22167,in0);
and and13266(N22164,in2,R0);
and and13267(N22165,R1,N22168);
and and13268(N22166,N22169,N22170);
and and13273(N22176,N22180,in0);
and and13274(N22177,in1,N22181);
and and13275(N22178,N22182,N22183);
and and13276(N22179,R4,N22184);
and and13281(N22189,N22193,N22194);
and and13282(N22190,N22195,R1);
and and13283(N22191,N22196,N22197);
and and13284(N22192,R4,R5);
and and13289(N22202,N22206,N22207);
and and13290(N22203,in1,N22208);
and and13291(N22204,R1,N22209);
and and13292(N22205,N22210,R4);
and and13297(N22215,N22219,in0);
and and13298(N22216,in2,R0);
and and13299(N22217,N22220,N22221);
and and13300(N22218,R4,N22222);
and and13305(N22228,N22232,N22233);
and and13306(N22229,N22234,N22235);
and and13307(N22230,R1,R2);
and and13308(N22231,R3,R4);
and and13313(N22240,N22244,in0);
and and13314(N22241,in1,N22245);
and and13315(N22242,N22246,R2);
and and13316(N22243,R3,R4);
and and13321(N22252,N22256,in0);
and and13322(N22253,R0,N22257);
and and13323(N22254,R2,R3);
and and13324(N22255,R4,N22258);
and and13329(N22264,N22268,N22269);
and and13330(N22265,N22270,R1);
and and13331(N22266,N22271,R3);
and and13332(N22267,R4,N22272);
and and13337(N22276,N22280,N22281);
and and13338(N22277,in2,R0);
and and13339(N22278,N22282,R2);
and and13340(N22279,N22283,R4);
and and13345(N22288,N22292,in1);
and and13346(N22289,N22293,R0);
and and13347(N22290,N22294,R2);
and and13348(N22291,R4,N22295);
and and13353(N22300,N22304,in0);
and and13354(N22301,in1,in2);
and and13355(N22302,N22305,R2);
and and13356(N22303,R4,N22306);
and and13361(N22312,N22316,in0);
and and13362(N22313,in1,in2);
and and13363(N22314,R1,R2);
and and13364(N22315,N22317,N22318);
and and13369(N22324,N22328,N22329);
and and13370(N22325,in2,N22330);
and and13371(N22326,R1,R2);
and and13372(N22327,R3,N22331);
and and13377(N22336,N22340,in0);
and and13378(N22337,in1,R0);
and and13379(N22338,R1,N22341);
and and13380(N22339,N22342,N22343);
and and13385(N22348,N22352,in0);
and and13386(N22349,in1,N22353);
and and13387(N22350,N22354,R1);
and and13388(N22351,R2,N22355);
and and13393(N22360,N22364,in0);
and and13394(N22361,N22365,R0);
and and13395(N22362,R1,N22366);
and and13396(N22363,N22367,R5);
and and13401(N22372,N22376,in0);
and and13402(N22373,N22377,R0);
and and13403(N22374,R1,R2);
and and13404(N22375,N22378,N22379);
and and13409(N22384,N22388,in1);
and and13410(N22385,N22389,R1);
and and13411(N22386,N22390,N22391);
and and13412(N22387,R4,R5);
and and13417(N22396,N22400,N22401);
and and13418(N22397,in1,R0);
and and13419(N22398,N22402,N22403);
and and13420(N22399,R3,N22404);
and and13425(N22408,N22412,N22413);
and and13426(N22409,in1,in2);
and and13427(N22410,N22414,N22415);
and and13428(N22411,R2,R5);
and and13433(N22420,N22424,in0);
and and13434(N22421,N22425,in2);
and and13435(N22422,R1,N22426);
and and13436(N22423,N22427,R5);
and and13441(N22432,N22436,N22437);
and and13442(N22433,in2,R0);
and and13443(N22434,N22438,R2);
and and13444(N22435,R3,N22439);
and and13449(N22444,N22448,N22449);
and and13450(N22445,in1,N22450);
and and13451(N22446,R0,R1);
and and13452(N22447,N22451,R4);
and and13457(N22456,N22460,N22461);
and and13458(N22457,N22462,R0);
and and13459(N22458,R1,R2);
and and13460(N22459,R4,N22463);
and and13465(N22468,N22472,in0);
and and13466(N22469,N22473,N22474);
and and13467(N22470,R1,N22475);
and and13468(N22471,R3,R4);
and and13473(N22480,N22484,in0);
and and13474(N22481,in1,N22485);
and and13475(N22482,R1,N22486);
and and13476(N22483,N22487,R4);
and and13481(N22492,N22496,in0);
and and13482(N22493,N22497,R1);
and and13483(N22494,N22498,N22499);
and and13484(N22495,R4,R5);
and and13489(N22504,N22508,in2);
and and13490(N22505,N22509,N22510);
and and13491(N22506,R2,N22511);
and and13492(N22507,R4,N22512);
and and13497(N22516,N22520,in1);
and and13498(N22517,in2,N22521);
and and13499(N22518,R1,R2);
and and13500(N22519,N22522,N22523);
and and13505(N22528,N22532,N22533);
and and13506(N22529,N22534,N22535);
and and13507(N22530,R1,R3);
and and13508(N22531,R4,R5);
and and13513(N22540,N22544,in0);
and and13514(N22541,in1,N22545);
and and13515(N22542,R1,R2);
and and13516(N22543,N22546,N22547);
and and13521(N22552,N22556,N22557);
and and13522(N22553,in2,R0);
and and13523(N22554,N22558,R2);
and and13524(N22555,R3,N22559);
and and13529(N22564,N22568,in0);
and and13530(N22565,in1,N22569);
and and13531(N22566,R0,N22570);
and and13532(N22567,R2,N22571);
and and13537(N22576,N22580,in0);
and and13538(N22577,N22581,R0);
and and13539(N22578,R1,R2);
and and13540(N22579,N22582,N22583);
and and13545(N22588,N22592,in0);
and and13546(N22589,N22593,N22594);
and and13547(N22590,R1,R2);
and and13548(N22591,N22595,R4);
and and13553(N22600,N22604,N22605);
and and13554(N22601,in1,N22606);
and and13555(N22602,R1,R2);
and and13556(N22603,N22607,R4);
and and13561(N22612,N22616,in1);
and and13562(N22613,N22617,R0);
and and13563(N22614,N22618,R2);
and and13564(N22615,N22619,R4);
and and13569(N22624,N22628,in0);
and and13570(N22625,N22629,R0);
and and13571(N22626,N22630,R2);
and and13572(N22627,N22631,R4);
and and13577(N22636,N22640,in0);
and and13578(N22637,N22641,N22642);
and and13579(N22638,R2,R3);
and and13580(N22639,R4,N22643);
and and13585(N22648,N22652,in0);
and and13586(N22649,N22653,R0);
and and13587(N22650,N22654,R3);
and and13588(N22651,R4,R5);
and and13593(N22660,N22664,in1);
and and13594(N22661,N22665,R0);
and and13595(N22662,N22666,R3);
and and13596(N22663,R4,N22667);
and and13601(N22672,N22676,N22677);
and and13602(N22673,N22678,in2);
and and13603(N22674,R0,R1);
and and13604(N22675,N22679,R3);
and and13609(N22684,N22688,N22689);
and and13610(N22685,N22690,in2);
and and13611(N22686,R0,R1);
and and13612(N22687,R3,N22691);
and and13617(N22696,N22700,in0);
and and13618(N22697,N22701,R0);
and and13619(N22698,N22702,R3);
and and13620(N22699,N22703,N22704);
and and13625(N22708,N22712,in0);
and and13626(N22709,in2,N22713);
and and13627(N22710,R2,N22714);
and and13628(N22711,N22715,R5);
and and13633(N22720,N22724,in1);
and and13634(N22721,in2,N22725);
and and13635(N22722,N22726,R3);
and and13636(N22723,R4,N22727);
and and13641(N22732,N22736,in0);
and and13642(N22733,in1,in2);
and and13643(N22734,N22737,R1);
and and13644(N22735,N22738,N22739);
and and13649(N22744,N22748,in0);
and and13650(N22745,N22749,N22750);
and and13651(N22746,N22751,R3);
and and13652(N22747,R4,N22752);
and and13657(N22756,N22760,in0);
and and13658(N22757,N22761,N22762);
and and13659(N22758,N22763,R3);
and and13660(N22759,R4,N22764);
and and13665(N22768,N22772,in0);
and and13666(N22769,N22773,N22774);
and and13667(N22770,R0,R1);
and and13668(N22771,N22775,R4);
and and13673(N22780,N22784,in2);
and and13674(N22781,N22785,N22786);
and and13675(N22782,R2,R3);
and and13676(N22783,N22787,N22788);
and and13681(N22792,N22796,in0);
and and13682(N22793,in1,in2);
and and13683(N22794,N22797,R1);
and and13684(N22795,N22798,N22799);
and and13689(N22804,N22808,in0);
and and13690(N22805,in2,N22809);
and and13691(N22806,N22810,R2);
and and13692(N22807,R3,N22811);
and and13697(N22816,N22820,in0);
and and13698(N22817,N22821,N22822);
and and13699(N22818,R0,R1);
and and13700(N22819,R2,R5);
and and13705(N22828,N22832,in0);
and and13706(N22829,N22833,in2);
and and13707(N22830,R0,R1);
and and13708(N22831,R2,R3);
and and13713(N22839,N22843,in0);
and and13714(N22840,in1,N22844);
and and13715(N22841,R0,R1);
and and13716(N22842,R2,R3);
and and13721(N22850,N22854,N22855);
and and13722(N22851,in1,in2);
and and13723(N22852,R0,R1);
and and13724(N22853,N22856,R3);
and and13729(N22861,N22865,N22866);
and and13730(N22862,in2,R0);
and and13731(N22863,N22867,R3);
and and13732(N22864,R4,R5);
and and13737(N22872,N22876,in0);
and and13738(N22873,N22877,R0);
and and13739(N22874,N22878,R3);
and and13740(N22875,R4,N22879);
and and13745(N22883,N22887,in0);
and and13746(N22884,in1,N22888);
and and13747(N22885,N22889,R2);
and and13748(N22886,R3,R5);
and and13753(N22894,N22898,in0);
and and13754(N22895,in1,in2);
and and13755(N22896,R1,N22899);
and and13756(N22897,N22900,N22901);
and and13761(N22905,N22909,in1);
and and13762(N22906,in2,R0);
and and13763(N22907,R1,N22910);
and and13764(N22908,N22911,R5);
and and13769(N22916,N22920,in1);
and and13770(N22917,in2,R0);
and and13771(N22918,R1,R2);
and and13772(N22919,N22921,N22922);
and and13777(N22927,N22931,in0);
and and13778(N22928,in1,N22932);
and and13779(N22929,R0,R1);
and and13780(N22930,R2,N22933);
and and13785(N22938,N22942,in0);
and and13786(N22939,N22943,R0);
and and13787(N22940,R1,R2);
and and13788(N22941,R3,N22944);
and and13793(N22949,N22953,in1);
and and13794(N22950,N22954,R0);
and and13795(N22951,R1,R2);
and and13796(N22952,R3,N22955);
and and13801(N22960,N22964,in0);
and and13802(N22961,in2,R0);
and and13803(N22962,R2,N22965);
and and13804(N22963,N22966,N22967);
and and13809(N22971,N22975,in0);
and and13810(N22972,in1,R0);
and and13811(N22973,R2,N22976);
and and13812(N22974,N22977,N22978);
and and13817(N22982,N22986,in0);
and and13818(N22983,in2,N22987);
and and13819(N22984,N22988,R2);
and and13820(N22985,R3,R4);
and and13825(N22993,N22997,in0);
and and13826(N22994,N22998,N22999);
and and13827(N22995,R1,R3);
and and13828(N22996,N23000,R5);
and and13833(N23004,N23008,in0);
and and13834(N23005,N23009,in2);
and and13835(N23006,R0,R1);
and and13836(N23007,N23010,R4);
and and13841(N23015,N23019,in0);
and and13842(N23016,in1,R0);
and and13843(N23017,R1,N23020);
and and13844(N23018,N23021,R4);
and and13849(N23026,N23030,in1);
and and13850(N23027,in2,R0);
and and13851(N23028,R1,N23031);
and and13852(N23029,N23032,R4);
and and13857(N23037,N23041,N23042);
and and13858(N23038,in2,R0);
and and13859(N23039,R1,N23043);
and and13860(N23040,R4,N23044);
and and13865(N23048,N23052,in1);
and and13866(N23049,N23053,R0);
and and13867(N23050,R1,R2);
and and13868(N23051,N23054,R4);
and and13873(N23059,N23063,in0);
and and13874(N23060,N23064,R0);
and and13875(N23061,R1,R2);
and and13876(N23062,N23065,R4);
and and13881(N23070,N23074,in0);
and and13882(N23071,in1,N23075);
and and13883(N23072,R1,R3);
and and13884(N23073,R4,N23076);
and and13889(N23081,N23085,in0);
and and13890(N23082,in1,in2);
and and13891(N23083,N23086,R1);
and and13892(N23084,R4,N23087);
and and13897(N23092,N23096,N23097);
and and13898(N23093,N23098,R1);
and and13899(N23094,N23099,R3);
and and13900(N23095,R4,R5);
and and13905(N23103,N23107,in0);
and and13906(N23104,in1,R0);
and and13907(N23105,N23108,R2);
and and13908(N23106,R3,N23109);
and and13913(N23114,N23118,in0);
and and13914(N23115,N23119,R1);
and and13915(N23116,R2,N23120);
and and13916(N23117,R4,R5);
and and13921(N23125,N23129,in0);
and and13922(N23126,in1,N23130);
and and13923(N23127,R0,R2);
and and13924(N23128,N23131,R4);
and and13929(N23136,N23140,in0);
and and13930(N23137,in1,N23141);
and and13931(N23138,R0,R1);
and and13932(N23139,R2,N23142);
and and13937(N23147,N23151,in1);
and and13938(N23148,in2,R0);
and and13939(N23149,R1,R2);
and and13940(N23150,N23152,N23153);
and and13945(N23158,N23162,in0);
and and13946(N23159,N23163,in2);
and and13947(N23160,N23164,R1);
and and13948(N23161,R2,N23165);
and and13953(N23169,N23173,in0);
and and13954(N23170,N23174,in2);
and and13955(N23171,R0,N23175);
and and13956(N23172,R3,R4);
and and13961(N23180,N23184,in1);
and and13962(N23181,in2,R0);
and and13963(N23182,R1,N23185);
and and13964(N23183,R4,R5);
and and13969(N23191,N23195,in0);
and and13970(N23192,N23196,R1);
and and13971(N23193,R2,R3);
and and13972(N23194,N23197,R5);
and and13977(N23202,N23206,N23207);
and and13978(N23203,in2,R1);
and and13979(N23204,R2,R3);
and and13980(N23205,N23208,R5);
and and13985(N23213,N23217,in0);
and and13986(N23214,in1,in2);
and and13987(N23215,N23218,R2);
and and13988(N23216,N23219,R4);
and and13993(N23224,N23228,in0);
and and13994(N23225,in1,in2);
and and13995(N23226,N23229,R1);
and and13996(N23227,R2,R5);
and and14001(N23235,N23239,in0);
and and14002(N23236,N23240,in2);
and and14003(N23237,R0,N23241);
and and14004(N23238,R3,R4);
and and14009(N23246,N23250,in0);
and and14010(N23247,in1,in2);
and and14011(N23248,R0,R1);
and and14012(N23249,R2,N23251);
and and14017(N23257,N23261,in0);
and and14018(N23258,N23262,R0);
and and14019(N23259,N23263,R3);
and and14020(N23260,R4,N23264);
and and14025(N23268,N23272,in1);
and and14026(N23269,in2,R0);
and and14027(N23270,N23273,N23274);
and and14028(N23271,R3,N23275);
and and14033(N23279,N23283,in0);
and and14034(N23280,in1,N23284);
and and14035(N23281,N23285,R1);
and and14036(N23282,R2,N23286);
and and14041(N23290,N23294,in1);
and and14042(N23291,in2,N23295);
and and14043(N23292,R1,N23296);
and and14044(N23293,R4,R5);
and and14049(N23301,N23305,in1);
and and14050(N23302,R0,N23306);
and and14051(N23303,R2,R3);
and and14052(N23304,R4,N23307);
and and14057(N23312,N23316,in2);
and and14058(N23313,R0,N23317);
and and14059(N23314,R2,N23318);
and and14060(N23315,R4,R5);
and and14065(N23323,N23327,in0);
and and14066(N23324,in2,R1);
and and14067(N23325,N23328,N23329);
and and14068(N23326,R4,R5);
and and14073(N23334,N23338,in0);
and and14074(N23335,N23339,in2);
and and14075(N23336,R1,N23340);
and and14076(N23337,R4,R5);
and and14081(N23345,N23349,in1);
and and14082(N23346,in2,N23350);
and and14083(N23347,R1,N23351);
and and14084(N23348,R4,R5);
and and14089(N23356,N23360,in0);
and and14090(N23357,in1,in2);
and and14091(N23358,R0,R1);
and and14092(N23359,N23361,N23362);
and and14097(N23367,N23371,in0);
and and14098(N23368,in1,in2);
and and14099(N23369,N23372,R1);
and and14100(N23370,R2,N23373);
and and14105(N23378,N23382,in0);
and and14106(N23379,in1,in2);
and and14107(N23380,R0,R2);
and and14108(N23381,N23383,N23384);
and and14113(N23389,N23393,in0);
and and14114(N23390,in1,N23394);
and and14115(N23391,N23395,R2);
and and14116(N23392,R3,R5);
and and14121(N23400,N23404,in0);
and and14122(N23401,in2,N23405);
and and14123(N23402,R1,R2);
and and14124(N23403,R3,R5);
and and14129(N23410,N23414,in0);
and and14130(N23411,N23415,R0);
and and14131(N23412,R1,R2);
and and14132(N23413,R3,R5);
and and14137(N23420,N23424,in0);
and and14138(N23421,in1,R0);
and and14139(N23422,N23425,R3);
and and14140(N23423,R4,R5);
and and14145(N23430,N23434,in1);
and and14146(N23431,N23435,R0);
and and14147(N23432,R1,R2);
and and14148(N23433,R3,R4);
and and14153(N23440,N23444,in0);
and and14154(N23441,N23445,R0);
and and14155(N23442,R1,R2);
and and14156(N23443,R3,R4);
and and14161(N23450,N23454,in0);
and and14162(N23451,N23455,R0);
and and14163(N23452,R2,R3);
and and14164(N23453,N23456,R5);
and and14169(N23460,N23464,N23465);
and and14170(N23461,in1,R0);
and and14171(N23462,R1,R3);
and and14172(N23463,N23466,R5);
and and14177(N23470,N23474,in0);
and and14178(N23471,N23475,R0);
and and14179(N23472,R1,R2);
and and14180(N23473,N23476,R5);
and and14185(N23480,N23484,N23485);
and and14186(N23481,in1,R0);
and and14187(N23482,R1,R2);
and and14188(N23483,N23486,R5);
and and14193(N23490,N23494,N23495);
and and14194(N23491,in2,R0);
and and14195(N23492,R1,R2);
and and14196(N23493,N23496,R5);
and and14201(N23500,N23504,in1);
and and14202(N23501,N23505,N23506);
and and14203(N23502,R1,R3);
and and14204(N23503,R4,R5);
and and14209(N23510,N23514,in0);
and and14210(N23511,N23515,in2);
and and14211(N23512,R1,R3);
and and14212(N23513,R4,R5);
and and14217(N23520,N23524,in0);
and and14218(N23521,N23525,N23526);
and and14219(N23522,R1,R2);
and and14220(N23523,R3,R4);
and and14225(N23530,N23534,in0);
and and14226(N23531,N23535,R1);
and and14227(N23532,R2,R3);
and and14228(N23533,N23536,R5);
and and14233(N23540,N23544,in0);
and and14234(N23541,in1,in2);
and and14235(N23542,R0,R1);
and and14236(N23543,N23545,R3);
and and14241(N23550,N23554,in0);
and and14242(N23551,in1,in2);
and and14243(N23552,R0,N23555);
and and14244(N23553,R2,R3);
and and14249(N23559,N23563,in0);
and and14250(N23560,in1,N23564);
and and14251(N23561,R2,R3);
and and14252(N23562,R4,R5);
and and14257(N23568,N23572,in0);
and and14258(N23569,N23573,R0);
and and14259(N23570,R1,R2);
and and14260(N23571,R3,R4);
and and14265(N23577,N23581,in0);
and and14266(N23578,in1,in2);
and and14267(N23579,R1,R2);
and and14268(N23580,R3,R4);
and and14273(N23586,N23590,in0);
and and14274(N23587,N23591,in2);
and and14275(N23588,R0,R1);
and and14276(N23589,R2,R5);
and and14281(N23595,N23599,in0);
and and14282(N23596,in1,in2);
and and14283(N23597,R1,R2);
and and14284(N23598,R3,R5);
and and14289(N23604,N23608,in0);
and and14290(N23605,in2,R0);
and and14291(N23606,R1,R2);
and and14292(N23607,R3,R4);
and and14297(N23613,N23617,in0);
and and14298(N23614,in1,N23618);
and and14299(N23615,R0,R1);
and and14300(N23616,R2,R3);
and and14305(N23622,N23626,in0);
and and14306(N23623,in2,R0);
and and14307(N23624,R1,R2);
and and14308(N23625,N23627,R5);
and and14313(N23631,N23635,in0);
and and14314(N23632,in1,R0);
and and14315(N23633,R1,R3);
and and14316(N23634,R4,R5);
and and14321(N23639,in0,N23643);
and and14322(N23640,N23644,N23645);
and and14323(N23641,N23646,N23647);
and and14324(N23642,N23648,N23649);
and and14328(N23653,N23657,N23658);
and and14329(N23654,N23659,N23660);
and and14330(N23655,R3,N23661);
and and14331(N23656,N23662,N23663);
and and14335(N23667,N23671,N23672);
and and14336(N23668,N23673,R3);
and and14337(N23669,N23674,N23675);
and and14338(N23670,N23676,R7);
and and14342(N23680,in0,N23684);
and and14343(N23681,N23685,N23686);
and and14344(N23682,N23687,N23688);
and and14345(N23683,N23689,R7);
and and14349(N23693,in0,N23697);
and and14350(N23694,N23698,N23699);
and and14351(N23695,N23700,N23701);
and and14352(N23696,R6,N23702);
and and14356(N23706,N23710,R0);
and and14357(N23707,R1,N23711);
and and14358(N23708,N23712,N23713);
and and14359(N23709,N23714,N23715);
and and14363(N23719,in0,N23723);
and and14364(N23720,N23724,R2);
and and14365(N23721,N23725,N23726);
and and14366(N23722,N23727,N23728);
and and14370(N23732,in0,N23736);
and and14371(N23733,N23737,N23738);
and and14372(N23734,R3,N23739);
and and14373(N23735,N23740,N23741);
and and14377(N23745,in0,N23749);
and and14378(N23746,R2,R3);
and and14379(N23747,N23750,N23751);
and and14380(N23748,N23752,N23753);
and and14384(N23757,in0,N23761);
and and14385(N23758,N23762,R2);
and and14386(N23759,N23763,N23764);
and and14387(N23760,R6,N23765);
and and14391(N23769,in0,N23773);
and and14392(N23770,N23774,N23775);
and and14393(N23771,R3,N23776);
and and14394(N23772,R5,N23777);
and and14398(N23781,in0,N23785);
and and14399(N23782,in2,N23786);
and and14400(N23783,R4,N23787);
and and14401(N23784,N23788,N23789);
and and14405(N23793,N23797,N23798);
and and14406(N23794,N23799,R3);
and and14407(N23795,N23800,R5);
and and14408(N23796,R6,N23801);
and and14412(N23805,N23809,N23810);
and and14413(N23806,R1,R2);
and and14414(N23807,N23811,N23812);
and and14415(N23808,N23813,R7);
and and14419(N23817,N23821,N23822);
and and14420(N23818,R1,R2);
and and14421(N23819,N23823,R5);
and and14422(N23820,N23824,N23825);
and and14426(N23829,R0,N23833);
and and14427(N23830,N23834,N23835);
and and14428(N23831,R4,R5);
and and14429(N23832,N23836,N23837);
and and14433(N23841,in0,in1);
and and14434(N23842,N23845,N23846);
and and14435(N23843,R3,N23847);
and and14436(N23844,N23848,N23849);
and and14440(N23853,N23857,in1);
and and14441(N23854,N23858,R0);
and and14442(N23855,R3,N23859);
and and14443(N23856,N23860,R7);
and and14447(N23864,in0,in1);
and and14448(N23865,in2,N23868);
and and14449(N23866,N23869,N23870);
and and14450(N23867,R6,N23871);
and and14454(N23875,N23879,N23880);
and and14455(N23876,N23881,R2);
and and14456(N23877,R3,R4);
and and14457(N23878,R5,N23882);
and and14461(N23886,in1,N23890);
and and14462(N23887,N23891,R1);
and and14463(N23888,R2,N23892);
and and14464(N23889,N23893,R6);
and and14468(N23897,in0,N23901);
and and14469(N23898,N23902,R1);
and and14470(N23899,R2,N23903);
and and14471(N23900,N23904,R6);
and and14475(N23908,in0,R0);
and and14476(N23909,R1,N23912);
and and14477(N23910,N23913,N23914);
and and14478(N23911,R6,N23915);
and and14482(N23919,in1,N23923);
and and14483(N23920,N23924,R3);
and and14484(N23921,N23925,R5);
and and14485(N23922,R6,N23926);
and and14489(N23930,in0,N23934);
and and14490(N23931,R1,R2);
and and14491(N23932,N23935,R5);
and and14492(N23933,N23936,N23937);
and and14496(N23941,in0,R0);
and and14497(N23942,R1,N23945);
and and14498(N23943,R3,N23946);
and and14499(N23944,N23947,R7);
and and14503(N23951,in0,N23955);
and and14504(N23952,N23956,R2);
and and14505(N23953,R3,R5);
and and14506(N23954,R6,N23957);
and and14510(N23961,in0,N23965);
and and14511(N23962,R0,N23966);
and and14512(N23963,R2,R3);
and and14513(N23964,R5,N23967);
and and14517(N23971,in2,N23975);
and and14518(N23972,R1,R3);
and and14519(N23973,R4,N23976);
and and14520(N23974,N23977,R7);
and and14524(N23981,R0,N23985);
and and14525(N23982,R2,N23986);
and and14526(N23983,R4,N23987);
and and14527(N23984,R6,R7);
and and14531(N23991,in0,R0);
and and14532(N23992,R1,N23995);
and and14533(N23993,N23996,N23997);
and and14534(N23994,R6,R7);
and and14538(N24001,in0,in2);
and and14539(N24002,R0,N24005);
and and14540(N24003,R2,N24006);
and and14541(N24004,R5,N24007);
and and14545(N24011,in0,in2);
and and14546(N24012,R0,N24015);
and and14547(N24013,R2,N24016);
and and14548(N24014,R4,N24017);
and and14552(N24021,in0,N24025);
and and14553(N24022,R0,R1);
and and14554(N24023,N24026,R3);
and and14555(N24024,N24027,R7);
and and14559(N24031,in1,N24035);
and and14560(N24032,N24036,R2);
and and14561(N24033,R3,R4);
and and14562(N24034,R5,N24037);
and and14566(N24041,N24045,N24046);
and and14567(N24042,R2,R3);
and and14568(N24043,R4,R5);
and and14569(N24044,R6,R7);
and and14573(N24050,in0,R0);
and and14574(N24051,R2,N24054);
and and14575(N24052,R4,N24055);
and and14576(N24053,R6,R7);
and and10683(N18117,N18124,N18125);
and and10684(N18118,N18126,N18127);
and and10692(N18135,N18142,R5);
and and10693(N18136,N18143,N18144);
and and10701(N18152,N18159,N18160);
and and10702(N18153,N18161,R7);
and and10710(N18169,N18176,N18177);
and and10711(N18170,N18178,R7);
and and10719(N18186,N18193,N18194);
and and10720(N18187,R6,N18195);
and and10728(N18203,R3,R5);
and and10729(N18204,N18211,N18212);
and and10737(N18220,N18227,N18228);
and and10738(N18221,N18229,R7);
and and10746(N18237,N18242,N18243);
and and10747(N18238,N18244,N18245);
and and10755(N18253,R4,R5);
and and10756(N18254,N18260,N18261);
and and10764(N18269,R4,N18275);
and and10765(N18270,N18276,N18277);
and and10773(N18285,R4,N18291);
and and10774(N18286,N18292,N18293);
and and10782(N18301,R4,N18307);
and and10783(N18302,N18308,N18309);
and and10791(N18317,N18323,N18324);
and and10792(N18318,N18325,R7);
and and10800(N18333,R4,N18339);
and and10801(N18334,N18340,N18341);
and and10809(N18349,N18355,R4);
and and10810(N18350,N18356,N18357);
and and10818(N18365,N18372,N18373);
and and10819(N18366,R6,R7);
and and10827(N18381,N18387,N18388);
and and10828(N18382,R6,N18389);
and and10836(N18397,N18402,N18403);
and and10837(N18398,N18404,N18405);
and and10845(N18413,N18418,N18419);
and and10846(N18414,N18420,N18421);
and and10854(N18429,R4,N18435);
and and10855(N18430,N18436,N18437);
and and10863(N18445,N18451,R5);
and and10864(N18446,N18452,N18453);
and and10872(N18461,N18467,R5);
and and10873(N18462,N18468,N18469);
and and10881(N18477,N18483,N18484);
and and10882(N18478,N18485,R7);
and and10890(N18493,N18499,R4);
and and10891(N18494,N18500,N18501);
and and10899(N18509,N18515,N18516);
and and10900(N18510,N18517,R7);
and and10908(N18525,N18531,N18532);
and and10909(N18526,N18533,R7);
and and10917(N18541,R4,N18548);
and and10918(N18542,N18549,R7);
and and10926(N18557,N18563,R5);
and and10927(N18558,R6,N18564);
and and10935(N18572,N18576,N18577);
and and10936(N18573,N18578,N18579);
and and10944(N18587,N18592,N18593);
and and10945(N18588,R6,N18594);
and and10953(N18602,N18606,N18607);
and and10954(N18603,N18608,N18609);
and and10962(N18617,N18623,R5);
and and10963(N18618,R6,N18624);
and and10971(N18632,N18637,N18638);
and and10972(N18633,R6,N18639);
and and10980(N18647,N18652,R5);
and and10981(N18648,N18653,N18654);
and and10989(N18662,N18667,R5);
and and10990(N18663,N18668,N18669);
and and10998(N18677,N18683,R5);
and and10999(N18678,R6,N18684);
and and11007(N18692,N18697,R4);
and and11008(N18693,N18698,N18699);
and and11016(N18707,N18713,R5);
and and11017(N18708,R6,N18714);
and and11025(N18722,N18728,N18729);
and and11026(N18723,R6,R7);
and and11034(N18737,N18741,N18742);
and and11035(N18738,N18743,N18744);
and and11043(N18752,N18756,N18757);
and and11044(N18753,N18758,N18759);
and and11052(N18767,N18771,N18772);
and and11053(N18768,N18773,N18774);
and and11061(N18782,R4,N18788);
and and11062(N18783,N18789,R7);
and and11070(N18797,R4,N18803);
and and11071(N18798,N18804,R7);
and and11079(N18812,N18818,R5);
and and11080(N18813,R6,N18819);
and and11088(N18827,N18832,R5);
and and11089(N18828,N18833,N18834);
and and11097(N18842,N18847,N18848);
and and11098(N18843,N18849,R7);
and and11106(N18857,R3,R5);
and and11107(N18858,N18863,N18864);
and and11115(N18872,N18877,N18878);
and and11116(N18873,R6,N18879);
and and11124(N18887,N18892,N18893);
and and11125(N18888,N18894,R7);
and and11133(N18902,R4,R5);
and and11134(N18903,N18908,N18909);
and and11142(N18917,R4,N18921);
and and11143(N18918,N18922,N18923);
and and11151(N18931,R4,N18935);
and and11152(N18932,N18936,N18937);
and and11160(N18945,N18949,N18950);
and and11161(N18946,R6,N18951);
and and11169(N18959,N18963,R5);
and and11170(N18960,N18964,N18965);
and and11178(N18973,R4,N18977);
and and11179(N18974,N18978,N18979);
and and11187(N18987,R4,R5);
and and11188(N18988,N18992,N18993);
and and11196(N19001,R4,R5);
and and11197(N19002,N19006,N19007);
and and11205(N19015,N19019,R5);
and and11206(N19016,N19020,N19021);
and and11214(N19029,R3,N19034);
and and11215(N19030,R5,N19035);
and and11223(N19043,R4,N19048);
and and11224(N19044,N19049,R7);
and and11232(N19057,R4,N19062);
and and11233(N19058,N19063,R7);
and and11241(N19071,R4,R5);
and and11242(N19072,N19076,N19077);
and and11250(N19085,R4,R5);
and and11251(N19086,N19090,N19091);
and and11259(N19099,R3,R4);
and and11260(N19100,N19105,R7);
and and11268(N19113,N19118,R5);
and and11269(N19114,R6,N19119);
and and11277(N19127,R4,R5);
and and11278(N19128,N19132,N19133);
and and11286(N19141,N19146,R5);
and and11287(N19142,N19147,R7);
and and11295(N19155,R4,R5);
and and11296(N19156,N19161,R7);
and and11304(N19169,N19173,R5);
and and11305(N19170,N19174,N19175);
and and11313(N19183,N19187,R5);
and and11314(N19184,N19188,N19189);
and and11322(N19197,R4,N19201);
and and11323(N19198,N19202,N19203);
and and11331(N19211,R4,R5);
and and11332(N19212,R6,N19217);
and and11340(N19225,N19230,N19231);
and and11341(N19226,R6,R7);
and and11349(N19239,N19244,N19245);
and and11350(N19240,R6,R7);
and and11358(N19253,N19258,N19259);
and and11359(N19254,R6,R7);
and and11367(N19267,N19272,R5);
and and11368(N19268,N19273,R7);
and and11376(N19281,N19286,R5);
and and11377(N19282,N19287,R7);
and and11385(N19295,N19300,R5);
and and11386(N19296,N19301,R7);
and and11394(N19309,R4,R5);
and and11395(N19310,N19315,R7);
and and11403(N19323,N19328,R5);
and and11404(N19324,N19329,R7);
and and11412(N19337,R4,N19342);
and and11413(N19338,N19343,R7);
and and11421(N19351,R4,N19356);
and and11422(N19352,R6,N19357);
and and11430(N19365,R4,N19369);
and and11431(N19366,N19370,N19371);
and and11439(N19379,R3,N19384);
and and11440(N19380,R5,N19385);
and and11448(N19393,R4,N19398);
and and11449(N19394,R6,N19399);
and and11457(N19407,R4,R5);
and and11458(N19408,R6,N19413);
and and11466(N19421,R4,N19427);
and and11467(N19422,R6,R7);
and and11475(N19435,R4,N19441);
and and11476(N19436,R6,R7);
and and11484(N19449,N19453,N19454);
and and11485(N19450,N19455,R7);
and and11493(N19463,N19467,N19468);
and and11494(N19464,N19469,R7);
and and11502(N19477,R3,N19482);
and and11503(N19478,R5,N19483);
and and11511(N19491,N19495,R5);
and and11512(N19492,N19496,N19497);
and and11520(N19505,R4,N19510);
and and11521(N19506,N19511,R7);
and and11529(N19519,R4,N19524);
and and11530(N19520,N19525,R7);
and and11538(N19533,N19538,R4);
and and11539(N19534,R5,N19539);
and and11547(N19547,R4,N19552);
and and11548(N19548,R6,N19553);
and and11556(N19561,R3,R4);
and and11557(N19562,R5,N19567);
and and11565(N19575,R4,R5);
and and11566(N19576,N19580,N19581);
and and11574(N19589,N19593,N19594);
and and11575(N19590,R5,N19595);
and and11583(N19603,N19608,N19609);
and and11584(N19604,R6,R7);
and and11592(N19617,R3,N19623);
and and11593(N19618,R5,R6);
and and11601(N19631,N19636,R4);
and and11602(N19632,N19637,R7);
and and11610(N19645,N19649,N19650);
and and11611(N19646,R5,N19651);
and and11619(N19659,N19663,R5);
and and11620(N19660,N19664,N19665);
and and11628(N19673,R3,R4);
and and11629(N19674,N19679,R7);
and and11637(N19687,R4,N19692);
and and11638(N19688,N19693,R7);
and and11646(N19701,R4,N19706);
and and11647(N19702,N19707,R7);
and and11655(N19715,R4,N19720);
and and11656(N19716,N19721,R7);
and and11664(N19729,N19733,N19734);
and and11665(N19730,R6,R7);
and and11673(N19742,R4,N19745);
and and11674(N19743,N19746,N19747);
and and11682(N19755,R3,R4);
and and11683(N19756,N19759,N19760);
and and11691(N19768,R4,R5);
and and11692(N19769,R6,R7);
and and11700(N19781,N19785,R5);
and and11701(N19782,N19786,R7);
and and11709(N19794,R3,R4);
and and11710(N19795,N19798,N19799);
and and11718(N19807,N19810,N19811);
and and11719(N19808,R6,N19812);
and and11727(N19820,R3,N19824);
and and11728(N19821,R6,N19825);
and and11736(N19833,R3,N19837);
and and11737(N19834,N19838,R6);
and and11745(N19846,R3,R5);
and and11746(N19847,R6,N19851);
and and11754(N19859,N19862,N19863);
and and11755(N19860,R6,N19864);
and and11763(N19872,R4,R5);
and and11764(N19873,R6,N19877);
and and11772(N19885,R4,R5);
and and11773(N19886,N19890,R7);
and and11781(N19898,R4,R5);
and and11782(N19899,N19903,R7);
and and11790(N19911,R4,R5);
and and11791(N19912,N19915,N19916);
and and11799(N19924,R4,R5);
and and11800(N19925,N19928,N19929);
and and11808(N19937,N19941,R5);
and and11809(N19938,R6,N19942);
and and11817(N19950,R4,R5);
and and11818(N19951,R6,N19955);
and and11826(N19963,N19968,R5);
and and11827(N19964,R6,R7);
and and11835(N19976,R4,R5);
and and11836(N19977,R6,N19981);
and and11844(N19989,R4,N19993);
and and11845(N19990,R6,N19994);
and and11853(N20002,R3,R4);
and and11854(N20003,N20007,R7);
and and11862(N20015,R4,N20020);
and and11863(N20016,R6,R7);
and and11871(N20028,R3,R4);
and and11872(N20029,N20032,N20033);
and and11880(N20041,R4,N20045);
and and11881(N20042,R6,N20046);
and and11889(N20054,R4,N20058);
and and11890(N20055,R6,N20059);
and and11898(N20067,R4,N20071);
and and11899(N20068,R6,N20072);
and and11907(N20080,R4,N20084);
and and11908(N20081,R6,N20085);
and and11916(N20093,N20098,R5);
and and11917(N20094,R6,R7);
and and11925(N20106,N20110,N20111);
and and11926(N20107,R6,R7);
and and11934(N20119,R4,R5);
and and11935(N20120,N20124,R7);
and and11943(N20132,R4,R5);
and and11944(N20133,N20137,R7);
and and11952(N20145,R3,R5);
and and11953(N20146,N20149,N20150);
and and11961(N20158,R4,N20163);
and and11962(N20159,R6,R7);
and and11970(N20171,R3,R4);
and and11971(N20172,R6,N20176);
and and11979(N20184,R4,R5);
and and11980(N20185,N20188,N20189);
and and11988(N20197,R4,R5);
and and11989(N20198,N20201,N20202);
and and11997(N20210,R4,R5);
and and11998(N20211,N20214,N20215);
and and12006(N20223,N20228,R4);
and and12007(N20224,R6,R7);
and and12015(N20236,R4,N20240);
and and12016(N20237,N20241,R7);
and and12024(N20249,N20252,R5);
and and12025(N20250,R6,N20253);
and and12033(N20261,R4,R5);
and and12034(N20262,N20264,N20265);
and and12042(N20273,R3,R5);
and and12043(N20274,N20277,R7);
and and12051(N20285,R3,R5);
and and12052(N20286,N20289,R7);
and and12060(N20297,R4,N20300);
and and12061(N20298,N20301,R7);
and and12069(N20309,R4,N20313);
and and12070(N20310,R6,R7);
and and12078(N20321,R4,N20324);
and and12079(N20322,R6,N20325);
and and12087(N20333,N20336,R5);
and and12088(N20334,N20337,R7);
and and12096(N20345,R4,R5);
and and12097(N20346,R6,N20349);
and and12105(N20357,N20360,N20361);
and and12106(N20358,R6,R7);
and and12114(N20369,R4,R5);
and and12115(N20370,N20373,R7);
and and12123(N20381,R4,R5);
and and12124(N20382,N20384,N20385);
and and12132(N20393,N20395,N20396);
and and12133(N20394,R6,N20397);
and and12141(N20405,N20408,R5);
and and12142(N20406,R6,N20409);
and and12150(N20417,R3,N20421);
and and12151(N20418,R5,R7);
and and12159(N20429,N20433,R5);
and and12160(N20430,R6,R7);
and and12168(N20441,R4,R5);
and and12169(N20442,N20444,N20445);
and and12177(N20453,N20455,R5);
and and12178(N20454,N20456,N20457);
and and12186(N20465,R3,N20468);
and and12187(N20466,R5,N20469);
and and12195(N20477,N20481,R5);
and and12196(N20478,R6,R7);
and and12204(N20489,R3,R5);
and and12205(N20490,R6,R7);
and and12213(N20501,N20504,N20505);
and and12214(N20502,R6,R7);
and and12222(N20513,R4,N20516);
and and12223(N20514,N20517,R7);
and and12231(N20525,R4,R5);
and and12232(N20526,R6,R7);
and and12240(N20537,R4,N20541);
and and12241(N20538,R6,R7);
and and12249(N20549,R4,N20553);
and and12250(N20550,R6,R7);
and and12258(N20561,R4,R5);
and and12259(N20562,N20565,R7);
and and12267(N20573,R3,R4);
and and12268(N20574,R5,R7);
and and12276(N20585,R4,R5);
and and12277(N20586,R6,N20589);
and and12285(N20597,R4,R5);
and and12286(N20598,N20601,R7);
and and12294(N20609,R3,R4);
and and12295(N20610,N20613,R6);
and and12303(N20621,R4,R5);
and and12304(N20622,N20624,N20625);
and and12312(N20633,N20636,N20637);
and and12313(N20634,R6,R7);
and and12321(N20645,R4,R5);
and and12322(N20646,N20648,N20649);
and and12330(N20657,R4,N20660);
and and12331(N20658,N20661,R7);
and and12339(N20669,N20671,N20672);
and and12340(N20670,R6,R7);
and and12348(N20680,R4,R5);
and and12349(N20681,R6,N20683);
and and12357(N20691,R3,R4);
and and12358(N20692,N20694,R6);
and and12366(N20702,R4,N20705);
and and12367(N20703,R6,R7);
and and12375(N20713,R3,R4);
and and12376(N20714,R6,R7);
and and12384(N20724,N20727,R4);
and and12385(N20725,R6,R7);
and and12393(N20735,N20737,R4);
and and12394(N20736,R5,R7);
and and12402(N20745,R4,R5);
and and12403(N20746,R6,R7);
and and12411(N20755,R4,R5);
and and12412(N20756,R6,R7);
and and12420(N20765,R3,N20767);
and and12421(N20766,R5,R7);
and and12429(N20775,R4,R5);
and and12430(N20776,R6,R7);
and and12438(N20785,R4,R5);
and and12439(N20786,R6,N20787);
and and12447(N20795,R3,R4);
and and12448(N20796,R5,N20797);
and and12456(N20805,R4,R5);
and and12457(N20806,R6,N20807);
and and12465(N20815,R4,R5);
and and12466(N20816,N20817,R7);
and and12474(N20825,R4,R5);
and and12475(N20826,R6,R7);
and and12483(N20835,R4,N20837);
and and12484(N20836,R6,R7);
and and12492(N20845,R3,R4);
and and12493(N20846,R5,R7);
and and12501(N20855,N20862,N20863);
and and12509(N20871,N20878,N20879);
and and12517(N20887,N20893,N20894);
and and12525(N20902,R6,N20909);
and and12533(N20917,N20923,N20924);
and and12541(N20932,R6,N20939);
and and12549(N20947,R6,N20954);
and and12557(N20962,N20968,N20969);
and and12565(N20977,N20983,N20984);
and and12573(N20992,N20998,N20999);
and and12581(N21007,N21013,N21014);
and and12589(N21022,N21028,N21029);
and and12597(N21037,N21043,N21044);
and and12605(N21052,R6,N21059);
and and12613(N21067,N21073,N21074);
and and12621(N21082,N21087,N21088);
and and12629(N21096,N21101,N21102);
and and12637(N21110,N21115,N21116);
and and12645(N21124,N21129,N21130);
and and12653(N21138,N21144,R7);
and and12661(N21152,N21158,R7);
and and12669(N21166,N21171,N21172);
and and12677(N21180,N21185,N21186);
and and12685(N21194,R6,N21200);
and and12693(N21208,R6,N21214);
and and12701(N21222,N21228,R7);
and and12709(N21236,N21242,R7);
and and12717(N21250,R6,N21256);
and and12725(N21264,N21269,N21270);
and and12733(N21278,N21283,N21284);
and and12741(N21292,N21297,N21298);
and and12749(N21306,N21311,N21312);
and and12757(N21320,N21326,R7);
and and12765(N21334,R6,N21340);
and and12773(N21348,N21353,N21354);
and and12781(N21362,N21367,N21368);
and and12789(N21376,N21381,N21382);
and and12797(N21390,R5,N21396);
and and12805(N21404,N21409,N21410);
and and12813(N21418,R6,N21424);
and and12821(N21432,N21438,R7);
and and12829(N21446,R6,N21452);
and and12837(N21460,N21465,N21466);
and and12845(N21474,N21479,N21480);
and and12853(N21488,N21493,N21494);
and and12861(N21502,R6,N21508);
and and12869(N21516,N21521,N21522);
and and12877(N21530,N21534,N21535);
and and12885(N21543,N21548,R7);
and and12893(N21556,N21560,N21561);
and and12901(N21569,R6,N21574);
and and12909(N21582,N21586,N21587);
and and12917(N21595,R6,N21600);
and and12925(N21608,R6,N21613);
and and12933(N21621,R6,N21626);
and and12941(N21634,N21639,R6);
and and12949(N21647,N21652,R7);
and and12957(N21660,N21664,N21665);
and and12965(N21673,N21677,N21678);
and and12973(N21686,R6,R7);
and and12981(N21699,R6,R7);
and and12989(N21712,R6,R7);
and and12997(N21725,N21730,R7);
and and13005(N21738,N21743,R7);
and and13013(N21751,R6,N21756);
and and13021(N21764,R6,N21769);
and and13029(N21777,R6,N21782);
and and13037(N21790,R6,N21795);
and and13045(N21803,N21807,N21808);
and and13053(N21816,R6,N21821);
and and13061(N21829,R6,N21834);
and and13069(N21842,R6,R7);
and and13077(N21855,R6,N21860);
and and13085(N21868,N21872,N21873);
and and13093(N21881,N21886,R7);
and and13101(N21894,N21899,R7);
and and13109(N21907,N21912,R7);
and and13117(N21920,N21925,R7);
and and13125(N21933,R6,R7);
and and13133(N21946,R6,R7);
and and13141(N21959,N21964,R6);
and and13149(N21972,N21977,R6);
and and13157(N21985,N21990,R7);
and and13165(N21998,N22003,R7);
and and13173(N22011,N22016,R7);
and and13181(N22024,N22029,R7);
and and13189(N22037,N22042,R7);
and and13197(N22050,N22055,R7);
and and13205(N22063,N22067,N22068);
and and13213(N22076,N22081,R7);
and and13221(N22089,N22094,R7);
and and13229(N22102,N22106,N22107);
and and13237(N22115,N22120,R7);
and and13245(N22128,N22132,N22133);
and and13253(N22141,N22146,R6);
and and13261(N22154,N22159,R7);
and and13269(N22167,N22171,N22172);
and and13277(N22180,R6,N22185);
and and13285(N22193,N22198,R7);
and and13293(N22206,N22211,R6);
and and13301(N22219,N22223,N22224);
and and13309(N22232,N22236,R7);
and and13317(N22244,N22247,N22248);
and and13325(N22256,N22259,N22260);
and and13333(N22268,R6,R7);
and and13341(N22280,R6,N22284);
and and13349(N22292,R6,N22296);
and and13357(N22304,N22307,N22308);
and and13365(N22316,N22319,N22320);
and and13373(N22328,N22332,R6);
and and13381(N22340,R5,N22344);
and and13389(N22352,R4,N22356);
and and13397(N22364,N22368,R7);
and and13405(N22376,R6,N22380);
and and13413(N22388,R6,N22392);
and and13421(N22400,R6,R7);
and and13429(N22412,N22416,R7);
and and13437(N22424,R6,N22428);
and and13445(N22436,R5,N22440);
and and13453(N22448,R6,N22452);
and and13461(N22460,N22464,R7);
and and13469(N22472,N22476,R7);
and and13477(N22484,N22488,R7);
and and13485(N22496,N22500,R7);
and and13493(N22508,R6,R7);
and and13501(N22520,N22524,R6);
and and13509(N22532,R6,N22536);
and and13517(N22544,N22548,R7);
and and13525(N22556,N22560,R7);
and and13533(N22568,R5,N22572);
and and13541(N22580,N22584,R7);
and and13549(N22592,R6,N22596);
and and13557(N22604,R6,N22608);
and and13565(N22616,R5,N22620);
and and13573(N22628,R5,N22632);
and and13581(N22640,R6,N22644);
and and13589(N22652,N22655,N22656);
and and13597(N22664,N22668,R7);
and and13605(N22676,N22680,R7);
and and13613(N22688,N22692,R7);
and and13621(N22700,R6,R7);
and and13629(N22712,N22716,R7);
and and13637(N22724,R6,N22728);
and and13645(N22736,R6,N22740);
and and13653(N22748,R6,R7);
and and13661(N22760,R6,R7);
and and13669(N22772,R6,N22776);
and and13677(N22784,R6,R7);
and and13685(N22796,R6,N22800);
and and13693(N22808,N22812,R7);
and and13701(N22820,N22823,N22824);
and and13709(N22832,N22834,N22835);
and and13717(N22843,N22845,N22846);
and and13725(N22854,R6,N22857);
and and13733(N22865,R6,N22868);
and and13741(N22876,R6,R7);
and and13749(N22887,R6,N22890);
and and13757(N22898,R6,R7);
and and13765(N22909,N22912,R7);
and and13773(N22920,R6,N22923);
and and13781(N22931,R6,N22934);
and and13789(N22942,R6,N22945);
and and13797(N22953,R6,N22956);
and and13805(N22964,R6,R7);
and and13813(N22975,R6,R7);
and and13821(N22986,R5,N22989);
and and13829(N22997,R6,R7);
and and13837(N23008,R6,N23011);
and and13845(N23019,R6,N23022);
and and13853(N23030,R6,N23033);
and and13861(N23041,R6,R7);
and and13869(N23052,N23055,R7);
and and13877(N23063,N23066,R7);
and and13885(N23074,N23077,R7);
and and13893(N23085,N23088,R7);
and and13901(N23096,R6,R7);
and and13909(N23107,N23110,R7);
and and13917(N23118,N23121,R7);
and and13925(N23129,N23132,R7);
and and13933(N23140,N23143,R7);
and and13941(N23151,N23154,R7);
and and13949(N23162,R4,R6);
and and13957(N23173,R5,N23176);
and and13965(N23184,N23186,N23187);
and and13973(N23195,R6,N23198);
and and13981(N23206,R6,N23209);
and and13989(N23217,N23220,R7);
and and13997(N23228,N23230,N23231);
and and14005(N23239,N23242,R7);
and and14013(N23250,N23252,N23253);
and and14021(N23261,R6,R7);
and and14029(N23272,R6,R7);
and and14037(N23283,R4,R6);
and and14045(N23294,R6,N23297);
and and14053(N23305,R6,N23308);
and and14061(N23316,R6,N23319);
and and14069(N23327,N23330,R7);
and and14077(N23338,N23341,R7);
and and14085(N23349,R6,N23352);
and and14093(N23360,R5,N23363);
and and14101(N23371,N23374,R6);
and and14109(N23382,R5,N23385);
and and14117(N23393,R6,N23396);
and and14125(N23404,N23406,R7);
and and14133(N23414,N23416,R7);
and and14141(N23424,N23426,R7);
and and14149(N23434,N23436,R7);
and and14157(N23444,N23446,R7);
and and14165(N23454,R6,R7);
and and14173(N23464,R6,R7);
and and14181(N23474,R6,R7);
and and14189(N23484,R6,R7);
and and14197(N23494,R6,R7);
and and14205(N23504,R6,R7);
and and14213(N23514,R6,N23516);
and and14221(N23524,R6,R7);
and and14229(N23534,R6,R7);
and and14237(N23544,N23546,R7);
and and14245(N23554,R5,R6);
and and14253(N23563,R6,R7);
and and14261(N23572,R5,R6);
and and14269(N23581,R6,N23582);
and and14277(N23590,R6,R7);
and and14285(N23599,R6,N23600);
and and14293(N23608,N23609,R7);
and and14301(N23617,R4,R7);
and and14309(N23626,R6,R7);
and and14317(N23635,R6,R7);
and and14577(N24427,N24428,N24429);
and and14586(N24444,N24445,N24446);
and and14595(N24461,N24462,N24463);
and and14604(N24478,N24479,N24480);
and and14613(N24495,N24496,N24497);
and and14622(N24512,N24513,N24514);
and and14631(N24529,N24530,N24531);
and and14640(N24546,N24547,N24548);
and and14649(N24563,N24564,N24565);
and and14658(N24579,N24580,N24581);
and and14667(N24595,N24596,N24597);
and and14676(N24611,N24612,N24613);
and and14685(N24627,N24628,N24629);
and and14694(N24643,N24644,N24645);
and and14703(N24659,N24660,N24661);
and and14712(N24675,N24676,N24677);
and and14721(N24691,N24692,N24693);
and and14730(N24707,N24708,N24709);
and and14739(N24723,N24724,N24725);
and and14748(N24739,N24740,N24741);
and and14757(N24755,N24756,N24757);
and and14766(N24771,N24772,N24773);
and and14775(N24787,N24788,N24789);
and and14784(N24803,N24804,N24805);
and and14793(N24819,N24820,N24821);
and and14802(N24835,N24836,N24837);
and and14811(N24851,N24852,N24853);
and and14820(N24867,N24868,N24869);
and and14829(N24882,N24883,N24884);
and and14838(N24897,N24898,N24899);
and and14847(N24912,N24913,N24914);
and and14856(N24927,N24928,N24929);
and and14865(N24942,N24943,N24944);
and and14874(N24957,N24958,N24959);
and and14883(N24972,N24973,N24974);
and and14892(N24987,N24988,N24989);
and and14901(N25002,N25003,N25004);
and and14910(N25017,N25018,N25019);
and and14919(N25032,N25033,N25034);
and and14928(N25047,N25048,N25049);
and and14937(N25062,N25063,N25064);
and and14946(N25077,N25078,N25079);
and and14955(N25092,N25093,N25094);
and and14964(N25107,N25108,N25109);
and and14973(N25122,N25123,N25124);
and and14982(N25137,N25138,N25139);
and and14991(N25152,N25153,N25154);
and and15000(N25167,N25168,N25169);
and and15009(N25182,N25183,N25184);
and and15018(N25197,N25198,N25199);
and and15027(N25212,N25213,N25214);
and and15036(N25227,N25228,N25229);
and and15045(N25242,N25243,N25244);
and and15054(N25257,N25258,N25259);
and and15063(N25271,N25272,N25273);
and and15072(N25285,N25286,N25287);
and and15081(N25299,N25300,N25301);
and and15090(N25313,N25314,N25315);
and and15099(N25327,N25328,N25329);
and and15108(N25341,N25342,N25343);
and and15117(N25355,N25356,N25357);
and and15126(N25369,N25370,N25371);
and and15135(N25383,N25384,N25385);
and and15144(N25397,N25398,N25399);
and and15153(N25411,N25412,N25413);
and and15162(N25425,N25426,N25427);
and and15171(N25439,N25440,N25441);
and and15180(N25453,N25454,N25455);
and and15189(N25467,N25468,N25469);
and and15198(N25481,N25482,N25483);
and and15207(N25495,N25496,N25497);
and and15216(N25509,N25510,N25511);
and and15225(N25523,N25524,N25525);
and and15234(N25537,N25538,N25539);
and and15243(N25551,N25552,N25553);
and and15252(N25565,N25566,N25567);
and and15261(N25579,N25580,N25581);
and and15270(N25593,N25594,N25595);
and and15279(N25607,N25608,N25609);
and and15288(N25621,N25622,N25623);
and and15297(N25635,N25636,N25637);
and and15306(N25649,N25650,N25651);
and and15315(N25663,N25664,N25665);
and and15324(N25677,N25678,N25679);
and and15333(N25691,N25692,N25693);
and and15342(N25705,N25706,N25707);
and and15351(N25719,N25720,N25721);
and and15360(N25733,N25734,N25735);
and and15369(N25747,N25748,N25749);
and and15378(N25761,N25762,N25763);
and and15387(N25775,N25776,N25777);
and and15396(N25789,N25790,N25791);
and and15405(N25803,N25804,N25805);
and and15414(N25817,N25818,N25819);
and and15423(N25831,N25832,N25833);
and and15432(N25845,N25846,N25847);
and and15441(N25859,N25860,N25861);
and and15450(N25873,N25874,N25875);
and and15459(N25887,N25888,N25889);
and and15468(N25901,N25902,N25903);
and and15477(N25915,N25916,N25917);
and and15486(N25929,N25930,N25931);
and and15495(N25943,N25944,N25945);
and and15504(N25957,N25958,N25959);
and and15513(N25971,N25972,N25973);
and and15522(N25985,N25986,N25987);
and and15531(N25999,N26000,N26001);
and and15540(N26013,N26014,N26015);
and and15549(N26027,N26028,N26029);
and and15558(N26041,N26042,N26043);
and and15567(N26055,N26056,N26057);
and and15576(N26069,N26070,N26071);
and and15585(N26083,N26084,N26085);
and and15594(N26097,N26098,N26099);
and and15603(N26111,N26112,N26113);
and and15612(N26125,N26126,N26127);
and and15621(N26139,N26140,N26141);
and and15630(N26152,N26153,N26154);
and and15639(N26165,N26166,N26167);
and and15648(N26178,N26179,N26180);
and and15657(N26191,N26192,N26193);
and and15666(N26204,N26205,N26206);
and and15675(N26217,N26218,N26219);
and and15684(N26230,N26231,N26232);
and and15693(N26243,N26244,N26245);
and and15702(N26256,N26257,N26258);
and and15711(N26269,N26270,N26271);
and and15720(N26282,N26283,N26284);
and and15729(N26295,N26296,N26297);
and and15738(N26308,N26309,N26310);
and and15747(N26321,N26322,N26323);
and and15756(N26334,N26335,N26336);
and and15765(N26347,N26348,N26349);
and and15774(N26360,N26361,N26362);
and and15783(N26373,N26374,N26375);
and and15792(N26386,N26387,N26388);
and and15801(N26399,N26400,N26401);
and and15810(N26412,N26413,N26414);
and and15819(N26425,N26426,N26427);
and and15828(N26438,N26439,N26440);
and and15837(N26451,N26452,N26453);
and and15846(N26464,N26465,N26466);
and and15855(N26477,N26478,N26479);
and and15864(N26490,N26491,N26492);
and and15873(N26503,N26504,N26505);
and and15882(N26515,N26516,N26517);
and and15891(N26527,N26528,N26529);
and and15900(N26539,N26540,N26541);
and and15909(N26551,N26552,N26553);
and and15918(N26563,N26564,N26565);
and and15927(N26575,N26576,N26577);
and and15936(N26587,N26588,N26589);
and and15945(N26599,N26600,N26601);
and and15954(N26611,N26612,N26613);
and and15963(N26623,N26624,N26625);
and and15972(N26635,N26636,N26637);
and and15981(N26647,N26648,N26649);
and and15990(N26659,N26660,N26661);
and and15999(N26671,N26672,N26673);
and and16008(N26683,N26684,N26685);
and and16017(N26695,N26696,N26697);
and and16026(N26707,N26708,N26709);
and and16035(N26719,N26720,N26721);
and and16044(N26731,N26732,N26733);
and and16053(N26743,N26744,N26745);
and and16062(N26755,N26756,N26757);
and and16071(N26767,N26768,N26769);
and and16080(N26779,N26780,N26781);
and and16089(N26791,N26792,N26793);
and and16098(N26803,N26804,N26805);
and and16107(N26815,N26816,N26817);
and and16116(N26827,N26828,N26829);
and and16125(N26839,N26840,N26841);
and and16134(N26851,N26852,N26853);
and and16143(N26863,N26864,N26865);
and and16152(N26875,N26876,N26877);
and and16161(N26887,N26888,N26889);
and and16170(N26899,N26900,N26901);
and and16179(N26911,N26912,N26913);
and and16188(N26923,N26924,N26925);
and and16197(N26935,N26936,N26937);
and and16206(N26947,N26948,N26949);
and and16215(N26959,N26960,N26961);
and and16224(N26971,N26972,N26973);
and and16233(N26982,N26983,N26984);
and and16242(N26993,N26994,N26995);
and and16251(N27004,N27005,N27006);
and and16260(N27015,N27016,N27017);
and and16269(N27026,N27027,N27028);
and and16278(N27037,N27038,N27039);
and and16287(N27048,N27049,N27050);
and and16296(N27059,N27060,N27061);
and and16305(N27070,N27071,N27072);
and and16314(N27081,N27082,N27083);
and and16323(N27092,N27093,N27094);
and and16332(N27103,N27104,N27105);
and and16341(N27114,N27115,N27116);
and and16350(N27125,N27126,N27127);
and and16359(N27136,N27137,N27138);
and and16368(N27147,N27148,N27149);
and and16377(N27157,N27158,N27159);
and and16386(N27167,N27168,N27169);
and and16395(N27177,N27178,N27179);
and and16404(N27187,N27188,N27189);
and and16413(N27197,N27198,N27199);
and and16421(N27213,N27214,N27215);
and and16429(N27229,N27230,N27231);
and and16437(N27245,N27246,N27247);
and and16445(N27260,N27261,N27262);
and and16453(N27275,N27276,N27277);
and and16461(N27290,N27291,N27292);
and and16469(N27305,N27306,N27307);
and and16477(N27320,N27321,N27322);
and and16485(N27335,N27336,N27337);
and and16493(N27350,N27351,N27352);
and and16501(N27365,N27366,N27367);
and and16509(N27380,N27381,N27382);
and and16517(N27395,N27396,N27397);
and and16525(N27410,N27411,N27412);
and and16533(N27424,N27425,N27426);
and and16541(N27438,N27439,N27440);
and and16549(N27452,N27453,N27454);
and and16557(N27466,N27467,N27468);
and and16565(N27480,N27481,N27482);
and and16573(N27494,N27495,N27496);
and and16581(N27508,N27509,N27510);
and and16589(N27522,N27523,N27524);
and and16597(N27536,N27537,N27538);
and and16605(N27550,N27551,N27552);
and and16613(N27564,N27565,N27566);
and and16621(N27578,N27579,N27580);
and and16629(N27592,N27593,N27594);
and and16637(N27606,N27607,N27608);
and and16645(N27620,N27621,N27622);
and and16653(N27634,N27635,N27636);
and and16661(N27648,N27649,N27650);
and and16669(N27662,N27663,N27664);
and and16677(N27676,N27677,N27678);
and and16685(N27690,N27691,N27692);
and and16693(N27704,N27705,N27706);
and and16701(N27718,N27719,N27720);
and and16709(N27732,N27733,N27734);
and and16717(N27746,N27747,N27748);
and and16725(N27759,N27760,N27761);
and and16733(N27772,N27773,N27774);
and and16741(N27785,N27786,N27787);
and and16749(N27798,N27799,N27800);
and and16757(N27811,N27812,N27813);
and and16765(N27824,N27825,N27826);
and and16773(N27837,N27838,N27839);
and and16781(N27850,N27851,N27852);
and and16789(N27863,N27864,N27865);
and and16797(N27876,N27877,N27878);
and and16805(N27889,N27890,N27891);
and and16813(N27902,N27903,N27904);
and and16821(N27915,N27916,N27917);
and and16829(N27928,N27929,N27930);
and and16837(N27941,N27942,N27943);
and and16845(N27954,N27955,N27956);
and and16853(N27967,N27968,N27969);
and and16861(N27980,N27981,N27982);
and and16869(N27993,N27994,N27995);
and and16877(N28006,N28007,N28008);
and and16885(N28019,N28020,N28021);
and and16893(N28032,N28033,N28034);
and and16901(N28045,N28046,N28047);
and and16909(N28058,N28059,N28060);
and and16917(N28071,N28072,N28073);
and and16925(N28084,N28085,N28086);
and and16933(N28097,N28098,N28099);
and and16941(N28110,N28111,N28112);
and and16949(N28123,N28124,N28125);
and and16957(N28136,N28137,N28138);
and and16965(N28149,N28150,N28151);
and and16973(N28162,N28163,N28164);
and and16981(N28174,N28175,N28176);
and and16989(N28186,N28187,N28188);
and and16997(N28198,N28199,N28200);
and and17005(N28210,N28211,N28212);
and and17013(N28222,N28223,N28224);
and and17021(N28234,N28235,N28236);
and and17029(N28246,N28247,N28248);
and and17037(N28258,N28259,N28260);
and and17045(N28270,N28271,N28272);
and and17053(N28282,N28283,N28284);
and and17061(N28294,N28295,N28296);
and and17069(N28306,N28307,N28308);
and and17077(N28318,N28319,N28320);
and and17085(N28330,N28331,N28332);
and and17093(N28342,N28343,N28344);
and and17101(N28354,N28355,N28356);
and and17109(N28366,N28367,N28368);
and and17117(N28378,N28379,N28380);
and and17125(N28390,N28391,N28392);
and and17133(N28402,N28403,N28404);
and and17141(N28414,N28415,N28416);
and and17149(N28426,N28427,N28428);
and and17157(N28438,N28439,N28440);
and and17165(N28450,N28451,N28452);
and and17173(N28462,N28463,N28464);
and and17181(N28474,N28475,N28476);
and and17189(N28486,N28487,N28488);
and and17197(N28498,N28499,N28500);
and and17205(N28510,N28511,N28512);
and and17213(N28522,N28523,N28524);
and and17221(N28534,N28535,N28536);
and and17229(N28546,N28547,N28548);
and and17237(N28558,N28559,N28560);
and and17245(N28570,N28571,N28572);
and and17253(N28582,N28583,N28584);
and and17261(N28594,N28595,N28596);
and and17269(N28606,N28607,N28608);
and and17277(N28618,N28619,N28620);
and and17285(N28630,N28631,N28632);
and and17293(N28642,N28643,N28644);
and and17301(N28654,N28655,N28656);
and and17309(N28665,N28666,N28667);
and and17317(N28676,N28677,N28678);
and and17325(N28687,N28688,N28689);
and and17333(N28698,N28699,N28700);
and and17341(N28709,N28710,N28711);
and and17349(N28720,N28721,N28722);
and and17357(N28731,N28732,N28733);
and and17365(N28742,N28743,N28744);
and and17373(N28753,N28754,N28755);
and and17381(N28764,N28765,N28766);
and and17389(N28775,N28776,N28777);
and and17397(N28786,N28787,N28788);
and and17405(N28797,N28798,N28799);
and and17413(N28808,N28809,N28810);
and and17421(N28819,N28820,N28821);
and and17429(N28830,N28831,N28832);
and and17437(N28841,N28842,N28843);
and and17445(N28852,N28853,N28854);
and and17453(N28863,N28864,N28865);
and and17461(N28874,N28875,N28876);
and and17469(N28885,N28886,N28887);
and and17477(N28896,N28897,N28898);
and and17485(N28907,N28908,N28909);
and and17493(N28918,N28919,N28920);
and and17501(N28929,N28930,N28931);
and and17509(N28939,N28940,N28941);
and and17517(N28949,N28950,N28951);
and and17525(N28959,N28960,N28961);
and and17533(N28969,N28970,N28971);
and and17541(N28979,N28980,N28981);
and and17549(N28989,N28990,N28991);
and and17557(N28999,N29000,N29001);
and and17565(N29009,N29010,N29011);
and and17573(N29019,N29020,N29021);
and and17581(N29029,N29030,N29031);
and and17589(N29039,N29040,N29041);
and and17597(N29049,N29050,N29051);
and and17605(N29058,N29059,N29060);
and and17612(N29071,N29072,N29073);
and and17619(N29084,N29085,N29086);
and and17626(N29097,N29098,N29099);
and and17633(N29109,N29110,N29111);
and and17640(N29121,N29122,N29123);
and and17647(N29133,N29134,N29135);
and and17654(N29145,N29146,N29147);
and and17661(N29157,N29158,N29159);
and and17668(N29168,N29169,N29170);
and and17675(N29179,N29180,N29181);
and and17682(N29190,N29191,N29192);
and and17689(N29201,N29202,N29203);
and and17696(N29212,N29213,N29214);
and and17703(N29223,N29224,N29225);
and and17710(N29234,N29235,N29236);
and and17717(N29244,N29245,N29246);
and and17724(N29254,N29255,N29256);
and and17731(N29263,N29264,N29265);
and and14578(N24428,N24430,N24431);
and and14579(N24429,N24432,N24433);
and and14587(N24445,N24447,N24448);
and and14588(N24446,N24449,N24450);
and and14596(N24462,N24464,N24465);
and and14597(N24463,N24466,N24467);
and and14605(N24479,N24481,N24482);
and and14606(N24480,N24483,N24484);
and and14614(N24496,N24498,N24499);
and and14615(N24497,N24500,N24501);
and and14623(N24513,N24515,N24516);
and and14624(N24514,N24517,N24518);
and and14632(N24530,N24532,N24533);
and and14633(N24531,N24534,N24535);
and and14641(N24547,N24549,N24550);
and and14642(N24548,N24551,N24552);
and and14650(N24564,N24566,N24567);
and and14651(N24565,N24568,N24569);
and and14659(N24580,N24582,N24583);
and and14660(N24581,N24584,N24585);
and and14668(N24596,N24598,N24599);
and and14669(N24597,N24600,N24601);
and and14677(N24612,N24614,N24615);
and and14678(N24613,N24616,N24617);
and and14686(N24628,N24630,N24631);
and and14687(N24629,N24632,N24633);
and and14695(N24644,N24646,N24647);
and and14696(N24645,N24648,N24649);
and and14704(N24660,N24662,N24663);
and and14705(N24661,N24664,N24665);
and and14713(N24676,N24678,N24679);
and and14714(N24677,N24680,N24681);
and and14722(N24692,N24694,N24695);
and and14723(N24693,N24696,N24697);
and and14731(N24708,N24710,N24711);
and and14732(N24709,N24712,N24713);
and and14740(N24724,N24726,N24727);
and and14741(N24725,N24728,N24729);
and and14749(N24740,N24742,N24743);
and and14750(N24741,N24744,N24745);
and and14758(N24756,N24758,N24759);
and and14759(N24757,N24760,N24761);
and and14767(N24772,N24774,N24775);
and and14768(N24773,N24776,N24777);
and and14776(N24788,N24790,N24791);
and and14777(N24789,N24792,N24793);
and and14785(N24804,N24806,N24807);
and and14786(N24805,N24808,N24809);
and and14794(N24820,N24822,N24823);
and and14795(N24821,N24824,N24825);
and and14803(N24836,N24838,N24839);
and and14804(N24837,N24840,N24841);
and and14812(N24852,N24854,N24855);
and and14813(N24853,N24856,N24857);
and and14821(N24868,N24870,N24871);
and and14822(N24869,N24872,N24873);
and and14830(N24883,N24885,N24886);
and and14831(N24884,N24887,N24888);
and and14839(N24898,N24900,N24901);
and and14840(N24899,N24902,N24903);
and and14848(N24913,N24915,N24916);
and and14849(N24914,N24917,N24918);
and and14857(N24928,N24930,N24931);
and and14858(N24929,N24932,N24933);
and and14866(N24943,N24945,N24946);
and and14867(N24944,N24947,N24948);
and and14875(N24958,N24960,N24961);
and and14876(N24959,N24962,N24963);
and and14884(N24973,N24975,N24976);
and and14885(N24974,N24977,N24978);
and and14893(N24988,N24990,N24991);
and and14894(N24989,N24992,N24993);
and and14902(N25003,N25005,N25006);
and and14903(N25004,N25007,N25008);
and and14911(N25018,N25020,N25021);
and and14912(N25019,N25022,N25023);
and and14920(N25033,N25035,N25036);
and and14921(N25034,N25037,N25038);
and and14929(N25048,N25050,N25051);
and and14930(N25049,N25052,N25053);
and and14938(N25063,N25065,N25066);
and and14939(N25064,N25067,N25068);
and and14947(N25078,N25080,N25081);
and and14948(N25079,N25082,N25083);
and and14956(N25093,N25095,N25096);
and and14957(N25094,N25097,N25098);
and and14965(N25108,N25110,N25111);
and and14966(N25109,N25112,N25113);
and and14974(N25123,N25125,N25126);
and and14975(N25124,N25127,N25128);
and and14983(N25138,N25140,N25141);
and and14984(N25139,N25142,N25143);
and and14992(N25153,N25155,N25156);
and and14993(N25154,N25157,N25158);
and and15001(N25168,N25170,N25171);
and and15002(N25169,N25172,N25173);
and and15010(N25183,N25185,N25186);
and and15011(N25184,N25187,N25188);
and and15019(N25198,N25200,N25201);
and and15020(N25199,N25202,N25203);
and and15028(N25213,N25215,N25216);
and and15029(N25214,N25217,N25218);
and and15037(N25228,N25230,N25231);
and and15038(N25229,N25232,N25233);
and and15046(N25243,N25245,N25246);
and and15047(N25244,N25247,N25248);
and and15055(N25258,N25260,N25261);
and and15056(N25259,N25262,N25263);
and and15064(N25272,N25274,N25275);
and and15065(N25273,N25276,N25277);
and and15073(N25286,N25288,N25289);
and and15074(N25287,N25290,N25291);
and and15082(N25300,N25302,N25303);
and and15083(N25301,N25304,N25305);
and and15091(N25314,N25316,N25317);
and and15092(N25315,N25318,N25319);
and and15100(N25328,N25330,N25331);
and and15101(N25329,N25332,N25333);
and and15109(N25342,N25344,N25345);
and and15110(N25343,N25346,N25347);
and and15118(N25356,N25358,N25359);
and and15119(N25357,N25360,N25361);
and and15127(N25370,N25372,N25373);
and and15128(N25371,N25374,N25375);
and and15136(N25384,N25386,N25387);
and and15137(N25385,N25388,N25389);
and and15145(N25398,N25400,N25401);
and and15146(N25399,N25402,N25403);
and and15154(N25412,N25414,N25415);
and and15155(N25413,N25416,N25417);
and and15163(N25426,N25428,N25429);
and and15164(N25427,N25430,N25431);
and and15172(N25440,N25442,N25443);
and and15173(N25441,N25444,N25445);
and and15181(N25454,N25456,N25457);
and and15182(N25455,N25458,N25459);
and and15190(N25468,N25470,N25471);
and and15191(N25469,N25472,N25473);
and and15199(N25482,N25484,N25485);
and and15200(N25483,N25486,N25487);
and and15208(N25496,N25498,N25499);
and and15209(N25497,N25500,N25501);
and and15217(N25510,N25512,N25513);
and and15218(N25511,N25514,N25515);
and and15226(N25524,N25526,N25527);
and and15227(N25525,N25528,N25529);
and and15235(N25538,N25540,N25541);
and and15236(N25539,N25542,N25543);
and and15244(N25552,N25554,N25555);
and and15245(N25553,N25556,N25557);
and and15253(N25566,N25568,N25569);
and and15254(N25567,N25570,N25571);
and and15262(N25580,N25582,N25583);
and and15263(N25581,N25584,N25585);
and and15271(N25594,N25596,N25597);
and and15272(N25595,N25598,N25599);
and and15280(N25608,N25610,N25611);
and and15281(N25609,N25612,N25613);
and and15289(N25622,N25624,N25625);
and and15290(N25623,N25626,N25627);
and and15298(N25636,N25638,N25639);
and and15299(N25637,N25640,N25641);
and and15307(N25650,N25652,N25653);
and and15308(N25651,N25654,N25655);
and and15316(N25664,N25666,N25667);
and and15317(N25665,N25668,N25669);
and and15325(N25678,N25680,N25681);
and and15326(N25679,N25682,N25683);
and and15334(N25692,N25694,N25695);
and and15335(N25693,N25696,N25697);
and and15343(N25706,N25708,N25709);
and and15344(N25707,N25710,N25711);
and and15352(N25720,N25722,N25723);
and and15353(N25721,N25724,N25725);
and and15361(N25734,N25736,N25737);
and and15362(N25735,N25738,N25739);
and and15370(N25748,N25750,N25751);
and and15371(N25749,N25752,N25753);
and and15379(N25762,N25764,N25765);
and and15380(N25763,N25766,N25767);
and and15388(N25776,N25778,N25779);
and and15389(N25777,N25780,N25781);
and and15397(N25790,N25792,N25793);
and and15398(N25791,N25794,N25795);
and and15406(N25804,N25806,N25807);
and and15407(N25805,N25808,N25809);
and and15415(N25818,N25820,N25821);
and and15416(N25819,N25822,N25823);
and and15424(N25832,N25834,N25835);
and and15425(N25833,N25836,N25837);
and and15433(N25846,N25848,N25849);
and and15434(N25847,N25850,N25851);
and and15442(N25860,N25862,N25863);
and and15443(N25861,N25864,N25865);
and and15451(N25874,N25876,N25877);
and and15452(N25875,N25878,N25879);
and and15460(N25888,N25890,N25891);
and and15461(N25889,N25892,N25893);
and and15469(N25902,N25904,N25905);
and and15470(N25903,N25906,N25907);
and and15478(N25916,N25918,N25919);
and and15479(N25917,N25920,N25921);
and and15487(N25930,N25932,N25933);
and and15488(N25931,N25934,N25935);
and and15496(N25944,N25946,N25947);
and and15497(N25945,N25948,N25949);
and and15505(N25958,N25960,N25961);
and and15506(N25959,N25962,N25963);
and and15514(N25972,N25974,N25975);
and and15515(N25973,N25976,N25977);
and and15523(N25986,N25988,N25989);
and and15524(N25987,N25990,N25991);
and and15532(N26000,N26002,N26003);
and and15533(N26001,N26004,N26005);
and and15541(N26014,N26016,N26017);
and and15542(N26015,N26018,N26019);
and and15550(N26028,N26030,N26031);
and and15551(N26029,N26032,N26033);
and and15559(N26042,N26044,N26045);
and and15560(N26043,N26046,N26047);
and and15568(N26056,N26058,N26059);
and and15569(N26057,N26060,N26061);
and and15577(N26070,N26072,N26073);
and and15578(N26071,N26074,N26075);
and and15586(N26084,N26086,N26087);
and and15587(N26085,N26088,N26089);
and and15595(N26098,N26100,N26101);
and and15596(N26099,N26102,N26103);
and and15604(N26112,N26114,N26115);
and and15605(N26113,N26116,N26117);
and and15613(N26126,N26128,N26129);
and and15614(N26127,N26130,N26131);
and and15622(N26140,N26142,N26143);
and and15623(N26141,N26144,N26145);
and and15631(N26153,N26155,N26156);
and and15632(N26154,N26157,N26158);
and and15640(N26166,N26168,N26169);
and and15641(N26167,N26170,N26171);
and and15649(N26179,N26181,N26182);
and and15650(N26180,N26183,N26184);
and and15658(N26192,N26194,N26195);
and and15659(N26193,N26196,N26197);
and and15667(N26205,N26207,N26208);
and and15668(N26206,N26209,N26210);
and and15676(N26218,N26220,N26221);
and and15677(N26219,N26222,N26223);
and and15685(N26231,N26233,N26234);
and and15686(N26232,N26235,N26236);
and and15694(N26244,N26246,N26247);
and and15695(N26245,N26248,N26249);
and and15703(N26257,N26259,N26260);
and and15704(N26258,N26261,N26262);
and and15712(N26270,N26272,N26273);
and and15713(N26271,N26274,N26275);
and and15721(N26283,N26285,N26286);
and and15722(N26284,N26287,N26288);
and and15730(N26296,N26298,N26299);
and and15731(N26297,N26300,N26301);
and and15739(N26309,N26311,N26312);
and and15740(N26310,N26313,N26314);
and and15748(N26322,N26324,N26325);
and and15749(N26323,N26326,N26327);
and and15757(N26335,N26337,N26338);
and and15758(N26336,N26339,N26340);
and and15766(N26348,N26350,N26351);
and and15767(N26349,N26352,N26353);
and and15775(N26361,N26363,N26364);
and and15776(N26362,N26365,N26366);
and and15784(N26374,N26376,N26377);
and and15785(N26375,N26378,N26379);
and and15793(N26387,N26389,N26390);
and and15794(N26388,N26391,N26392);
and and15802(N26400,N26402,N26403);
and and15803(N26401,N26404,N26405);
and and15811(N26413,N26415,N26416);
and and15812(N26414,N26417,N26418);
and and15820(N26426,N26428,N26429);
and and15821(N26427,N26430,N26431);
and and15829(N26439,N26441,N26442);
and and15830(N26440,N26443,N26444);
and and15838(N26452,N26454,N26455);
and and15839(N26453,N26456,N26457);
and and15847(N26465,N26467,N26468);
and and15848(N26466,N26469,N26470);
and and15856(N26478,N26480,N26481);
and and15857(N26479,N26482,N26483);
and and15865(N26491,N26493,N26494);
and and15866(N26492,N26495,N26496);
and and15874(N26504,N26506,N26507);
and and15875(N26505,N26508,N26509);
and and15883(N26516,N26518,N26519);
and and15884(N26517,N26520,N26521);
and and15892(N26528,N26530,N26531);
and and15893(N26529,N26532,N26533);
and and15901(N26540,N26542,N26543);
and and15902(N26541,N26544,N26545);
and and15910(N26552,N26554,N26555);
and and15911(N26553,N26556,N26557);
and and15919(N26564,N26566,N26567);
and and15920(N26565,N26568,N26569);
and and15928(N26576,N26578,N26579);
and and15929(N26577,N26580,N26581);
and and15937(N26588,N26590,N26591);
and and15938(N26589,N26592,N26593);
and and15946(N26600,N26602,N26603);
and and15947(N26601,N26604,N26605);
and and15955(N26612,N26614,N26615);
and and15956(N26613,N26616,N26617);
and and15964(N26624,N26626,N26627);
and and15965(N26625,N26628,N26629);
and and15973(N26636,N26638,N26639);
and and15974(N26637,N26640,N26641);
and and15982(N26648,N26650,N26651);
and and15983(N26649,N26652,N26653);
and and15991(N26660,N26662,N26663);
and and15992(N26661,N26664,N26665);
and and16000(N26672,N26674,N26675);
and and16001(N26673,N26676,N26677);
and and16009(N26684,N26686,N26687);
and and16010(N26685,N26688,N26689);
and and16018(N26696,N26698,N26699);
and and16019(N26697,N26700,N26701);
and and16027(N26708,N26710,N26711);
and and16028(N26709,N26712,N26713);
and and16036(N26720,N26722,N26723);
and and16037(N26721,N26724,N26725);
and and16045(N26732,N26734,N26735);
and and16046(N26733,N26736,N26737);
and and16054(N26744,N26746,N26747);
and and16055(N26745,N26748,N26749);
and and16063(N26756,N26758,N26759);
and and16064(N26757,N26760,N26761);
and and16072(N26768,N26770,N26771);
and and16073(N26769,N26772,N26773);
and and16081(N26780,N26782,N26783);
and and16082(N26781,N26784,N26785);
and and16090(N26792,N26794,N26795);
and and16091(N26793,N26796,N26797);
and and16099(N26804,N26806,N26807);
and and16100(N26805,N26808,N26809);
and and16108(N26816,N26818,N26819);
and and16109(N26817,N26820,N26821);
and and16117(N26828,N26830,N26831);
and and16118(N26829,N26832,N26833);
and and16126(N26840,N26842,N26843);
and and16127(N26841,N26844,N26845);
and and16135(N26852,N26854,N26855);
and and16136(N26853,N26856,N26857);
and and16144(N26864,N26866,N26867);
and and16145(N26865,N26868,N26869);
and and16153(N26876,N26878,N26879);
and and16154(N26877,N26880,N26881);
and and16162(N26888,N26890,N26891);
and and16163(N26889,N26892,N26893);
and and16171(N26900,N26902,N26903);
and and16172(N26901,N26904,N26905);
and and16180(N26912,N26914,N26915);
and and16181(N26913,N26916,N26917);
and and16189(N26924,N26926,N26927);
and and16190(N26925,N26928,N26929);
and and16198(N26936,N26938,N26939);
and and16199(N26937,N26940,N26941);
and and16207(N26948,N26950,N26951);
and and16208(N26949,N26952,N26953);
and and16216(N26960,N26962,N26963);
and and16217(N26961,N26964,N26965);
and and16225(N26972,N26974,N26975);
and and16226(N26973,N26976,N26977);
and and16234(N26983,N26985,N26986);
and and16235(N26984,N26987,N26988);
and and16243(N26994,N26996,N26997);
and and16244(N26995,N26998,N26999);
and and16252(N27005,N27007,N27008);
and and16253(N27006,N27009,N27010);
and and16261(N27016,N27018,N27019);
and and16262(N27017,N27020,N27021);
and and16270(N27027,N27029,N27030);
and and16271(N27028,N27031,N27032);
and and16279(N27038,N27040,N27041);
and and16280(N27039,N27042,N27043);
and and16288(N27049,N27051,N27052);
and and16289(N27050,N27053,N27054);
and and16297(N27060,N27062,N27063);
and and16298(N27061,N27064,N27065);
and and16306(N27071,N27073,N27074);
and and16307(N27072,N27075,N27076);
and and16315(N27082,N27084,N27085);
and and16316(N27083,N27086,N27087);
and and16324(N27093,N27095,N27096);
and and16325(N27094,N27097,N27098);
and and16333(N27104,N27106,N27107);
and and16334(N27105,N27108,N27109);
and and16342(N27115,N27117,N27118);
and and16343(N27116,N27119,N27120);
and and16351(N27126,N27128,N27129);
and and16352(N27127,N27130,N27131);
and and16360(N27137,N27139,N27140);
and and16361(N27138,N27141,N27142);
and and16369(N27148,N27150,N27151);
and and16370(N27149,N27152,N27153);
and and16378(N27158,N27160,N27161);
and and16379(N27159,N27162,N27163);
and and16387(N27168,N27170,N27171);
and and16388(N27169,N27172,N27173);
and and16396(N27178,N27180,N27181);
and and16397(N27179,N27182,N27183);
and and16405(N27188,N27190,N27191);
and and16406(N27189,N27192,N27193);
and and16414(N27198,N27200,N27201);
and and16415(N27199,N27202,N27203);
and and16422(N27214,N27216,N27217);
and and16423(N27215,N27218,N27219);
and and16430(N27230,N27232,N27233);
and and16431(N27231,N27234,N27235);
and and16438(N27246,N27248,N27249);
and and16439(N27247,N27250,N27251);
and and16446(N27261,N27263,N27264);
and and16447(N27262,N27265,N27266);
and and16454(N27276,N27278,N27279);
and and16455(N27277,N27280,N27281);
and and16462(N27291,N27293,N27294);
and and16463(N27292,N27295,N27296);
and and16470(N27306,N27308,N27309);
and and16471(N27307,N27310,N27311);
and and16478(N27321,N27323,N27324);
and and16479(N27322,N27325,N27326);
and and16486(N27336,N27338,N27339);
and and16487(N27337,N27340,N27341);
and and16494(N27351,N27353,N27354);
and and16495(N27352,N27355,N27356);
and and16502(N27366,N27368,N27369);
and and16503(N27367,N27370,N27371);
and and16510(N27381,N27383,N27384);
and and16511(N27382,N27385,N27386);
and and16518(N27396,N27398,N27399);
and and16519(N27397,N27400,N27401);
and and16526(N27411,N27413,N27414);
and and16527(N27412,N27415,N27416);
and and16534(N27425,N27427,N27428);
and and16535(N27426,N27429,N27430);
and and16542(N27439,N27441,N27442);
and and16543(N27440,N27443,N27444);
and and16550(N27453,N27455,N27456);
and and16551(N27454,N27457,N27458);
and and16558(N27467,N27469,N27470);
and and16559(N27468,N27471,N27472);
and and16566(N27481,N27483,N27484);
and and16567(N27482,N27485,N27486);
and and16574(N27495,N27497,N27498);
and and16575(N27496,N27499,N27500);
and and16582(N27509,N27511,N27512);
and and16583(N27510,N27513,N27514);
and and16590(N27523,N27525,N27526);
and and16591(N27524,N27527,N27528);
and and16598(N27537,N27539,N27540);
and and16599(N27538,N27541,N27542);
and and16606(N27551,N27553,N27554);
and and16607(N27552,N27555,N27556);
and and16614(N27565,N27567,N27568);
and and16615(N27566,N27569,N27570);
and and16622(N27579,N27581,N27582);
and and16623(N27580,N27583,N27584);
and and16630(N27593,N27595,N27596);
and and16631(N27594,N27597,N27598);
and and16638(N27607,N27609,N27610);
and and16639(N27608,N27611,N27612);
and and16646(N27621,N27623,N27624);
and and16647(N27622,N27625,N27626);
and and16654(N27635,N27637,N27638);
and and16655(N27636,N27639,N27640);
and and16662(N27649,N27651,N27652);
and and16663(N27650,N27653,N27654);
and and16670(N27663,N27665,N27666);
and and16671(N27664,N27667,N27668);
and and16678(N27677,N27679,N27680);
and and16679(N27678,N27681,N27682);
and and16686(N27691,N27693,N27694);
and and16687(N27692,N27695,N27696);
and and16694(N27705,N27707,N27708);
and and16695(N27706,N27709,N27710);
and and16702(N27719,N27721,N27722);
and and16703(N27720,N27723,N27724);
and and16710(N27733,N27735,N27736);
and and16711(N27734,N27737,N27738);
and and16718(N27747,N27749,N27750);
and and16719(N27748,N27751,N27752);
and and16726(N27760,N27762,N27763);
and and16727(N27761,N27764,N27765);
and and16734(N27773,N27775,N27776);
and and16735(N27774,N27777,N27778);
and and16742(N27786,N27788,N27789);
and and16743(N27787,N27790,N27791);
and and16750(N27799,N27801,N27802);
and and16751(N27800,N27803,N27804);
and and16758(N27812,N27814,N27815);
and and16759(N27813,N27816,N27817);
and and16766(N27825,N27827,N27828);
and and16767(N27826,N27829,N27830);
and and16774(N27838,N27840,N27841);
and and16775(N27839,N27842,N27843);
and and16782(N27851,N27853,N27854);
and and16783(N27852,N27855,N27856);
and and16790(N27864,N27866,N27867);
and and16791(N27865,N27868,N27869);
and and16798(N27877,N27879,N27880);
and and16799(N27878,N27881,N27882);
and and16806(N27890,N27892,N27893);
and and16807(N27891,N27894,N27895);
and and16814(N27903,N27905,N27906);
and and16815(N27904,N27907,N27908);
and and16822(N27916,N27918,N27919);
and and16823(N27917,N27920,N27921);
and and16830(N27929,N27931,N27932);
and and16831(N27930,N27933,N27934);
and and16838(N27942,N27944,N27945);
and and16839(N27943,N27946,N27947);
and and16846(N27955,N27957,N27958);
and and16847(N27956,N27959,N27960);
and and16854(N27968,N27970,N27971);
and and16855(N27969,N27972,N27973);
and and16862(N27981,N27983,N27984);
and and16863(N27982,N27985,N27986);
and and16870(N27994,N27996,N27997);
and and16871(N27995,N27998,N27999);
and and16878(N28007,N28009,N28010);
and and16879(N28008,N28011,N28012);
and and16886(N28020,N28022,N28023);
and and16887(N28021,N28024,N28025);
and and16894(N28033,N28035,N28036);
and and16895(N28034,N28037,N28038);
and and16902(N28046,N28048,N28049);
and and16903(N28047,N28050,N28051);
and and16910(N28059,N28061,N28062);
and and16911(N28060,N28063,N28064);
and and16918(N28072,N28074,N28075);
and and16919(N28073,N28076,N28077);
and and16926(N28085,N28087,N28088);
and and16927(N28086,N28089,N28090);
and and16934(N28098,N28100,N28101);
and and16935(N28099,N28102,N28103);
and and16942(N28111,N28113,N28114);
and and16943(N28112,N28115,N28116);
and and16950(N28124,N28126,N28127);
and and16951(N28125,N28128,N28129);
and and16958(N28137,N28139,N28140);
and and16959(N28138,N28141,N28142);
and and16966(N28150,N28152,N28153);
and and16967(N28151,N28154,N28155);
and and16974(N28163,N28165,N28166);
and and16975(N28164,N28167,N28168);
and and16982(N28175,N28177,N28178);
and and16983(N28176,N28179,N28180);
and and16990(N28187,N28189,N28190);
and and16991(N28188,N28191,N28192);
and and16998(N28199,N28201,N28202);
and and16999(N28200,N28203,N28204);
and and17006(N28211,N28213,N28214);
and and17007(N28212,N28215,N28216);
and and17014(N28223,N28225,N28226);
and and17015(N28224,N28227,N28228);
and and17022(N28235,N28237,N28238);
and and17023(N28236,N28239,N28240);
and and17030(N28247,N28249,N28250);
and and17031(N28248,N28251,N28252);
and and17038(N28259,N28261,N28262);
and and17039(N28260,N28263,N28264);
and and17046(N28271,N28273,N28274);
and and17047(N28272,N28275,N28276);
and and17054(N28283,N28285,N28286);
and and17055(N28284,N28287,N28288);
and and17062(N28295,N28297,N28298);
and and17063(N28296,N28299,N28300);
and and17070(N28307,N28309,N28310);
and and17071(N28308,N28311,N28312);
and and17078(N28319,N28321,N28322);
and and17079(N28320,N28323,N28324);
and and17086(N28331,N28333,N28334);
and and17087(N28332,N28335,N28336);
and and17094(N28343,N28345,N28346);
and and17095(N28344,N28347,N28348);
and and17102(N28355,N28357,N28358);
and and17103(N28356,N28359,N28360);
and and17110(N28367,N28369,N28370);
and and17111(N28368,N28371,N28372);
and and17118(N28379,N28381,N28382);
and and17119(N28380,N28383,N28384);
and and17126(N28391,N28393,N28394);
and and17127(N28392,N28395,N28396);
and and17134(N28403,N28405,N28406);
and and17135(N28404,N28407,N28408);
and and17142(N28415,N28417,N28418);
and and17143(N28416,N28419,N28420);
and and17150(N28427,N28429,N28430);
and and17151(N28428,N28431,N28432);
and and17158(N28439,N28441,N28442);
and and17159(N28440,N28443,N28444);
and and17166(N28451,N28453,N28454);
and and17167(N28452,N28455,N28456);
and and17174(N28463,N28465,N28466);
and and17175(N28464,N28467,N28468);
and and17182(N28475,N28477,N28478);
and and17183(N28476,N28479,N28480);
and and17190(N28487,N28489,N28490);
and and17191(N28488,N28491,N28492);
and and17198(N28499,N28501,N28502);
and and17199(N28500,N28503,N28504);
and and17206(N28511,N28513,N28514);
and and17207(N28512,N28515,N28516);
and and17214(N28523,N28525,N28526);
and and17215(N28524,N28527,N28528);
and and17222(N28535,N28537,N28538);
and and17223(N28536,N28539,N28540);
and and17230(N28547,N28549,N28550);
and and17231(N28548,N28551,N28552);
and and17238(N28559,N28561,N28562);
and and17239(N28560,N28563,N28564);
and and17246(N28571,N28573,N28574);
and and17247(N28572,N28575,N28576);
and and17254(N28583,N28585,N28586);
and and17255(N28584,N28587,N28588);
and and17262(N28595,N28597,N28598);
and and17263(N28596,N28599,N28600);
and and17270(N28607,N28609,N28610);
and and17271(N28608,N28611,N28612);
and and17278(N28619,N28621,N28622);
and and17279(N28620,N28623,N28624);
and and17286(N28631,N28633,N28634);
and and17287(N28632,N28635,N28636);
and and17294(N28643,N28645,N28646);
and and17295(N28644,N28647,N28648);
and and17302(N28655,N28657,N28658);
and and17303(N28656,N28659,N28660);
and and17310(N28666,N28668,N28669);
and and17311(N28667,N28670,N28671);
and and17318(N28677,N28679,N28680);
and and17319(N28678,N28681,N28682);
and and17326(N28688,N28690,N28691);
and and17327(N28689,N28692,N28693);
and and17334(N28699,N28701,N28702);
and and17335(N28700,N28703,N28704);
and and17342(N28710,N28712,N28713);
and and17343(N28711,N28714,N28715);
and and17350(N28721,N28723,N28724);
and and17351(N28722,N28725,N28726);
and and17358(N28732,N28734,N28735);
and and17359(N28733,N28736,N28737);
and and17366(N28743,N28745,N28746);
and and17367(N28744,N28747,N28748);
and and17374(N28754,N28756,N28757);
and and17375(N28755,N28758,N28759);
and and17382(N28765,N28767,N28768);
and and17383(N28766,N28769,N28770);
and and17390(N28776,N28778,N28779);
and and17391(N28777,N28780,N28781);
and and17398(N28787,N28789,N28790);
and and17399(N28788,N28791,N28792);
and and17406(N28798,N28800,N28801);
and and17407(N28799,N28802,N28803);
and and17414(N28809,N28811,N28812);
and and17415(N28810,N28813,N28814);
and and17422(N28820,N28822,N28823);
and and17423(N28821,N28824,N28825);
and and17430(N28831,N28833,N28834);
and and17431(N28832,N28835,N28836);
and and17438(N28842,N28844,N28845);
and and17439(N28843,N28846,N28847);
and and17446(N28853,N28855,N28856);
and and17447(N28854,N28857,N28858);
and and17454(N28864,N28866,N28867);
and and17455(N28865,N28868,N28869);
and and17462(N28875,N28877,N28878);
and and17463(N28876,N28879,N28880);
and and17470(N28886,N28888,N28889);
and and17471(N28887,N28890,N28891);
and and17478(N28897,N28899,N28900);
and and17479(N28898,N28901,N28902);
and and17486(N28908,N28910,N28911);
and and17487(N28909,N28912,N28913);
and and17494(N28919,N28921,N28922);
and and17495(N28920,N28923,N28924);
and and17502(N28930,N28932,N28933);
and and17503(N28931,N28934,N28935);
and and17510(N28940,N28942,N28943);
and and17511(N28941,N28944,N28945);
and and17518(N28950,N28952,N28953);
and and17519(N28951,N28954,N28955);
and and17526(N28960,N28962,N28963);
and and17527(N28961,N28964,N28965);
and and17534(N28970,N28972,N28973);
and and17535(N28971,N28974,N28975);
and and17542(N28980,N28982,N28983);
and and17543(N28981,N28984,N28985);
and and17550(N28990,N28992,N28993);
and and17551(N28991,N28994,N28995);
and and17558(N29000,N29002,N29003);
and and17559(N29001,N29004,N29005);
and and17566(N29010,N29012,N29013);
and and17567(N29011,N29014,N29015);
and and17574(N29020,N29022,N29023);
and and17575(N29021,N29024,N29025);
and and17582(N29030,N29032,N29033);
and and17583(N29031,N29034,N29035);
and and17590(N29040,N29042,N29043);
and and17591(N29041,N29044,N29045);
and and17598(N29050,N29052,N29053);
and and17599(N29051,N29054,N29055);
and and17606(N29059,N29061,N29062);
and and17607(N29060,N29063,N29064);
and and17613(N29072,N29074,N29075);
and and17614(N29073,N29076,N29077);
and and17620(N29085,N29087,N29088);
and and17621(N29086,N29089,N29090);
and and17627(N29098,N29100,N29101);
and and17628(N29099,N29102,N29103);
and and17634(N29110,N29112,N29113);
and and17635(N29111,N29114,N29115);
and and17641(N29122,N29124,N29125);
and and17642(N29123,N29126,N29127);
and and17648(N29134,N29136,N29137);
and and17649(N29135,N29138,N29139);
and and17655(N29146,N29148,N29149);
and and17656(N29147,N29150,N29151);
and and17662(N29158,N29160,N29161);
and and17663(N29159,N29162,N29163);
and and17669(N29169,N29171,N29172);
and and17670(N29170,N29173,N29174);
and and17676(N29180,N29182,N29183);
and and17677(N29181,N29184,N29185);
and and17683(N29191,N29193,N29194);
and and17684(N29192,N29195,N29196);
and and17690(N29202,N29204,N29205);
and and17691(N29203,N29206,N29207);
and and17697(N29213,N29215,N29216);
and and17698(N29214,N29217,N29218);
and and17704(N29224,N29226,N29227);
and and17705(N29225,N29228,N29229);
and and17711(N29235,N29237,N29238);
and and17712(N29236,N29239,N29240);
and and17718(N29245,N29247,N29248);
and and17719(N29246,N29249,N29250);
and and17725(N29255,N29257,N29258);
and and17726(N29256,N29259,N29260);
and and17732(N29264,N29266,N29267);
and and17733(N29265,N29268,in0);
and and14580(N24430,N24434,N24435);
and and14581(N24431,N24436,N24437);
and and14582(N24432,N24438,N24439);
and and14583(N24433,N24440,R2);
and and14589(N24447,N24451,N24452);
and and14590(N24448,N24453,in1);
and and14591(N24449,in2,N24454);
and and14592(N24450,N24455,N24456);
and and14598(N24464,N24468,N24469);
and and14599(N24465,N24470,N24471);
and and14600(N24466,in2,N24472);
and and14601(N24467,N24473,N24474);
and and14607(N24481,N24485,N24486);
and and14608(N24482,N24487,in1);
and and14609(N24483,N24488,N24489);
and and14610(N24484,R2,N24490);
and and14616(N24498,N24502,N24503);
and and14617(N24499,N24504,N24505);
and and14618(N24500,in2,N24506);
and and14619(N24501,N24507,R2);
and and14625(N24515,N24519,N24520);
and and14626(N24516,N24521,N24522);
and and14627(N24517,N24523,R0);
and and14628(N24518,N24524,N24525);
and and14634(N24532,N24536,N24537);
and and14635(N24533,N24538,N24539);
and and14636(N24534,N24540,N24541);
and and14637(N24535,R1,N24542);
and and14643(N24549,N24553,N24554);
and and14644(N24550,N24555,N24556);
and and14645(N24551,N24557,N24558);
and and14646(N24552,R1,N24559);
and and14652(N24566,N24570,N24571);
and and14653(N24567,N24572,N24573);
and and14654(N24568,N24574,R1);
and and14655(N24569,N24575,R3);
and and14661(N24582,N24586,N24587);
and and14662(N24583,N24588,in2);
and and14663(N24584,N24589,N24590);
and and14664(N24585,N24591,R3);
and and14670(N24598,N24602,N24603);
and and14671(N24599,in0,in2);
and and14672(N24600,N24604,N24605);
and and14673(N24601,N24606,N24607);
and and14679(N24614,N24618,N24619);
and and14680(N24615,N24620,in2);
and and14681(N24616,N24621,N24622);
and and14682(N24617,N24623,R3);
and and14688(N24630,N24634,N24635);
and and14689(N24631,N24636,N24637);
and and14690(N24632,R0,N24638);
and and14691(N24633,R2,N24639);
and and14697(N24646,N24650,N24651);
and and14698(N24647,N24652,N24653);
and and14699(N24648,R0,R1);
and and14700(N24649,R2,N24654);
and and14706(N24662,N24666,N24667);
and and14707(N24663,N24668,N24669);
and and14708(N24664,R0,R1);
and and14709(N24665,N24670,N24671);
and and14715(N24678,N24682,N24683);
and and14716(N24679,N24684,N24685);
and and14717(N24680,N24686,N24687);
and and14718(N24681,N24688,R2);
and and14724(N24694,N24698,N24699);
and and14725(N24695,N24700,N24701);
and and14726(N24696,in2,N24702);
and and14727(N24697,N24703,N24704);
and and14733(N24710,N24714,N24715);
and and14734(N24711,N24716,N24717);
and and14735(N24712,N24718,R1);
and and14736(N24713,N24719,N24720);
and and14742(N24726,N24730,N24731);
and and14743(N24727,N24732,N24733);
and and14744(N24728,in2,N24734);
and and14745(N24729,R1,N24735);
and and14751(N24742,N24746,N24747);
and and14752(N24743,N24748,N24749);
and and14753(N24744,in2,R1);
and and14754(N24745,N24750,N24751);
and and14760(N24758,N24762,N24763);
and and14761(N24759,N24764,N24765);
and and14762(N24760,in2,R0);
and and14763(N24761,N24766,N24767);
and and14769(N24774,N24778,N24779);
and and14770(N24775,N24780,N24781);
and and14771(N24776,N24782,N24783);
and and14772(N24777,R1,R2);
and and14778(N24790,N24794,N24795);
and and14779(N24791,N24796,in1);
and and14780(N24792,in2,N24797);
and and14781(N24793,N24798,R3);
and and14787(N24806,N24810,N24811);
and and14788(N24807,N24812,in1);
and and14789(N24808,N24813,N24814);
and and14790(N24809,R1,N24815);
and and14796(N24822,N24826,N24827);
and and14797(N24823,N24828,N24829);
and and14798(N24824,in2,N24830);
and and14799(N24825,R1,N24831);
and and14805(N24838,N24842,N24843);
and and14806(N24839,N24844,in1);
and and14807(N24840,in2,R0);
and and14808(N24841,N24845,N24846);
and and14814(N24854,N24858,N24859);
and and14815(N24855,N24860,N24861);
and and14816(N24856,N24862,R1);
and and14817(N24857,R2,N24863);
and and14823(N24870,N24874,N24875);
and and14824(N24871,in0,N24876);
and and14825(N24872,R0,N24877);
and and14826(N24873,R2,R3);
and and14832(N24885,N24889,N24890);
and and14833(N24886,N24891,N24892);
and and14834(N24887,N24893,R1);
and and14835(N24888,N24894,R3);
and and14841(N24900,N24904,N24905);
and and14842(N24901,N24906,in1);
and and14843(N24902,in2,N24907);
and and14844(N24903,N24908,R2);
and and14850(N24915,N24919,N24920);
and and14851(N24916,N24921,N24922);
and and14852(N24917,R0,N24923);
and and14853(N24918,R2,R3);
and and14859(N24930,N24934,N24935);
and and14860(N24931,N24936,N24937);
and and14861(N24932,R0,N24938);
and and14862(N24933,N24939,R3);
and and14868(N24945,N24949,N24950);
and and14869(N24946,N24951,in1);
and and14870(N24947,N24952,N24953);
and and14871(N24948,R1,N24954);
and and14877(N24960,N24964,N24965);
and and14878(N24961,N24966,N24967);
and and14879(N24962,R0,R1);
and and14880(N24963,N24968,N24969);
and and14886(N24975,N24979,N24980);
and and14887(N24976,N24981,N24982);
and and14888(N24977,N24983,N24984);
and and14889(N24978,R1,N24985);
and and14895(N24990,N24994,N24995);
and and14896(N24991,in0,N24996);
and and14897(N24992,N24997,N24998);
and and14898(N24993,R2,N24999);
and and14904(N25005,N25009,N25010);
and and14905(N25006,in1,N25011);
and and14906(N25007,N25012,N25013);
and and14907(N25008,R2,N25014);
and and14913(N25020,N25024,N25025);
and and14914(N25021,in0,N25026);
and and14915(N25022,in2,N25027);
and and14916(N25023,N25028,R2);
and and14922(N25035,N25039,N25040);
and and14923(N25036,N25041,in2);
and and14924(N25037,N25042,N25043);
and and14925(N25038,R2,R3);
and and14931(N25050,N25054,N25055);
and and14932(N25051,N25056,N25057);
and and14933(N25052,R0,N25058);
and and14934(N25053,R2,N25059);
and and14940(N25065,N25069,N25070);
and and14941(N25066,N25071,N25072);
and and14942(N25067,N25073,R0);
and and14943(N25068,N25074,R3);
and and14949(N25080,N25084,N25085);
and and14950(N25081,in0,in2);
and and14951(N25082,N25086,N25087);
and and14952(N25083,N25088,N25089);
and and14958(N25095,N25099,N25100);
and and14959(N25096,N25101,in1);
and and14960(N25097,in2,N25102);
and and14961(N25098,N25103,N25104);
and and14967(N25110,N25114,N25115);
and and14968(N25111,N25116,in1);
and and14969(N25112,N25117,R1);
and and14970(N25113,N25118,N25119);
and and14976(N25125,N25129,N25130);
and and14977(N25126,in0,N25131);
and and14978(N25127,in2,N25132);
and and14979(N25128,N25133,N25134);
and and14985(N25140,N25144,N25145);
and and14986(N25141,N25146,in1);
and and14987(N25142,in2,N25147);
and and14988(N25143,N25148,R3);
and and14994(N25155,N25159,N25160);
and and14995(N25156,N25161,N25162);
and and14996(N25157,N25163,R1);
and and14997(N25158,N25164,R3);
and and15003(N25170,N25174,N25175);
and and15004(N25171,N25176,N25177);
and and15005(N25172,N25178,N25179);
and and15006(N25173,R2,N25180);
and and15012(N25185,N25189,N25190);
and and15013(N25186,N25191,N25192);
and and15014(N25187,N25193,N25194);
and and15015(N25188,N25195,R2);
and and15021(N25200,N25204,N25205);
and and15022(N25201,N25206,in1);
and and15023(N25202,N25207,N25208);
and and15024(N25203,N25209,R2);
and and15030(N25215,N25219,N25220);
and and15031(N25216,N25221,in2);
and and15032(N25217,R0,N25222);
and and15033(N25218,R2,N25223);
and and15039(N25230,N25234,N25235);
and and15040(N25231,N25236,in1);
and and15041(N25232,N25237,R0);
and and15042(N25233,N25238,R2);
and and15048(N25245,N25249,N25250);
and and15049(N25246,N25251,N25252);
and and15050(N25247,N25253,R0);
and and15051(N25248,N25254,R3);
and and15057(N25260,N25264,N25265);
and and15058(N25261,N25266,N25267);
and and15059(N25262,R0,R1);
and and15060(N25263,N25268,R3);
and and15066(N25274,N25278,N25279);
and and15067(N25275,in0,in1);
and and15068(N25276,in2,N25280);
and and15069(N25277,N25281,R3);
and and15075(N25288,N25292,N25293);
and and15076(N25289,N25294,in1);
and and15077(N25290,N25295,R0);
and and15078(N25291,N25296,R2);
and and15084(N25302,N25306,N25307);
and and15085(N25303,N25308,in2);
and and15086(N25304,N25309,R1);
and and15087(N25305,N25310,R3);
and and15093(N25316,N25320,N25321);
and and15094(N25317,N25322,in2);
and and15095(N25318,N25323,R1);
and and15096(N25319,R2,N25324);
and and15102(N25330,N25334,N25335);
and and15103(N25331,N25336,N25337);
and and15104(N25332,N25338,R1);
and and15105(N25333,R2,R3);
and and15111(N25344,N25348,N25349);
and and15112(N25345,N25350,N25351);
and and15113(N25346,R0,R1);
and and15114(N25347,R2,N25352);
and and15120(N25358,N25362,N25363);
and and15121(N25359,N25364,in2);
and and15122(N25360,N25365,R1);
and and15123(N25361,R2,N25366);
and and15129(N25372,N25376,N25377);
and and15130(N25373,N25378,in1);
and and15131(N25374,in2,R0);
and and15132(N25375,N25379,R2);
and and15138(N25386,N25390,N25391);
and and15139(N25387,in0,N25392);
and and15140(N25388,R0,R1);
and and15141(N25389,N25393,R3);
and and15147(N25400,N25404,N25405);
and and15148(N25401,N25406,in2);
and and15149(N25402,R0,R1);
and and15150(N25403,N25407,R3);
and and15156(N25414,N25418,N25419);
and and15157(N25415,in0,in1);
and and15158(N25416,N25420,N25421);
and and15159(N25417,R1,N25422);
and and15165(N25428,N25432,N25433);
and and15166(N25429,N25434,in1);
and and15167(N25430,in2,N25435);
and and15168(N25431,R1,N25436);
and and15174(N25442,N25446,N25447);
and and15175(N25443,N25448,in2);
and and15176(N25444,N25449,R1);
and and15177(N25445,N25450,N25451);
and and15183(N25456,N25460,N25461);
and and15184(N25457,in0,in2);
and and15185(N25458,N25462,N25463);
and and15186(N25459,R2,N25464);
and and15192(N25470,N25474,N25475);
and and15193(N25471,N25476,N25477);
and and15194(N25472,N25478,R0);
and and15195(N25473,N25479,R2);
and and15201(N25484,N25488,N25489);
and and15202(N25485,N25490,N25491);
and and15203(N25486,N25492,N25493);
and and15204(N25487,R2,R3);
and and15210(N25498,N25502,N25503);
and and15211(N25499,N25504,N25505);
and and15212(N25500,R0,N25506);
and and15213(N25501,N25507,R3);
and and15219(N25512,N25516,N25517);
and and15220(N25513,N25518,in1);
and and15221(N25514,N25519,R1);
and and15222(N25515,R2,R3);
and and15228(N25526,N25530,N25531);
and and15229(N25527,N25532,N25533);
and and15230(N25528,in2,R1);
and and15231(N25529,R2,N25534);
and and15237(N25540,N25544,N25545);
and and15238(N25541,N25546,in1);
and and15239(N25542,N25547,R1);
and and15240(N25543,R2,N25548);
and and15246(N25554,N25558,N25559);
and and15247(N25555,in1,in2);
and and15248(N25556,R0,R1);
and and15249(N25557,N25560,N25561);
and and15255(N25568,N25572,N25573);
and and15256(N25569,N25574,N25575);
and and15257(N25570,R0,N25576);
and and15258(N25571,N25577,R3);
and and15264(N25582,N25586,N25587);
and and15265(N25583,in0,in2);
and and15266(N25584,R0,N25588);
and and15267(N25585,N25589,R3);
and and15273(N25596,N25600,N25601);
and and15274(N25597,in0,in2);
and and15275(N25598,N25602,N25603);
and and15276(N25599,R2,R3);
and and15282(N25610,N25614,N25615);
and and15283(N25611,in0,in1);
and and15284(N25612,N25616,N25617);
and and15285(N25613,N25618,R2);
and and15291(N25624,N25628,N25629);
and and15292(N25625,N25630,N25631);
and and15293(N25626,N25632,R0);
and and15294(N25627,N25633,R3);
and and15300(N25638,N25642,N25643);
and and15301(N25639,N25644,in1);
and and15302(N25640,N25645,R1);
and and15303(N25641,R2,R3);
and and15309(N25652,N25656,N25657);
and and15310(N25653,in1,N25658);
and and15311(N25654,R0,R1);
and and15312(N25655,N25659,N25660);
and and15318(N25666,N25670,N25671);
and and15319(N25667,N25672,N25673);
and and15320(N25668,in2,R0);
and and15321(N25669,R1,R2);
and and15327(N25680,N25684,N25685);
and and15328(N25681,in0,in1);
and and15329(N25682,N25686,N25687);
and and15330(N25683,N25688,R3);
and and15336(N25694,N25698,N25699);
and and15337(N25695,in0,in1);
and and15338(N25696,N25700,N25701);
and and15339(N25697,N25702,R3);
and and15345(N25708,N25712,N25713);
and and15346(N25709,N25714,N25715);
and and15347(N25710,in2,N25716);
and and15348(N25711,R1,R3);
and and15354(N25722,N25726,N25727);
and and15355(N25723,in1,N25728);
and and15356(N25724,N25729,R1);
and and15357(N25725,N25730,R3);
and and15363(N25736,N25740,N25741);
and and15364(N25737,N25742,in1);
and and15365(N25738,N25743,N25744);
and and15366(N25739,N25745,R2);
and and15372(N25750,N25754,N25755);
and and15373(N25751,N25756,N25757);
and and15374(N25752,in2,N25758);
and and15375(N25753,N25759,R2);
and and15381(N25764,N25768,N25769);
and and15382(N25765,in1,in2);
and and15383(N25766,N25770,N25771);
and and15384(N25767,R2,N25772);
and and15390(N25778,N25782,N25783);
and and15391(N25779,N25784,in1);
and and15392(N25780,in2,N25785);
and and15393(N25781,R1,N25786);
and and15399(N25792,N25796,N25797);
and and15400(N25793,in0,in1);
and and15401(N25794,in2,N25798);
and and15402(N25795,R1,N25799);
and and15408(N25806,N25810,N25811);
and and15409(N25807,N25812,in1);
and and15410(N25808,N25813,N25814);
and and15411(N25809,N25815,R3);
and and15417(N25820,N25824,N25825);
and and15418(N25821,in0,N25826);
and and15419(N25822,N25827,R0);
and and15420(N25823,N25828,R2);
and and15426(N25834,N25838,N25839);
and and15427(N25835,in1,N25840);
and and15428(N25836,N25841,R1);
and and15429(N25837,R2,R3);
and and15435(N25848,N25852,N25853);
and and15436(N25849,N25854,in1);
and and15437(N25850,in2,R0);
and and15438(N25851,N25855,R3);
and and15444(N25862,N25866,N25867);
and and15445(N25863,N25868,N25869);
and and15446(N25864,N25870,R0);
and and15447(N25865,R1,N25871);
and and15453(N25876,N25880,N25881);
and and15454(N25877,in0,in2);
and and15455(N25878,N25882,R1);
and and15456(N25879,N25883,N25884);
and and15462(N25890,N25894,N25895);
and and15463(N25891,N25896,in2);
and and15464(N25892,N25897,R1);
and and15465(N25893,N25898,N25899);
and and15471(N25904,N25908,N25909);
and and15472(N25905,N25910,N25911);
and and15473(N25906,in2,N25912);
and and15474(N25907,N25913,R2);
and and15480(N25918,N25922,N25923);
and and15481(N25919,N25924,in1);
and and15482(N25920,N25925,N25926);
and and15483(N25921,R2,N25927);
and and15489(N25932,N25936,N25937);
and and15490(N25933,N25938,N25939);
and and15491(N25934,in2,N25940);
and and15492(N25935,R2,R3);
and and15498(N25946,N25950,N25951);
and and15499(N25947,N25952,N25953);
and and15500(N25948,in2,R0);
and and15501(N25949,N25954,R2);
and and15507(N25960,N25964,N25965);
and and15508(N25961,N25966,in1);
and and15509(N25962,in2,N25967);
and and15510(N25963,R2,R3);
and and15516(N25974,N25978,N25979);
and and15517(N25975,N25980,in1);
and and15518(N25976,R0,R1);
and and15519(N25977,N25981,R3);
and and15525(N25988,N25992,N25993);
and and15526(N25989,N25994,in1);
and and15527(N25990,in2,R0);
and and15528(N25991,R1,N25995);
and and15534(N26002,N26006,N26007);
and and15535(N26003,N26008,in1);
and and15536(N26004,N26009,R0);
and and15537(N26005,R1,R2);
and and15543(N26016,N26020,N26021);
and and15544(N26017,N26022,in1);
and and15545(N26018,R0,N26023);
and and15546(N26019,N26024,R3);
and and15552(N26030,N26034,N26035);
and and15553(N26031,N26036,N26037);
and and15554(N26032,in2,R0);
and and15555(N26033,N26038,N26039);
and and15561(N26044,N26048,N26049);
and and15562(N26045,N26050,N26051);
and and15563(N26046,N26052,R0);
and and15564(N26047,R1,R2);
and and15570(N26058,N26062,N26063);
and and15571(N26059,N26064,in1);
and and15572(N26060,N26065,R0);
and and15573(N26061,R1,R2);
and and15579(N26072,N26076,N26077);
and and15580(N26073,N26078,in1);
and and15581(N26074,in2,N26079);
and and15582(N26075,R1,R2);
and and15588(N26086,N26090,N26091);
and and15589(N26087,in0,in1);
and and15590(N26088,N26092,N26093);
and and15591(N26089,R1,R2);
and and15597(N26100,N26104,N26105);
and and15598(N26101,N26106,N26107);
and and15599(N26102,R0,N26108);
and and15600(N26103,R2,R3);
and and15606(N26114,N26118,N26119);
and and15607(N26115,N26120,in2);
and and15608(N26116,N26121,N26122);
and and15609(N26117,R2,R3);
and and15615(N26128,N26132,N26133);
and and15616(N26129,in1,N26134);
and and15617(N26130,N26135,N26136);
and and15618(N26131,R2,R3);
and and15624(N26142,N26146,N26147);
and and15625(N26143,N26148,in1);
and and15626(N26144,in2,R0);
and and15627(N26145,R1,R2);
and and15633(N26155,N26159,N26160);
and and15634(N26156,in0,in1);
and and15635(N26157,N26161,R0);
and and15636(N26158,R1,N26162);
and and15642(N26168,N26172,N26173);
and and15643(N26169,in1,N26174);
and and15644(N26170,R0,N26175);
and and15645(N26171,R2,R3);
and and15651(N26181,N26185,N26186);
and and15652(N26182,N26187,N26188);
and and15653(N26183,in2,N26189);
and and15654(N26184,R2,R3);
and and15660(N26194,N26198,N26199);
and and15661(N26195,in0,in1);
and and15662(N26196,in2,N26200);
and and15663(N26197,R2,N26201);
and and15669(N26207,N26211,N26212);
and and15670(N26208,in1,N26213);
and and15671(N26209,R0,N26214);
and and15672(N26210,R2,R3);
and and15678(N26220,N26224,N26225);
and and15679(N26221,N26226,N26227);
and and15680(N26222,in2,R0);
and and15681(N26223,R2,N26228);
and and15687(N26233,N26237,N26238);
and and15688(N26234,in0,in1);
and and15689(N26235,N26239,R1);
and and15690(N26236,R2,N26240);
and and15696(N26246,N26250,N26251);
and and15697(N26247,in0,N26252);
and and15698(N26248,in2,R0);
and and15699(N26249,N26253,R2);
and and15705(N26259,N26263,N26264);
and and15706(N26260,in1,in2);
and and15707(N26261,N26265,R1);
and and15708(N26262,N26266,N26267);
and and15714(N26272,N26276,N26277);
and and15715(N26273,in0,in1);
and and15716(N26274,R0,N26278);
and and15717(N26275,R2,N26279);
and and15723(N26285,N26289,N26290);
and and15724(N26286,N26291,in1);
and and15725(N26287,in2,N26292);
and and15726(N26288,N26293,R2);
and and15732(N26298,N26302,N26303);
and and15733(N26299,in0,N26304);
and and15734(N26300,in2,R0);
and and15735(N26301,R2,R3);
and and15741(N26311,N26315,N26316);
and and15742(N26312,N26317,in1);
and and15743(N26313,N26318,R0);
and and15744(N26314,R1,N26319);
and and15750(N26324,N26328,N26329);
and and15751(N26325,N26330,in2);
and and15752(N26326,R0,R1);
and and15753(N26327,N26331,N26332);
and and15759(N26337,N26341,N26342);
and and15760(N26338,N26343,N26344);
and and15761(N26339,in2,R0);
and and15762(N26340,N26345,R2);
and and15768(N26350,N26354,N26355);
and and15769(N26351,N26356,in1);
and and15770(N26352,N26357,R0);
and and15771(N26353,N26358,R2);
and and15777(N26363,N26367,N26368);
and and15778(N26364,in0,N26369);
and and15779(N26365,N26370,R0);
and and15780(N26366,R1,N26371);
and and15786(N26376,N26380,N26381);
and and15787(N26377,N26382,in2);
and and15788(N26378,R0,R1);
and and15789(N26379,N26383,R3);
and and15795(N26389,N26393,N26394);
and and15796(N26390,N26395,N26396);
and and15797(N26391,N26397,R0);
and and15798(N26392,R1,R2);
and and15804(N26402,N26406,N26407);
and and15805(N26403,in0,in1);
and and15806(N26404,N26408,N26409);
and and15807(N26405,R2,R3);
and and15813(N26415,N26419,N26420);
and and15814(N26416,in0,in1);
and and15815(N26417,in2,N26421);
and and15816(N26418,R1,N26422);
and and15822(N26428,N26432,N26433);
and and15823(N26429,in0,N26434);
and and15824(N26430,N26435,N26436);
and and15825(N26431,R1,R3);
and and15831(N26441,N26445,N26446);
and and15832(N26442,N26447,in1);
and and15833(N26443,N26448,N26449);
and and15834(N26444,R1,R3);
and and15840(N26454,N26458,N26459);
and and15841(N26455,N26460,in1);
and and15842(N26456,in2,R0);
and and15843(N26457,R1,R2);
and and15849(N26467,N26471,N26472);
and and15850(N26468,in0,N26473);
and and15851(N26469,in2,R1);
and and15852(N26470,R2,N26474);
and and15858(N26480,N26484,N26485);
and and15859(N26481,in0,in2);
and and15860(N26482,R0,R1);
and and15861(N26483,R2,N26486);
and and15867(N26493,N26497,N26498);
and and15868(N26494,N26499,in1);
and and15869(N26495,in2,N26500);
and and15870(N26496,N26501,R2);
and and15876(N26506,N26510,N26511);
and and15877(N26507,N26512,in2);
and and15878(N26508,R0,R1);
and and15879(N26509,N26513,R3);
and and15885(N26518,N26522,N26523);
and and15886(N26519,in1,in2);
and and15887(N26520,R0,R1);
and and15888(N26521,N26524,R3);
and and15894(N26530,N26534,N26535);
and and15895(N26531,in0,N26536);
and and15896(N26532,in2,R0);
and and15897(N26533,R1,N26537);
and and15903(N26542,N26546,N26547);
and and15904(N26543,N26548,in2);
and and15905(N26544,N26549,R1);
and and15906(N26545,R2,R3);
and and15912(N26554,N26558,N26559);
and and15913(N26555,N26560,in1);
and and15914(N26556,in2,R0);
and and15915(N26557,R1,R3);
and and15921(N26566,N26570,N26571);
and and15922(N26567,N26572,in1);
and and15923(N26568,in2,R1);
and and15924(N26569,R2,N26573);
and and15930(N26578,N26582,N26583);
and and15931(N26579,N26584,in1);
and and15932(N26580,in2,R0);
and and15933(N26581,R1,R2);
and and15939(N26590,N26594,N26595);
and and15940(N26591,in0,in1);
and and15941(N26592,in2,N26596);
and and15942(N26593,R1,R2);
and and15948(N26602,N26606,N26607);
and and15949(N26603,in0,in1);
and and15950(N26604,in2,R0);
and and15951(N26605,R1,N26608);
and and15957(N26614,N26618,N26619);
and and15958(N26615,in0,in1);
and and15959(N26616,N26620,N26621);
and and15960(N26617,R2,R3);
and and15966(N26626,N26630,N26631);
and and15967(N26627,N26632,in1);
and and15968(N26628,in2,R0);
and and15969(N26629,N26633,R3);
and and15975(N26638,N26642,N26643);
and and15976(N26639,in0,in2);
and and15977(N26640,R0,N26644);
and and15978(N26641,N26645,R3);
and and15984(N26650,N26654,N26655);
and and15985(N26651,in0,in1);
and and15986(N26652,N26656,R0);
and and15987(N26653,N26657,R3);
and and15993(N26662,N26666,N26667);
and and15994(N26663,in0,in1);
and and15995(N26664,in2,R1);
and and15996(N26665,R2,N26668);
and and16002(N26674,N26678,N26679);
and and16003(N26675,N26680,in2);
and and16004(N26676,R0,R1);
and and16005(N26677,R2,R3);
and and16011(N26686,N26690,N26691);
and and16012(N26687,in1,in2);
and and16013(N26688,R0,R1);
and and16014(N26689,R2,R3);
and and16020(N26698,N26702,N26703);
and and16021(N26699,in0,in1);
and and16022(N26700,in2,R0);
and and16023(N26701,R1,N26704);
and and16029(N26710,N26714,N26715);
and and16030(N26711,N26716,in1);
and and16031(N26712,in2,R1);
and and16032(N26713,R2,R3);
and and16038(N26722,N26726,N26727);
and and16039(N26723,in0,in1);
and and16040(N26724,in2,N26728);
and and16041(N26725,R2,R3);
and and16047(N26734,N26738,N26739);
and and16048(N26735,N26740,in2);
and and16049(N26736,N26741,N26742);
and and16050(N26737,R2,R3);
and and16056(N26746,N26750,N26751);
and and16057(N26747,in0,in1);
and and16058(N26748,in2,N26752);
and and16059(N26749,R1,N26753);
and and16065(N26758,N26762,N26763);
and and16066(N26759,in0,in1);
and and16067(N26760,in2,N26764);
and and16068(N26761,N26765,R2);
and and16074(N26770,N26774,N26775);
and and16075(N26771,in0,N26776);
and and16076(N26772,R0,R1);
and and16077(N26773,R2,R3);
and and16083(N26782,N26786,N26787);
and and16084(N26783,N26788,in1);
and and16085(N26784,in2,N26789);
and and16086(N26785,R1,R2);
and and16092(N26794,N26798,N26799);
and and16093(N26795,in1,in2);
and and16094(N26796,R0,R1);
and and16095(N26797,R2,R3);
and and16101(N26806,N26810,N26811);
and and16102(N26807,N26812,N26813);
and and16103(N26808,R0,R1);
and and16104(N26809,R2,R3);
and and16110(N26818,N26822,N26823);
and and16111(N26819,N26824,in1);
and and16112(N26820,in2,R0);
and and16113(N26821,R1,R3);
and and16119(N26830,N26834,N26835);
and and16120(N26831,N26836,in1);
and and16121(N26832,in2,R0);
and and16122(N26833,R2,N26837);
and and16128(N26842,N26846,N26847);
and and16129(N26843,in1,N26848);
and and16130(N26844,N26849,R1);
and and16131(N26845,R2,R3);
and and16137(N26854,N26858,N26859);
and and16138(N26855,in0,N26860);
and and16139(N26856,N26861,R1);
and and16140(N26857,R2,R3);
and and16146(N26866,N26870,N26871);
and and16147(N26867,N26872,in1);
and and16148(N26868,N26873,R0);
and and16149(N26869,R1,R2);
and and16155(N26878,N26882,N26883);
and and16156(N26879,in0,N26884);
and and16157(N26880,in2,R1);
and and16158(N26881,N26885,R3);
and and16164(N26890,N26894,N26895);
and and16165(N26891,in0,in1);
and and16166(N26892,N26896,R1);
and and16167(N26893,N26897,R3);
and and16173(N26902,N26906,N26907);
and and16174(N26903,in0,in2);
and and16175(N26904,N26908,R1);
and and16176(N26905,N26909,R3);
and and16182(N26914,N26918,N26919);
and and16183(N26915,N26920,in1);
and and16184(N26916,in2,R0);
and and16185(N26917,R1,R2);
and and16191(N26926,N26930,N26931);
and and16192(N26927,N26932,in1);
and and16193(N26928,in2,N26933);
and and16194(N26929,R1,R2);
and and16200(N26938,N26942,N26943);
and and16201(N26939,in0,in2);
and and16202(N26940,R0,N26944);
and and16203(N26941,R2,R3);
and and16209(N26950,N26954,N26955);
and and16210(N26951,in0,in1);
and and16211(N26952,N26956,R0);
and and16212(N26953,R2,R3);
and and16218(N26962,N26966,N26967);
and and16219(N26963,in0,in1);
and and16220(N26964,in2,N26968);
and and16221(N26965,R2,R3);
and and16227(N26974,N26978,N26979);
and and16228(N26975,N26980,in2);
and and16229(N26976,R0,R1);
and and16230(N26977,N26981,R3);
and and16236(N26985,N26989,N26990);
and and16237(N26986,in0,N26991);
and and16238(N26987,R0,R1);
and and16239(N26988,N26992,R3);
and and16245(N26996,N27000,N27001);
and and16246(N26997,in0,in2);
and and16247(N26998,R0,R1);
and and16248(N26999,N27002,R3);
and and16254(N27007,N27011,N27012);
and and16255(N27008,in0,in1);
and and16256(N27009,N27013,R0);
and and16257(N27010,R1,N27014);
and and16263(N27018,N27022,N27023);
and and16264(N27019,in0,in1);
and and16265(N27020,in2,N27024);
and and16266(N27021,N27025,R2);
and and16272(N27029,N27033,N27034);
and and16273(N27030,N27035,in1);
and and16274(N27031,N27036,R0);
and and16275(N27032,R2,R3);
and and16281(N27040,N27044,N27045);
and and16282(N27041,in0,in1);
and and16283(N27042,in2,R0);
and and16284(N27043,R1,R2);
and and16290(N27051,N27055,N27056);
and and16291(N27052,N27057,N27058);
and and16292(N27053,in2,R0);
and and16293(N27054,R1,R2);
and and16299(N27062,N27066,N27067);
and and16300(N27063,N27068,in1);
and and16301(N27064,N27069,R0);
and and16302(N27065,R1,R2);
and and16308(N27073,N27077,N27078);
and and16309(N27074,N27079,N27080);
and and16310(N27075,in2,R1);
and and16311(N27076,R2,R3);
and and16317(N27084,N27088,N27089);
and and16318(N27085,in0,N27090);
and and16319(N27086,in2,R0);
and and16320(N27087,R1,R2);
and and16326(N27095,N27099,N27100);
and and16327(N27096,N27101,in1);
and and16328(N27097,in2,R0);
and and16329(N27098,R1,R2);
and and16335(N27106,N27110,N27111);
and and16336(N27107,in0,in1);
and and16337(N27108,in2,R0);
and and16338(N27109,R1,R2);
and and16344(N27117,N27121,N27122);
and and16345(N27118,in0,in1);
and and16346(N27119,in2,R0);
and and16347(N27120,R1,R2);
and and16353(N27128,N27132,N27133);
and and16354(N27129,N27134,in1);
and and16355(N27130,in2,R0);
and and16356(N27131,R1,R2);
and and16362(N27139,N27143,N27144);
and and16363(N27140,in0,in1);
and and16364(N27141,in2,N27145);
and and16365(N27142,R2,R3);
and and16371(N27150,N27154,N27155);
and and16372(N27151,in0,in1);
and and16373(N27152,in2,R0);
and and16374(N27153,R1,R2);
and and16380(N27160,N27164,N27165);
and and16381(N27161,in0,in1);
and and16382(N27162,in2,R1);
and and16383(N27163,R2,N27166);
and and16389(N27170,N27174,N27175);
and and16390(N27171,in0,in2);
and and16391(N27172,R0,N27176);
and and16392(N27173,R2,R3);
and and16398(N27180,N27184,N27185);
and and16399(N27181,in1,in2);
and and16400(N27182,R0,N27186);
and and16401(N27183,R2,R3);
and and16407(N27190,N27194,N27195);
and and16408(N27191,in1,in2);
and and16409(N27192,R0,R1);
and and16410(N27193,R2,N27196);
and and16416(N27200,N27204,N27205);
and and16417(N27201,N27206,N27207);
and and16418(N27202,N27208,N27209);
and and16419(N27203,N27210,N27211);
and and16424(N27216,N27220,N27221);
and and16425(N27217,N27222,N27223);
and and16426(N27218,N27224,R3);
and and16427(N27219,N27225,N27226);
and and16432(N27232,N27236,N27237);
and and16433(N27233,N27238,N27239);
and and16434(N27234,R0,N27240);
and and16435(N27235,N27241,N27242);
and and16440(N27248,N27252,in1);
and and16441(N27249,N27253,R1);
and and16442(N27250,N27254,N27255);
and and16443(N27251,N27256,N27257);
and and16448(N27263,N27267,in0);
and and16449(N27264,N27268,R1);
and and16450(N27265,N27269,N27270);
and and16451(N27266,N27271,N27272);
and and16456(N27278,N27282,N27283);
and and16457(N27279,N27284,N27285);
and and16458(N27280,N27286,R2);
and and16459(N27281,R3,N27287);
and and16464(N27293,N27297,N27298);
and and16465(N27294,in2,N27299);
and and16466(N27295,N27300,N27301);
and and16467(N27296,N27302,N27303);
and and16472(N27308,N27312,N27313);
and and16473(N27309,N27314,N27315);
and and16474(N27310,N27316,R2);
and and16475(N27311,N27317,N27318);
and and16480(N27323,N27327,N27328);
and and16481(N27324,N27329,N27330);
and and16482(N27325,N27331,N27332);
and and16483(N27326,R4,N27333);
and and16488(N27338,N27342,N27343);
and and16489(N27339,N27344,in2);
and and16490(N27340,R0,N27345);
and and16491(N27341,N27346,N27347);
and and16496(N27353,N27357,N27358);
and and16497(N27354,in1,N27359);
and and16498(N27355,R0,N27360);
and and16499(N27356,N27361,N27362);
and and16504(N27368,N27372,N27373);
and and16505(N27369,in1,N27374);
and and16506(N27370,R1,N27375);
and and16507(N27371,N27376,N27377);
and and16512(N27383,N27387,in0);
and and16513(N27384,N27388,N27389);
and and16514(N27385,N27390,N27391);
and and16515(N27386,N27392,N27393);
and and16520(N27398,N27402,N27403);
and and16521(N27399,N27404,N27405);
and and16522(N27400,R2,N27406);
and and16523(N27401,N27407,N27408);
and and16528(N27413,N27417,N27418);
and and16529(N27414,in1,N27419);
and and16530(N27415,N27420,N27421);
and and16531(N27416,R4,N27422);
and and16536(N27427,N27431,N27432);
and and16537(N27428,in1,N27433);
and and16538(N27429,N27434,N27435);
and and16539(N27430,R3,R4);
and and16544(N27441,N27445,in0);
and and16545(N27442,N27446,N27447);
and and16546(N27443,N27448,R3);
and and16547(N27444,R4,N27449);
and and16552(N27455,N27459,in0);
and and16553(N27456,N27460,N27461);
and and16554(N27457,R2,N27462);
and and16555(N27458,R4,N27463);
and and16560(N27469,N27473,N27474);
and and16561(N27470,N27475,N27476);
and and16562(N27471,N27477,R3);
and and16563(N27472,R4,R5);
and and16568(N27483,N27487,N27488);
and and16569(N27484,in2,N27489);
and and16570(N27485,R1,R2);
and and16571(N27486,N27490,N27491);
and and16576(N27497,N27501,in1);
and and16577(N27498,N27502,N27503);
and and16578(N27499,R2,N27504);
and and16579(N27500,N27505,N27506);
and and16584(N27511,N27515,in0);
and and16585(N27512,N27516,N27517);
and and16586(N27513,R2,N27518);
and and16587(N27514,N27519,N27520);
and and16592(N27525,N27529,N27530);
and and16593(N27526,in1,N27531);
and and16594(N27527,N27532,N27533);
and and16595(N27528,R3,N27534);
and and16600(N27539,N27543,in1);
and and16601(N27540,N27544,N27545);
and and16602(N27541,R1,N27546);
and and16603(N27542,N27547,N27548);
and and16608(N27553,N27557,N27558);
and and16609(N27554,N27559,N27560);
and and16610(N27555,N27561,R3);
and and16611(N27556,N27562,R5);
and and16616(N27567,N27571,in1);
and and16617(N27568,N27572,R0);
and and16618(N27569,R1,N27573);
and and16619(N27570,N27574,N27575);
and and16624(N27581,N27585,in0);
and and16625(N27582,N27586,R0);
and and16626(N27583,R1,N27587);
and and16627(N27584,N27588,N27589);
and and16632(N27595,N27599,in1);
and and16633(N27596,N27600,N27601);
and and16634(N27597,N27602,R2);
and and16635(N27598,N27603,N27604);
and and16640(N27609,N27613,in0);
and and16641(N27610,N27614,N27615);
and and16642(N27611,N27616,R2);
and and16643(N27612,N27617,N27618);
and and16648(N27623,N27627,in0);
and and16649(N27624,N27628,R1);
and and16650(N27625,N27629,N27630);
and and16651(N27626,N27631,R5);
and and16656(N27637,N27641,in0);
and and16657(N27638,N27642,N27643);
and and16658(N27639,N27644,R3);
and and16659(N27640,N27645,R5);
and and16664(N27651,N27655,N27656);
and and16665(N27652,N27657,N27658);
and and16666(N27653,N27659,R3);
and and16667(N27654,N27660,R5);
and and16672(N27665,N27669,N27670);
and and16673(N27666,in1,N27671);
and and16674(N27667,R0,N27672);
and and16675(N27668,R4,N27673);
and and16680(N27679,N27683,N27684);
and and16681(N27680,N27685,N27686);
and and16682(N27681,R2,R3);
and and16683(N27682,N27687,N27688);
and and16688(N27693,N27697,N27698);
and and16689(N27694,N27699,N27700);
and and16690(N27695,R0,R1);
and and16691(N27696,N27701,N27702);
and and16696(N27707,N27711,in0);
and and16697(N27708,N27712,R1);
and and16698(N27709,N27713,N27714);
and and16699(N27710,N27715,R5);
and and16704(N27721,N27725,N27726);
and and16705(N27722,in1,N27727);
and and16706(N27723,N27728,R1);
and and16707(N27724,N27729,N27730);
and and16712(N27735,N27739,N27740);
and and16713(N27736,in1,N27741);
and and16714(N27737,R0,R1);
and and16715(N27738,N27742,N27743);
and and16720(N27749,N27753,N27754);
and and16721(N27750,in2,R0);
and and16722(N27751,R1,R3);
and and16723(N27752,N27755,N27756);
and and16728(N27762,N27766,N27767);
and and16729(N27763,in2,R0);
and and16730(N27764,N27768,N27769);
and and16731(N27765,R3,N27770);
and and16736(N27775,N27779,N27780);
and and16737(N27776,N27781,R0);
and and16738(N27777,N27782,R2);
and and16739(N27778,N27783,R4);
and and16744(N27788,N27792,N27793);
and and16745(N27789,in2,R0);
and and16746(N27790,N27794,N27795);
and and16747(N27791,R3,N27796);
and and16752(N27801,N27805,in0);
and and16753(N27802,N27806,R1);
and and16754(N27803,N27807,R3);
and and16755(N27804,N27808,N27809);
and and16760(N27814,N27818,N27819);
and and16761(N27815,N27820,R0);
and and16762(N27816,R1,N27821);
and and16763(N27817,R3,N27822);
and and16768(N27827,N27831,in0);
and and16769(N27828,N27832,R0);
and and16770(N27829,N27833,N27834);
and and16771(N27830,R3,N27835);
and and16776(N27840,N27844,N27845);
and and16777(N27841,N27846,in2);
and and16778(N27842,R1,R2);
and and16779(N27843,R4,N27847);
and and16784(N27853,N27857,in0);
and and16785(N27854,N27858,N27859);
and and16786(N27855,R1,N27860);
and and16787(N27856,N27861,N27862);
and and16792(N27866,N27870,in0);
and and16793(N27867,N27871,N27872);
and and16794(N27868,N27873,R3);
and and16795(N27869,N27874,R5);
and and16800(N27879,N27883,in0);
and and16801(N27880,N27884,N27885);
and and16802(N27881,N27886,R3);
and and16803(N27882,N27887,N27888);
and and16808(N27892,N27896,in0);
and and16809(N27893,N27897,N27898);
and and16810(N27894,R2,N27899);
and and16811(N27895,N27900,R5);
and and16816(N27905,N27909,in1);
and and16817(N27906,in2,N27910);
and and16818(N27907,R2,N27911);
and and16819(N27908,N27912,N27913);
and and16824(N27918,N27922,in0);
and and16825(N27919,R0,N27923);
and and16826(N27920,N27924,N27925);
and and16827(N27921,R4,N27926);
and and16832(N27931,N27935,N27936);
and and16833(N27932,in1,in2);
and and16834(N27933,N27937,R1);
and and16835(N27934,R4,N27938);
and and16840(N27944,N27948,in0);
and and16841(N27945,N27949,N27950);
and and16842(N27946,R1,N27951);
and and16843(N27947,R4,N27952);
and and16848(N27957,N27961,N27962);
and and16849(N27958,in1,in2);
and and16850(N27959,R0,N27963);
and and16851(N27960,N27964,N27965);
and and16856(N27970,N27974,in0);
and and16857(N27971,N27975,N27976);
and and16858(N27972,R1,R2);
and and16859(N27973,N27977,N27978);
and and16864(N27983,N27987,N27988);
and and16865(N27984,N27989,R0);
and and16866(N27985,R1,R2);
and and16867(N27986,N27990,N27991);
and and16872(N27996,N28000,N28001);
and and16873(N27997,N28002,R0);
and and16874(N27998,R1,N28003);
and and16875(N27999,N28004,R4);
and and16880(N28009,N28013,in0);
and and16881(N28010,N28014,N28015);
and and16882(N28011,N28016,R2);
and and16883(N28012,N28017,R4);
and and16888(N28022,N28026,in0);
and and16889(N28023,N28027,N28028);
and and16890(N28024,R1,R2);
and and16891(N28025,N28029,N28030);
and and16896(N28035,N28039,in0);
and and16897(N28036,in2,R0);
and and16898(N28037,R1,N28040);
and and16899(N28038,N28041,N28042);
and and16904(N28048,N28052,in0);
and and16905(N28049,N28053,N28054);
and and16906(N28050,R1,N28055);
and and16907(N28051,R3,N28056);
and and16912(N28061,N28065,in0);
and and16913(N28062,in1,N28066);
and and16914(N28063,N28067,R3);
and and16915(N28064,N28068,R5);
and and16920(N28074,N28078,N28079);
and and16921(N28075,in2,N28080);
and and16922(N28076,N28081,R3);
and and16923(N28077,N28082,R5);
and and16928(N28087,N28091,in0);
and and16929(N28088,N28092,N28093);
and and16930(N28089,N28094,R3);
and and16931(N28090,N28095,N28096);
and and16936(N28100,N28104,in0);
and and16937(N28101,N28105,N28106);
and and16938(N28102,R1,R2);
and and16939(N28103,N28107,N28108);
and and16944(N28113,N28117,N28118);
and and16945(N28114,N28119,R0);
and and16946(N28115,R1,N28120);
and and16947(N28116,N28121,R4);
and and16952(N28126,N28130,N28131);
and and16953(N28127,N28132,N28133);
and and16954(N28128,R0,R1);
and and16955(N28129,N28134,R3);
and and16960(N28139,N28143,in0);
and and16961(N28140,N28144,N28145);
and and16962(N28141,N28146,R2);
and and16963(N28142,N28147,R4);
and and16968(N28152,N28156,in0);
and and16969(N28153,N28157,N28158);
and and16970(N28154,N28159,N28160);
and and16971(N28155,R2,R4);
and and16976(N28165,N28169,in0);
and and16977(N28166,N28170,R1);
and and16978(N28167,R2,R3);
and and16979(N28168,R4,N28171);
and and16984(N28177,N28181,in0);
and and16985(N28178,R0,R1);
and and16986(N28179,N28182,N28183);
and and16987(N28180,N28184,R5);
and and16992(N28189,N28193,in0);
and and16993(N28190,N28194,R0);
and and16994(N28191,R1,R2);
and and16995(N28192,R3,N28195);
and and17000(N28201,N28205,in0);
and and17001(N28202,N28206,R1);
and and17002(N28203,N28207,R3);
and and17003(N28204,R4,R5);
and and17008(N28213,N28217,N28218);
and and17009(N28214,N28219,R1);
and and17010(N28215,R2,R3);
and and17011(N28216,N28220,R5);
and and17016(N28225,N28229,in0);
and and17017(N28226,in1,in2);
and and17018(N28227,N28230,N28231);
and and17019(N28228,R3,R4);
and and17024(N28237,N28241,N28242);
and and17025(N28238,in2,N28243);
and and17026(N28239,R1,R3);
and and17027(N28240,R4,N28244);
and and17032(N28249,N28253,in0);
and and17033(N28250,R0,N28254);
and and17034(N28251,N28255,R3);
and and17035(N28252,N28256,R5);
and and17040(N28261,N28265,in0);
and and17041(N28262,N28266,R1);
and and17042(N28263,N28267,R3);
and and17043(N28264,N28268,R5);
and and17048(N28273,N28277,N28278);
and and17049(N28274,in1,N28279);
and and17050(N28275,R2,R3);
and and17051(N28276,N28280,R5);
and and17056(N28285,N28289,N28290);
and and17057(N28286,in1,in2);
and and17058(N28287,R1,N28291);
and and17059(N28288,N28292,N28293);
and and17064(N28297,N28301,in0);
and and17065(N28298,in2,N28302);
and and17066(N28299,R1,N28303);
and and17067(N28300,N28304,N28305);
and and17072(N28309,N28313,in0);
and and17073(N28310,in1,in2);
and and17074(N28311,N28314,R1);
and and17075(N28312,N28315,N28316);
and and17080(N28321,N28325,N28326);
and and17081(N28322,N28327,R0);
and and17082(N28323,R1,R2);
and and17083(N28324,R3,N28328);
and and17088(N28333,N28337,in1);
and and17089(N28334,in2,N28338);
and and17090(N28335,N28339,R3);
and and17091(N28336,N28340,N28341);
and and17096(N28345,N28349,in0);
and and17097(N28346,N28350,R0);
and and17098(N28347,N28351,R2);
and and17099(N28348,N28352,N28353);
and and17104(N28357,N28361,in0);
and and17105(N28358,N28362,N28363);
and and17106(N28359,N28364,R2);
and and17107(N28360,R3,R4);
and and17112(N28369,N28373,in0);
and and17113(N28370,in1,N28374);
and and17114(N28371,R2,N28375);
and and17115(N28372,N28376,R5);
and and17120(N28381,N28385,N28386);
and and17121(N28382,N28387,N28388);
and and17122(N28383,R1,N28389);
and and17123(N28384,R3,R5);
and and17128(N28393,N28397,N28398);
and and17129(N28394,N28399,R1);
and and17130(N28395,R2,N28400);
and and17131(N28396,R4,R5);
and and17136(N28405,N28409,N28410);
and and17137(N28406,R0,R1);
and and17138(N28407,R2,N28411);
and and17139(N28408,R4,N28412);
and and17144(N28417,N28421,in0);
and and17145(N28418,N28422,N28423);
and and17146(N28419,R1,R2);
and and17147(N28420,R3,N28424);
and and17152(N28429,N28433,N28434);
and and17153(N28430,N28435,R1);
and and17154(N28431,R2,R3);
and and17155(N28432,R4,N28436);
and and17160(N28441,N28445,N28446);
and and17161(N28442,N28447,R0);
and and17162(N28443,N28448,R2);
and and17163(N28444,R4,N28449);
and and17168(N28453,N28457,N28458);
and and17169(N28454,N28459,in2);
and and17170(N28455,R0,R1);
and and17171(N28456,N28460,N28461);
and and17176(N28465,N28469,N28470);
and and17177(N28466,N28471,in2);
and and17178(N28467,R0,R1);
and and17179(N28468,R3,N28472);
and and17184(N28477,N28481,in0);
and and17185(N28478,N28482,N28483);
and and17186(N28479,R1,R2);
and and17187(N28480,R4,N28484);
and and17192(N28489,N28493,in0);
and and17193(N28490,N28494,R0);
and and17194(N28491,N28495,R2);
and and17195(N28492,N28496,R4);
and and17200(N28501,N28505,in0);
and and17201(N28502,N28506,N28507);
and and17202(N28503,R2,R3);
and and17203(N28504,R4,N28508);
and and17208(N28513,N28517,in0);
and and17209(N28514,N28518,R0);
and and17210(N28515,R1,R2);
and and17211(N28516,N28519,R5);
and and17216(N28525,N28529,N28530);
and and17217(N28526,N28531,N28532);
and and17218(N28527,R1,R2);
and and17219(N28528,R3,N28533);
and and17224(N28537,N28541,in1);
and and17225(N28538,in2,N28542);
and and17226(N28539,R2,N28543);
and and17227(N28540,R4,N28544);
and and17232(N28549,N28553,N28554);
and and17233(N28550,N28555,in2);
and and17234(N28551,R0,N28556);
and and17235(N28552,R3,R4);
and and17240(N28561,N28565,in2);
and and17241(N28562,R0,N28566);
and and17242(N28563,N28567,R3);
and and17243(N28564,N28568,R5);
and and17248(N28573,N28577,in0);
and and17249(N28574,R0,R1);
and and17250(N28575,N28578,R3);
and and17251(N28576,N28579,N28580);
and and17256(N28585,N28589,in0);
and and17257(N28586,N28590,N28591);
and and17258(N28587,N28592,R2);
and and17259(N28588,R3,R4);
and and17264(N28597,N28601,N28602);
and and17265(N28598,N28603,N28604);
and and17266(N28599,R0,R1);
and and17267(N28600,R2,R3);
and and17272(N28609,N28613,in1);
and and17273(N28610,N28614,R0);
and and17274(N28611,R1,N28615);
and and17275(N28612,R3,R4);
and and17280(N28621,N28625,in0);
and and17281(N28622,in1,R0);
and and17282(N28623,N28626,N28627);
and and17283(N28624,R4,R5);
and and17288(N28633,N28637,N28638);
and and17289(N28634,N28639,in2);
and and17290(N28635,R0,R1);
and and17291(N28636,R2,R4);
and and17296(N28645,N28649,N28650);
and and17297(N28646,N28651,R0);
and and17298(N28647,R1,R2);
and and17299(N28648,N28652,R4);
and and17304(N28657,N28661,in0);
and and17305(N28658,in1,in2);
and and17306(N28659,R0,R1);
and and17307(N28660,R3,N28662);
and and17312(N28668,N28672,in0);
and and17313(N28669,in2,R0);
and and17314(N28670,R1,R3);
and and17315(N28671,R4,N28673);
and and17320(N28679,N28683,in0);
and and17321(N28680,N28684,N28685);
and and17322(N28681,R1,R3);
and and17323(N28682,R4,N28686);
and and17328(N28690,N28694,in1);
and and17329(N28691,N28695,R1);
and and17330(N28692,N28696,R3);
and and17331(N28693,R4,N28697);
and and17336(N28701,N28705,N28706);
and and17337(N28702,in1,in2);
and and17338(N28703,R0,N28707);
and and17339(N28704,R2,R4);
and and17344(N28712,N28716,in0);
and and17345(N28713,N28717,R0);
and and17346(N28714,R2,R3);
and and17347(N28715,N28718,R5);
and and17352(N28723,N28727,in1);
and and17353(N28724,R0,N28728);
and and17354(N28725,R2,N28729);
and and17355(N28726,R4,R5);
and and17360(N28734,N28738,in0);
and and17361(N28735,N28739,R0);
and and17362(N28736,R1,R2);
and and17363(N28737,R3,N28740);
and and17368(N28745,N28749,in0);
and and17369(N28746,in1,R0);
and and17370(N28747,N28750,R2);
and and17371(N28748,R3,N28751);
and and17376(N28756,N28760,in1);
and and17377(N28757,R0,R1);
and and17378(N28758,R2,N28761);
and and17379(N28759,R4,N28762);
and and17384(N28767,N28771,in0);
and and17385(N28768,R0,R1);
and and17386(N28769,R2,N28772);
and and17387(N28770,R4,N28773);
and and17392(N28778,N28782,in0);
and and17393(N28779,N28783,R1);
and and17394(N28780,N28784,R3);
and and17395(N28781,R4,R5);
and and17400(N28789,N28793,in0);
and and17401(N28790,N28794,N28795);
and and17402(N28791,R1,R2);
and and17403(N28792,N28796,R4);
and and17408(N28800,N28804,N28805);
and and17409(N28801,in1,in2);
and and17410(N28802,R0,R1);
and and17411(N28803,N28806,R4);
and and17416(N28811,N28815,N28816);
and and17417(N28812,in1,R0);
and and17418(N28813,R1,R3);
and and17419(N28814,N28817,N28818);
and and17424(N28822,N28826,in0);
and and17425(N28823,in1,in2);
and and17426(N28824,N28827,R1);
and and17427(N28825,N28828,N28829);
and and17432(N28833,N28837,in0);
and and17433(N28834,N28838,R0);
and and17434(N28835,R1,N28839);
and and17435(N28836,R4,R5);
and and17440(N28844,N28848,in0);
and and17441(N28845,in1,N28849);
and and17442(N28846,R0,R1);
and and17443(N28847,R2,R3);
and and17448(N28855,N28859,in0);
and and17449(N28856,in1,R0);
and and17450(N28857,R2,N28860);
and and17451(N28858,N28861,R5);
and and17456(N28866,N28870,in0);
and and17457(N28867,in2,N28871);
and and17458(N28868,R1,R2);
and and17459(N28869,R3,N28872);
and and17464(N28877,N28881,in0);
and and17465(N28878,in2,R0);
and and17466(N28879,R1,N28882);
and and17467(N28880,N28883,R4);
and and17472(N28888,N28892,in2);
and and17473(N28889,N28893,R1);
and and17474(N28890,R2,R3);
and and17475(N28891,R4,N28894);
and and17480(N28899,N28903,in0);
and and17481(N28900,in1,in2);
and and17482(N28901,N28904,R2);
and and17483(N28902,R3,N28905);
and and17488(N28910,N28914,N28915);
and and17489(N28911,N28916,N28917);
and and17490(N28912,R1,R3);
and and17491(N28913,R4,R5);
and and17496(N28921,N28925,in0);
and and17497(N28922,N28926,N28927);
and and17498(N28923,R1,R2);
and and17499(N28924,N28928,R4);
and and17504(N28932,N28936,in0);
and and17505(N28933,in2,N28937);
and and17506(N28934,R2,R3);
and and17507(N28935,R4,R5);
and and17512(N28942,N28946,in0);
and and17513(N28943,R0,R1);
and and17514(N28944,R2,N28947);
and and17515(N28945,R4,R5);
and and17520(N28952,N28956,in0);
and and17521(N28953,N28957,N28958);
and and17522(N28954,R2,R3);
and and17523(N28955,R4,R5);
and and17528(N28962,N28966,N28967);
and and17529(N28963,in1,in2);
and and17530(N28964,N28968,R1);
and and17531(N28965,R3,R5);
and and17536(N28972,N28976,in0);
and and17537(N28973,R0,N28977);
and and17538(N28974,R2,R3);
and and17539(N28975,N28978,R5);
and and17544(N28982,N28986,in0);
and and17545(N28983,R0,R1);
and and17546(N28984,R2,R3);
and and17547(N28985,N28987,N28988);
and and17552(N28992,N28996,N28997);
and and17553(N28993,N28998,in2);
and and17554(N28994,R0,R1);
and and17555(N28995,R2,R5);
and and17560(N29002,N29006,in0);
and and17561(N29003,R0,N29007);
and and17562(N29004,R2,R3);
and and17563(N29005,R4,R5);
and and17568(N29012,N29016,in1);
and and17569(N29013,N29017,R0);
and and17570(N29014,R1,R2);
and and17571(N29015,N29018,R4);
and and17576(N29022,N29026,in0);
and and17577(N29023,R0,R1);
and and17578(N29024,R2,R3);
and and17579(N29025,N29027,R5);
and and17584(N29032,N29036,in0);
and and17585(N29033,N29037,R0);
and and17586(N29034,R1,R2);
and and17587(N29035,N29038,R4);
and and17592(N29042,N29046,in0);
and and17593(N29043,N29047,R1);
and and17594(N29044,R2,R3);
and and17595(N29045,R4,N29048);
and and17600(N29052,N29056,in0);
and and17601(N29053,in1,in2);
and and17602(N29054,R0,R1);
and and17603(N29055,N29057,R3);
and and17608(N29061,N29065,N29066);
and and17609(N29062,N29067,N29068);
and and17610(N29063,R4,R5);
and and17611(N29064,N29069,N29070);
and and17615(N29074,in0,N29078);
and and17616(N29075,N29079,N29080);
and and17617(N29076,N29081,N29082);
and and17618(N29077,R6,N29083);
and and17622(N29087,in0,N29091);
and and17623(N29088,N29092,N29093);
and and17624(N29089,N29094,N29095);
and and17625(N29090,R6,N29096);
and and17629(N29100,in0,N29104);
and and17630(N29101,R1,N29105);
and and17631(N29102,R3,N29106);
and and17632(N29103,N29107,N29108);
and and17636(N29112,N29116,R0);
and and17637(N29113,R1,N29117);
and and17638(N29114,R3,N29118);
and and17639(N29115,N29119,N29120);
and and17643(N29124,in0,N29128);
and and17644(N29125,R1,R2);
and and17645(N29126,N29129,N29130);
and and17646(N29127,N29131,N29132);
and and17650(N29136,in0,R0);
and and17651(N29137,N29140,N29141);
and and17652(N29138,N29142,N29143);
and and17653(N29139,R6,N29144);
and and17657(N29148,R0,N29152);
and and17658(N29149,N29153,N29154);
and and17659(N29150,R4,R5);
and and17660(N29151,N29155,N29156);
and and17664(N29160,in0,in1);
and and17665(N29161,N29164,R2);
and and17666(N29162,R3,N29165);
and and17667(N29163,N29166,N29167);
and and17671(N29171,in0,N29175);
and and17672(N29172,R2,R3);
and and17673(N29173,N29176,N29177);
and and17674(N29174,R6,N29178);
and and17678(N29182,in0,R0);
and and17679(N29183,R2,N29186);
and and17680(N29184,R4,N29187);
and and17681(N29185,N29188,N29189);
and and17685(N29193,in0,N29197);
and and17686(N29194,N29198,R3);
and and17687(N29195,R4,N29199);
and and17688(N29196,N29200,R7);
and and17692(N29204,in0,R0);
and and17693(N29205,N29208,N29209);
and and17694(N29206,R3,R4);
and and17695(N29207,N29210,N29211);
and and17699(N29215,in0,N29219);
and and17700(N29216,R1,N29220);
and and17701(N29217,N29221,R4);
and and17702(N29218,R6,N29222);
and and17706(N29226,in0,N29230);
and and17707(N29227,R1,N29231);
and and17708(N29228,N29232,R4);
and and17709(N29229,R6,N29233);
and and17713(N29237,in0,N29241);
and and17714(N29238,R0,R1);
and and17715(N29239,N29242,R5);
and and17716(N29240,N29243,R7);
and and17720(N29247,in0,R0);
and and17721(N29248,N29251,R2);
and and17722(N29249,R4,N29252);
and and17723(N29250,N29253,R7);
and and17727(N29257,in0,R0);
and and17728(N29258,R1,N29261);
and and17729(N29259,R3,R4);
and and17730(N29260,R5,N29262);
and and17734(N29266,R0,N29269);
and and17735(N29267,N29270,R4);
and and17736(N29268,N29271,N29272);
and and14584(N24434,N24441,R5);
and and14585(N24435,N24442,N24443);
and and14593(N24451,N24457,N24458);
and and14594(N24452,N24459,N24460);
and and14602(N24468,N24475,R4);
and and14603(N24469,N24476,N24477);
and and14611(N24485,N24491,N24492);
and and14612(N24486,N24493,N24494);
and and14620(N24502,N24508,N24509);
and and14621(N24503,N24510,N24511);
and and14629(N24519,R4,N24526);
and and14630(N24520,N24527,N24528);
and and14638(N24536,N24543,N24544);
and and14639(N24537,N24545,R7);
and and14647(N24553,R3,N24560);
and and14648(N24554,N24561,N24562);
and and14656(N24570,R4,N24576);
and and14657(N24571,N24577,N24578);
and and14665(N24586,N24592,N24593);
and and14666(N24587,N24594,R7);
and and14674(N24602,N24608,N24609);
and and14675(N24603,N24610,R7);
and and14683(N24618,R4,N24624);
and and14684(N24619,N24625,N24626);
and and14692(N24634,N24640,N24641);
and and14693(N24635,N24642,R7);
and and14701(N24650,N24655,N24656);
and and14702(N24651,N24657,N24658);
and and14710(N24666,N24672,R5);
and and14711(N24667,N24673,N24674);
and and14719(N24682,N24689,R5);
and and14720(N24683,N24690,R7);
and and14728(N24698,R4,N24705);
and and14729(N24699,R6,N24706);
and and14737(N24714,N24721,R5);
and and14738(N24715,R6,N24722);
and and14746(N24730,N24736,R5);
and and14747(N24731,N24737,N24738);
and and14755(N24746,R4,N24752);
and and14756(N24747,N24753,N24754);
and and14764(N24762,N24768,N24769);
and and14765(N24763,N24770,R7);
and and14773(N24778,N24784,N24785);
and and14774(N24779,N24786,R7);
and and14782(N24794,N24799,N24800);
and and14783(N24795,N24801,N24802);
and and14791(N24810,N24816,N24817);
and and14792(N24811,N24818,R7);
and and14800(N24826,N24832,N24833);
and and14801(N24827,N24834,R7);
and and14809(N24842,N24847,N24848);
and and14810(N24843,N24849,N24850);
and and14818(N24858,N24864,R5);
and and14819(N24859,N24865,N24866);
and and14827(N24874,N24878,N24879);
and and14828(N24875,N24880,N24881);
and and14836(N24889,N24895,N24896);
and and14837(N24890,R6,R7);
and and14845(N24904,N24909,R5);
and and14846(N24905,N24910,N24911);
and and14854(N24919,R4,N24924);
and and14855(N24920,N24925,N24926);
and and14863(N24934,R4,N24940);
and and14864(N24935,R6,N24941);
and and14872(N24949,N24955,R4);
and and14873(N24950,R5,N24956);
and and14881(N24964,R4,N24970);
and and14882(N24965,N24971,R7);
and and14890(N24979,R3,R4);
and and14891(N24980,N24986,R6);
and and14899(N24994,R4,R5);
and and14900(N24995,N25000,N25001);
and and14908(N25009,R4,R5);
and and14909(N25010,N25015,N25016);
and and14917(N25024,R3,N25029);
and and14918(N25025,N25030,N25031);
and and14926(N25039,N25044,N25045);
and and14927(N25040,R6,N25046);
and and14935(N25054,N25060,R5);
and and14936(N25055,N25061,R7);
and and14944(N25069,N25075,N25076);
and and14945(N25070,R6,R7);
and and14953(N25084,R4,N25090);
and and14954(N25085,R6,N25091);
and and14962(N25099,R4,N25105);
and and14963(N25100,R6,N25106);
and and14971(N25114,N25120,R5);
and and14972(N25115,R6,N25121);
and and14980(N25129,R3,R5);
and and14981(N25130,N25135,N25136);
and and14989(N25144,N25149,R5);
and and14990(N25145,N25150,N25151);
and and14998(N25159,R4,N25165);
and and14999(N25160,N25166,R7);
and and15007(N25174,R4,N25181);
and and15008(N25175,R6,R7);
and and15016(N25189,R3,N25196);
and and15017(N25190,R6,R7);
and and15025(N25204,R3,N25210);
and and15026(N25205,N25211,R7);
and and15034(N25219,N25224,R5);
and and15035(N25220,N25225,N25226);
and and15043(N25234,N25239,R5);
and and15044(N25235,N25240,N25241);
and and15052(N25249,R4,R5);
and and15053(N25250,N25255,N25256);
and and15061(N25264,N25269,R5);
and and15062(N25265,R6,N25270);
and and15070(N25278,N25282,N25283);
and and15071(N25279,N25284,R7);
and and15079(N25292,R3,R4);
and and15080(N25293,N25297,N25298);
and and15088(N25306,R4,R5);
and and15089(N25307,N25311,N25312);
and and15097(N25320,R4,N25325);
and and15098(N25321,N25326,R7);
and and15106(N25334,N25339,N25340);
and and15107(N25335,R6,R7);
and and15115(N25348,N25353,R5);
and and15116(N25349,R6,N25354);
and and15124(N25362,R4,R5);
and and15125(N25363,N25367,N25368);
and and15133(N25376,N25380,N25381);
and and15134(N25377,N25382,R7);
and and15142(N25390,N25394,N25395);
and and15143(N25391,R6,N25396);
and and15151(N25404,N25408,N25409);
and and15152(N25405,R6,N25410);
and and15160(N25418,R3,N25423);
and and15161(N25419,N25424,R7);
and and15169(N25432,R3,N25437);
and and15170(N25433,N25438,R7);
and and15178(N25446,R4,N25452);
and and15179(N25447,R6,R7);
and and15187(N25460,R4,R5);
and and15188(N25461,N25465,N25466);
and and15196(N25474,R3,R5);
and and15197(N25475,R6,N25480);
and and15205(N25488,R4,R5);
and and15206(N25489,N25494,R7);
and and15214(N25502,R4,R5);
and and15215(N25503,R6,N25508);
and and15223(N25516,N25520,N25521);
and and15224(N25517,R6,N25522);
and and15232(N25530,N25535,R5);
and and15233(N25531,N25536,R7);
and and15241(N25544,N25549,R5);
and and15242(N25545,N25550,R7);
and and15250(N25558,N25562,R5);
and and15251(N25559,N25563,N25564);
and and15259(N25572,R4,R5);
and and15260(N25573,N25578,R7);
and and15268(N25586,N25590,N25591);
and and15269(N25587,N25592,R7);
and and15277(N25600,N25604,R5);
and and15278(N25601,N25605,N25606);
and and15286(N25614,R3,N25619);
and and15287(N25615,R5,N25620);
and and15295(N25628,R4,N25634);
and and15296(N25629,R6,R7);
and and15304(N25642,N25646,R5);
and and15305(N25643,N25647,N25648);
and and15313(N25656,N25661,R5);
and and15314(N25657,N25662,R7);
and and15322(N25670,N25674,N25675);
and and15323(N25671,R6,N25676);
and and15331(N25684,N25689,R5);
and and15332(N25685,N25690,R7);
and and15340(N25698,N25703,N25704);
and and15341(N25699,R6,R7);
and and15349(N25712,N25717,R5);
and and15350(N25713,N25718,R7);
and and15358(N25726,N25731,R5);
and and15359(N25727,N25732,R7);
and and15367(N25740,R4,R5);
and and15368(N25741,N25746,R7);
and and15376(N25754,R4,R5);
and and15377(N25755,N25760,R7);
and and15385(N25768,N25773,R5);
and and15386(N25769,N25774,R7);
and and15394(N25782,N25787,R5);
and and15395(N25783,R6,N25788);
and and15403(N25796,N25800,R5);
and and15404(N25797,N25801,N25802);
and and15412(N25810,R4,N25816);
and and15413(N25811,R6,R7);
and and15421(N25824,R3,N25829);
and and15422(N25825,R5,N25830);
and and15430(N25838,N25842,N25843);
and and15431(N25839,N25844,R7);
and and15439(N25852,R4,N25856);
and and15440(N25853,N25857,N25858);
and and15448(N25866,R3,R4);
and and15449(N25867,R6,N25872);
and and15457(N25880,R4,N25885);
and and15458(N25881,N25886,R7);
and and15466(N25894,R4,R5);
and and15467(N25895,N25900,R7);
and and15475(N25908,R4,N25914);
and and15476(N25909,R6,R7);
and and15484(N25922,R4,N25928);
and and15485(N25923,R6,R7);
and and15493(N25936,N25941,N25942);
and and15494(N25937,R6,R7);
and and15502(N25950,R3,N25955);
and and15503(N25951,N25956,R7);
and and15511(N25964,N25968,N25969);
and and15512(N25965,N25970,R7);
and and15520(N25978,N25982,R5);
and and15521(N25979,N25983,N25984);
and and15529(N25992,N25996,N25997);
and and15530(N25993,R6,N25998);
and and15538(N26006,N26010,N26011);
and and15539(N26007,N26012,R7);
and and15547(N26020,R4,R5);
and and15548(N26021,N26025,N26026);
and and15556(N26034,R3,R4);
and and15557(N26035,R5,N26040);
and and15565(N26048,N26053,R4);
and and15566(N26049,R5,N26054);
and and15574(N26062,N26066,R5);
and and15575(N26063,N26067,N26068);
and and15583(N26076,N26080,R5);
and and15584(N26077,N26081,N26082);
and and15592(N26090,N26094,R5);
and and15593(N26091,N26095,N26096);
and and15601(N26104,R4,R5);
and and15602(N26105,N26109,N26110);
and and15610(N26118,R4,N26123);
and and15611(N26119,N26124,R7);
and and15619(N26132,R4,N26137);
and and15620(N26133,N26138,R7);
and and15628(N26146,R3,N26149);
and and15629(N26147,N26150,N26151);
and and15637(N26159,R3,N26163);
and and15638(N26160,R6,N26164);
and and15646(N26172,N26176,R5);
and and15647(N26173,N26177,R7);
and and15655(N26185,R4,R5);
and and15656(N26186,R6,N26190);
and and15664(N26198,R4,N26202);
and and15665(N26199,R6,N26203);
and and15673(N26211,N26215,N26216);
and and15674(N26212,R6,R7);
and and15682(N26224,R4,R5);
and and15683(N26225,N26229,R7);
and and15691(N26237,N26241,R5);
and and15692(N26238,R6,N26242);
and and15700(N26250,N26254,R5);
and and15701(N26251,N26255,R7);
and and15709(N26263,R4,R5);
and and15710(N26264,R6,N26268);
and and15718(N26276,N26280,N26281);
and and15719(N26277,R6,R7);
and and15727(N26289,R3,R4);
and and15728(N26290,R5,N26294);
and and15736(N26302,N26305,R5);
and and15737(N26303,N26306,N26307);
and and15745(N26315,R4,N26320);
and and15746(N26316,R6,R7);
and and15754(N26328,R4,N26333);
and and15755(N26329,R6,R7);
and and15763(N26341,R3,R4);
and and15764(N26342,R6,N26346);
and and15772(N26354,R3,R4);
and and15773(N26355,R6,N26359);
and and15781(N26367,R3,R4);
and and15782(N26368,N26372,R6);
and and15790(N26380,R4,N26384);
and and15791(N26381,R6,N26385);
and and15799(N26393,N26398,R5);
and and15800(N26394,R6,R7);
and and15808(N26406,N26410,N26411);
and and15809(N26407,R6,R7);
and and15817(N26419,N26423,R4);
and and15818(N26420,N26424,R6);
and and15826(N26432,R4,R5);
and and15827(N26433,N26437,R7);
and and15835(N26445,R4,R5);
and and15836(N26446,N26450,R7);
and and15844(N26458,N26461,N26462);
and and15845(N26459,N26463,R7);
and and15853(N26471,R4,N26475);
and and15854(N26472,R6,N26476);
and and15862(N26484,N26487,R5);
and and15863(N26485,N26488,N26489);
and and15871(N26497,R3,R4);
and and15872(N26498,N26502,R7);
and and15880(N26510,R4,R5);
and and15881(N26511,N26514,R7);
and and15889(N26522,N26525,R5);
and and15890(N26523,R6,N26526);
and and15898(N26534,R3,R5);
and and15899(N26535,R6,N26538);
and and15907(N26546,R4,R5);
and and15908(N26547,N26550,R7);
and and15916(N26558,N26561,R5);
and and15917(N26559,N26562,R7);
and and15925(N26570,R4,N26574);
and and15926(N26571,R6,R7);
and and15934(N26582,N26585,R5);
and and15935(N26583,R6,N26586);
and and15943(N26594,N26597,R4);
and and15944(N26595,R5,N26598);
and and15952(N26606,R3,N26609);
and and15953(N26607,R6,N26610);
and and15961(N26618,R4,R5);
and and15962(N26619,N26622,R7);
and and15970(N26630,R4,R5);
and and15971(N26631,R6,N26634);
and and15979(N26642,R4,R5);
and and15980(N26643,R6,N26646);
and and15988(N26654,R4,R5);
and and15989(N26655,R6,N26658);
and and15997(N26666,N26669,R5);
and and15998(N26667,N26670,R7);
and and16006(N26678,R4,N26681);
and and16007(N26679,N26682,R7);
and and16015(N26690,N26692,N26693);
and and16016(N26691,N26694,R7);
and and16024(N26702,N26705,R5);
and and16025(N26703,N26706,R7);
and and16033(N26714,R4,R5);
and and16034(N26715,N26717,N26718);
and and16042(N26726,N26729,R5);
and and16043(N26727,N26730,R7);
and and16051(N26738,R4,R5);
and and16052(N26739,R6,R7);
and and16060(N26750,R3,R5);
and and16061(N26751,N26754,R7);
and and16069(N26762,R4,R5);
and and16070(N26763,N26766,R7);
and and16078(N26774,R4,R5);
and and16079(N26775,N26777,N26778);
and and16087(N26786,R4,R5);
and and16088(N26787,R6,N26790);
and and16096(N26798,N26800,R5);
and and16097(N26799,N26801,N26802);
and and16105(N26810,R4,R5);
and and16106(N26811,R6,N26814);
and and16114(N26822,R4,N26825);
and and16115(N26823,R6,N26826);
and and16123(N26834,R4,N26838);
and and16124(N26835,R6,R7);
and and16132(N26846,R4,R5);
and and16133(N26847,R6,N26850);
and and16141(N26858,R4,R5);
and and16142(N26859,R6,N26862);
and and16150(N26870,N26874,R5);
and and16151(N26871,R6,R7);
and and16159(N26882,R4,R5);
and and16160(N26883,N26886,R7);
and and16168(N26894,R4,R5);
and and16169(N26895,N26898,R7);
and and16177(N26906,R4,R5);
and and16178(N26907,R6,N26910);
and and16186(N26918,N26921,R4);
and and16187(N26919,R5,N26922);
and and16195(N26930,R3,R5);
and and16196(N26931,R6,N26934);
and and16204(N26942,R4,R5);
and and16205(N26943,N26945,N26946);
and and16213(N26954,R4,R5);
and and16214(N26955,N26957,N26958);
and and16222(N26966,R4,N26969);
and and16223(N26967,N26970,R7);
and and16231(N26978,R4,R5);
and and16232(N26979,R6,R7);
and and16240(N26989,R4,R5);
and and16241(N26990,R6,R7);
and and16249(N27000,R4,N27003);
and and16250(N27001,R6,R7);
and and16258(N27011,R3,R4);
and and16259(N27012,R6,R7);
and and16267(N27022,R3,R4);
and and16268(N27023,R5,R6);
and and16276(N27033,R4,R5);
and and16277(N27034,R6,R7);
and and16285(N27044,N27046,R4);
and and16286(N27045,N27047,R6);
and and16294(N27055,R3,R4);
and and16295(N27056,R5,R7);
and and16303(N27066,R3,R4);
and and16304(N27067,R5,R7);
and and16312(N27077,R4,R5);
and and16313(N27078,R6,R7);
and and16321(N27088,N27091,R4);
and and16322(N27089,R6,R7);
and and16330(N27099,R3,R4);
and and16331(N27100,N27102,R6);
and and16339(N27110,R3,R4);
and and16340(N27111,N27112,N27113);
and and16348(N27121,R3,R4);
and and16349(N27122,N27123,N27124);
and and16357(N27132,R3,N27135);
and and16358(N27133,R5,R7);
and and16366(N27143,R4,R5);
and and16367(N27144,R6,N27146);
and and16375(N27154,N27156,R4);
and and16376(N27155,R5,R7);
and and16384(N27164,R4,R5);
and and16385(N27165,R6,R7);
and and16393(N27174,R4,R5);
and and16394(N27175,R6,R7);
and and16402(N27184,R4,R5);
and and16403(N27185,R6,R7);
and and16411(N27194,R4,R5);
and and16412(N27195,R6,R7);
and and16420(N27204,N27212,R7);
and and16428(N27220,N27227,N27228);
and and16436(N27236,N27243,N27244);
and and16444(N27252,N27258,N27259);
and and16452(N27267,N27273,N27274);
and and16460(N27282,N27288,N27289);
and and16468(N27297,R6,N27304);
and and16476(N27312,R6,N27319);
and and16484(N27327,R6,N27334);
and and16492(N27342,N27348,N27349);
and and16500(N27357,N27363,N27364);
and and16508(N27372,N27378,N27379);
and and16516(N27387,N27394,R7);
and and16524(N27402,R6,N27409);
and and16532(N27417,N27423,R7);
and and16540(N27431,N27436,N27437);
and and16548(N27445,N27450,N27451);
and and16556(N27459,N27464,N27465);
and and16564(N27473,N27478,N27479);
and and16572(N27487,N27492,N27493);
and and16580(N27501,N27507,R7);
and and16588(N27515,N27521,R7);
and and16596(N27529,R6,N27535);
and and16604(N27543,R6,N27549);
and and16612(N27557,N27563,R7);
and and16620(N27571,N27576,N27577);
and and16628(N27585,N27590,N27591);
and and16636(N27599,R6,N27605);
and and16644(N27613,R6,N27619);
and and16652(N27627,N27632,N27633);
and and16660(N27641,N27646,N27647);
and and16668(N27655,R6,N27661);
and and16676(N27669,N27674,N27675);
and and16684(N27683,N27689,R7);
and and16692(N27697,N27703,R6);
and and16700(N27711,N27716,N27717);
and and16708(N27725,R6,N27731);
and and16716(N27739,N27744,N27745);
and and16724(N27753,N27757,N27758);
and and16732(N27766,R5,N27771);
and and16740(N27779,R6,N27784);
and and16748(N27792,R6,N27797);
and and16756(N27805,N27810,R7);
and and16764(N27818,N27823,R7);
and and16772(N27831,N27836,R7);
and and16780(N27844,N27848,N27849);
and and16788(N27857,R6,R7);
and and16796(N27870,N27875,R7);
and and16804(N27883,R6,R7);
and and16812(N27896,N27901,R7);
and and16820(N27909,R6,N27914);
and and16828(N27922,R6,N27927);
and and16836(N27935,N27939,N27940);
and and16844(N27948,N27953,R7);
and and16852(N27961,N27966,R7);
and and16860(N27974,N27979,R6);
and and16868(N27987,N27992,R7);
and and16876(N28000,R5,N28005);
and and16884(N28013,N28018,R7);
and and16892(N28026,R5,N28031);
and and16900(N28039,N28043,N28044);
and and16908(N28052,N28057,R7);
and and16916(N28065,N28069,N28070);
and and16924(N28078,R6,N28083);
and and16932(N28091,R6,R7);
and and16940(N28104,N28109,R6);
and and16948(N28117,R5,N28122);
and and16956(N28130,N28135,R7);
and and16964(N28143,N28148,R7);
and and16972(N28156,N28161,R7);
and and16980(N28169,N28172,N28173);
and and16988(N28181,R6,N28185);
and and16996(N28193,N28196,N28197);
and and17004(N28205,N28208,N28209);
and and17012(N28217,N28221,R7);
and and17020(N28229,N28232,N28233);
and and17028(N28241,R6,N28245);
and and17036(N28253,R6,N28257);
and and17044(N28265,R6,N28269);
and and17052(N28277,R6,N28281);
and and17060(N28289,R6,R7);
and and17068(N28301,R6,R7);
and and17076(N28313,N28317,R6);
and and17084(N28325,R6,N28329);
and and17092(N28337,R6,R7);
and and17100(N28349,R6,R7);
and and17108(N28361,R5,N28365);
and and17116(N28373,N28377,R7);
and and17124(N28385,R6,R7);
and and17132(N28397,R6,N28401);
and and17140(N28409,R6,N28413);
and and17148(N28421,N28425,R7);
and and17156(N28433,R6,N28437);
and and17164(N28445,R6,R7);
and and17172(N28457,R6,R7);
and and17180(N28469,R5,N28473);
and and17188(N28481,R6,N28485);
and and17196(N28493,R5,N28497);
and and17204(N28505,R6,N28509);
and and17212(N28517,N28520,N28521);
and and17220(N28529,R5,R6);
and and17228(N28541,N28545,R7);
and and17236(N28553,N28557,R7);
and and17244(N28565,N28569,R7);
and and17252(N28577,N28581,R7);
and and17260(N28589,R5,N28593);
and and17268(N28601,N28605,R6);
and and17276(N28613,N28616,N28617);
and and17284(N28625,N28628,N28629);
and and17292(N28637,N28640,N28641);
and and17300(N28649,N28653,R6);
and and17308(N28661,N28663,N28664);
and and17316(N28672,N28674,N28675);
and and17324(N28683,R6,R7);
and and17332(N28694,R6,R7);
and and17340(N28705,R6,N28708);
and and17348(N28716,R6,N28719);
and and17356(N28727,N28730,R7);
and and17364(N28738,N28741,R7);
and and17372(N28749,R5,N28752);
and and17380(N28760,N28763,R7);
and and17388(N28771,N28774,R7);
and and17396(N28782,R6,N28785);
and and17404(N28793,R5,R7);
and and17412(N28804,R5,N28807);
and and17420(N28815,R6,R7);
and and17428(N28826,R6,R7);
and and17436(N28837,N28840,R7);
and and17444(N28848,N28850,N28851);
and and17452(N28859,N28862,R7);
and and17460(N28870,N28873,R7);
and and17468(N28881,R6,N28884);
and and17476(N28892,R6,N28895);
and and17484(N28903,N28906,R6);
and and17492(N28914,R6,R7);
and and17500(N28925,R5,R7);
and and17508(N28936,N28938,R7);
and and17516(N28946,R6,N28948);
and and17524(N28956,R6,R7);
and and17532(N28966,R6,R7);
and and17540(N28976,R6,R7);
and and17548(N28986,R6,R7);
and and17556(N28996,R6,R7);
and and17564(N29006,N29008,R7);
and and17572(N29016,R6,R7);
and and17580(N29026,R6,N29028);
and and17588(N29036,R5,R6);
and and17596(N29046,R6,R7);
and and17604(N29056,R4,R5);
and and17737(N29434,N29435,N29436);
and and17747(N29452,N29453,N29454);
and and17757(N29470,N29471,N29472);
and and17767(N29487,N29488,N29489);
and and17777(N29504,N29505,N29506);
and and17787(N29520,N29521,N29522);
and and17797(N29536,N29537,N29538);
and and17807(N29550,N29551,N29552);
and and17816(N29568,N29569,N29570);
and and17825(N29586,N29587,N29588);
and and17834(N29604,N29605,N29606);
and and17843(N29621,N29622,N29623);
and and17852(N29638,N29639,N29640);
and and17861(N29655,N29656,N29657);
and and17870(N29672,N29673,N29674);
and and17879(N29689,N29690,N29691);
and and17888(N29706,N29707,N29708);
and and17897(N29722,N29723,N29724);
and and17906(N29738,N29739,N29740);
and and17915(N29754,N29755,N29756);
and and17924(N29770,N29771,N29772);
and and17933(N29786,N29787,N29788);
and and17942(N29802,N29803,N29804);
and and17951(N29818,N29819,N29820);
and and17960(N29834,N29835,N29836);
and and17969(N29850,N29851,N29852);
and and17978(N29866,N29867,N29868);
and and17987(N29882,N29883,N29884);
and and17996(N29898,N29899,N29900);
and and18005(N29914,N29915,N29916);
and and18014(N29930,N29931,N29932);
and and18023(N29946,N29947,N29948);
and and18032(N29962,N29963,N29964);
and and18041(N29978,N29979,N29980);
and and18050(N29994,N29995,N29996);
and and18059(N30009,N30010,N30011);
and and18068(N30024,N30025,N30026);
and and18077(N30039,N30040,N30041);
and and18086(N30054,N30055,N30056);
and and18095(N30069,N30070,N30071);
and and18104(N30084,N30085,N30086);
and and18113(N30099,N30100,N30101);
and and18122(N30114,N30115,N30116);
and and18131(N30129,N30130,N30131);
and and18140(N30144,N30145,N30146);
and and18149(N30159,N30160,N30161);
and and18158(N30174,N30175,N30176);
and and18167(N30189,N30190,N30191);
and and18176(N30204,N30205,N30206);
and and18185(N30219,N30220,N30221);
and and18194(N30234,N30235,N30236);
and and18203(N30249,N30250,N30251);
and and18212(N30264,N30265,N30266);
and and18221(N30279,N30280,N30281);
and and18230(N30294,N30295,N30296);
and and18239(N30309,N30310,N30311);
and and18248(N30324,N30325,N30326);
and and18257(N30339,N30340,N30341);
and and18266(N30354,N30355,N30356);
and and18275(N30369,N30370,N30371);
and and18284(N30384,N30385,N30386);
and and18293(N30399,N30400,N30401);
and and18302(N30414,N30415,N30416);
and and18311(N30429,N30430,N30431);
and and18320(N30444,N30445,N30446);
and and18329(N30459,N30460,N30461);
and and18338(N30474,N30475,N30476);
and and18347(N30488,N30489,N30490);
and and18356(N30502,N30503,N30504);
and and18365(N30516,N30517,N30518);
and and18374(N30530,N30531,N30532);
and and18383(N30544,N30545,N30546);
and and18392(N30558,N30559,N30560);
and and18401(N30572,N30573,N30574);
and and18410(N30586,N30587,N30588);
and and18419(N30600,N30601,N30602);
and and18428(N30614,N30615,N30616);
and and18437(N30628,N30629,N30630);
and and18446(N30642,N30643,N30644);
and and18455(N30656,N30657,N30658);
and and18464(N30670,N30671,N30672);
and and18473(N30684,N30685,N30686);
and and18482(N30698,N30699,N30700);
and and18491(N30712,N30713,N30714);
and and18500(N30726,N30727,N30728);
and and18509(N30740,N30741,N30742);
and and18518(N30754,N30755,N30756);
and and18527(N30768,N30769,N30770);
and and18536(N30782,N30783,N30784);
and and18545(N30796,N30797,N30798);
and and18554(N30810,N30811,N30812);
and and18563(N30824,N30825,N30826);
and and18572(N30838,N30839,N30840);
and and18581(N30852,N30853,N30854);
and and18590(N30866,N30867,N30868);
and and18599(N30880,N30881,N30882);
and and18608(N30894,N30895,N30896);
and and18617(N30908,N30909,N30910);
and and18626(N30922,N30923,N30924);
and and18635(N30936,N30937,N30938);
and and18644(N30950,N30951,N30952);
and and18653(N30964,N30965,N30966);
and and18662(N30977,N30978,N30979);
and and18671(N30990,N30991,N30992);
and and18680(N31003,N31004,N31005);
and and18689(N31016,N31017,N31018);
and and18698(N31029,N31030,N31031);
and and18707(N31042,N31043,N31044);
and and18716(N31055,N31056,N31057);
and and18725(N31068,N31069,N31070);
and and18734(N31081,N31082,N31083);
and and18743(N31094,N31095,N31096);
and and18752(N31107,N31108,N31109);
and and18761(N31120,N31121,N31122);
and and18770(N31133,N31134,N31135);
and and18779(N31146,N31147,N31148);
and and18788(N31159,N31160,N31161);
and and18797(N31172,N31173,N31174);
and and18806(N31185,N31186,N31187);
and and18815(N31198,N31199,N31200);
and and18824(N31211,N31212,N31213);
and and18833(N31224,N31225,N31226);
and and18842(N31237,N31238,N31239);
and and18851(N31249,N31250,N31251);
and and18860(N31261,N31262,N31263);
and and18869(N31273,N31274,N31275);
and and18878(N31285,N31286,N31287);
and and18887(N31297,N31298,N31299);
and and18896(N31309,N31310,N31311);
and and18905(N31321,N31322,N31323);
and and18914(N31333,N31334,N31335);
and and18923(N31345,N31346,N31347);
and and18932(N31357,N31358,N31359);
and and18941(N31367,N31368,N31369);
and and18950(N31377,N31378,N31379);
and and18959(N31387,N31388,N31389);
and and18968(N31397,N31398,N31399);
and and18977(N31407,N31408,N31409);
and and18985(N31423,N31424,N31425);
and and18993(N31439,N31440,N31441);
and and19001(N31455,N31456,N31457);
and and19009(N31470,N31471,N31472);
and and19017(N31485,N31486,N31487);
and and19025(N31500,N31501,N31502);
and and19033(N31514,N31515,N31516);
and and19041(N31528,N31529,N31530);
and and19049(N31542,N31543,N31544);
and and19057(N31556,N31557,N31558);
and and19065(N31570,N31571,N31572);
and and19073(N31584,N31585,N31586);
and and19081(N31597,N31598,N31599);
and and19089(N31610,N31611,N31612);
and and19097(N31623,N31624,N31625);
and and19105(N31635,N31636,N31637);
and and19113(N31647,N31648,N31649);
and and19121(N31659,N31660,N31661);
and and19129(N31671,N31672,N31673);
and and19137(N31683,N31684,N31685);
and and19145(N31694,N31695,N31696);
and and19153(N31705,N31706,N31707);
and and19161(N31716,N31717,N31718);
and and19169(N31726,N31727,N31728);
and and17738(N29435,N29437,N29438);
and and17739(N29436,N29439,N29440);
and and17748(N29453,N29455,N29456);
and and17749(N29454,N29457,N29458);
and and17758(N29471,N29473,N29474);
and and17759(N29472,N29475,N29476);
and and17768(N29488,N29490,N29491);
and and17769(N29489,N29492,N29493);
and and17778(N29505,N29507,N29508);
and and17779(N29506,N29509,N29510);
and and17788(N29521,N29523,N29524);
and and17789(N29522,N29525,N29526);
and and17798(N29537,N29539,N29540);
and and17799(N29538,N29541,N29542);
and and17808(N29551,N29553,N29554);
and and17809(N29552,N29555,N29556);
and and17817(N29569,N29571,N29572);
and and17818(N29570,N29573,N29574);
and and17826(N29587,N29589,N29590);
and and17827(N29588,N29591,N29592);
and and17835(N29605,N29607,N29608);
and and17836(N29606,N29609,N29610);
and and17844(N29622,N29624,N29625);
and and17845(N29623,N29626,N29627);
and and17853(N29639,N29641,N29642);
and and17854(N29640,N29643,N29644);
and and17862(N29656,N29658,N29659);
and and17863(N29657,N29660,N29661);
and and17871(N29673,N29675,N29676);
and and17872(N29674,N29677,N29678);
and and17880(N29690,N29692,N29693);
and and17881(N29691,N29694,N29695);
and and17889(N29707,N29709,N29710);
and and17890(N29708,N29711,N29712);
and and17898(N29723,N29725,N29726);
and and17899(N29724,N29727,N29728);
and and17907(N29739,N29741,N29742);
and and17908(N29740,N29743,N29744);
and and17916(N29755,N29757,N29758);
and and17917(N29756,N29759,N29760);
and and17925(N29771,N29773,N29774);
and and17926(N29772,N29775,N29776);
and and17934(N29787,N29789,N29790);
and and17935(N29788,N29791,N29792);
and and17943(N29803,N29805,N29806);
and and17944(N29804,N29807,N29808);
and and17952(N29819,N29821,N29822);
and and17953(N29820,N29823,N29824);
and and17961(N29835,N29837,N29838);
and and17962(N29836,N29839,N29840);
and and17970(N29851,N29853,N29854);
and and17971(N29852,N29855,N29856);
and and17979(N29867,N29869,N29870);
and and17980(N29868,N29871,N29872);
and and17988(N29883,N29885,N29886);
and and17989(N29884,N29887,N29888);
and and17997(N29899,N29901,N29902);
and and17998(N29900,N29903,N29904);
and and18006(N29915,N29917,N29918);
and and18007(N29916,N29919,N29920);
and and18015(N29931,N29933,N29934);
and and18016(N29932,N29935,N29936);
and and18024(N29947,N29949,N29950);
and and18025(N29948,N29951,N29952);
and and18033(N29963,N29965,N29966);
and and18034(N29964,N29967,N29968);
and and18042(N29979,N29981,N29982);
and and18043(N29980,N29983,N29984);
and and18051(N29995,N29997,N29998);
and and18052(N29996,N29999,N30000);
and and18060(N30010,N30012,N30013);
and and18061(N30011,N30014,N30015);
and and18069(N30025,N30027,N30028);
and and18070(N30026,N30029,N30030);
and and18078(N30040,N30042,N30043);
and and18079(N30041,N30044,N30045);
and and18087(N30055,N30057,N30058);
and and18088(N30056,N30059,N30060);
and and18096(N30070,N30072,N30073);
and and18097(N30071,N30074,N30075);
and and18105(N30085,N30087,N30088);
and and18106(N30086,N30089,N30090);
and and18114(N30100,N30102,N30103);
and and18115(N30101,N30104,N30105);
and and18123(N30115,N30117,N30118);
and and18124(N30116,N30119,N30120);
and and18132(N30130,N30132,N30133);
and and18133(N30131,N30134,N30135);
and and18141(N30145,N30147,N30148);
and and18142(N30146,N30149,N30150);
and and18150(N30160,N30162,N30163);
and and18151(N30161,N30164,N30165);
and and18159(N30175,N30177,N30178);
and and18160(N30176,N30179,N30180);
and and18168(N30190,N30192,N30193);
and and18169(N30191,N30194,N30195);
and and18177(N30205,N30207,N30208);
and and18178(N30206,N30209,N30210);
and and18186(N30220,N30222,N30223);
and and18187(N30221,N30224,N30225);
and and18195(N30235,N30237,N30238);
and and18196(N30236,N30239,N30240);
and and18204(N30250,N30252,N30253);
and and18205(N30251,N30254,N30255);
and and18213(N30265,N30267,N30268);
and and18214(N30266,N30269,N30270);
and and18222(N30280,N30282,N30283);
and and18223(N30281,N30284,N30285);
and and18231(N30295,N30297,N30298);
and and18232(N30296,N30299,N30300);
and and18240(N30310,N30312,N30313);
and and18241(N30311,N30314,N30315);
and and18249(N30325,N30327,N30328);
and and18250(N30326,N30329,N30330);
and and18258(N30340,N30342,N30343);
and and18259(N30341,N30344,N30345);
and and18267(N30355,N30357,N30358);
and and18268(N30356,N30359,N30360);
and and18276(N30370,N30372,N30373);
and and18277(N30371,N30374,N30375);
and and18285(N30385,N30387,N30388);
and and18286(N30386,N30389,N30390);
and and18294(N30400,N30402,N30403);
and and18295(N30401,N30404,N30405);
and and18303(N30415,N30417,N30418);
and and18304(N30416,N30419,N30420);
and and18312(N30430,N30432,N30433);
and and18313(N30431,N30434,N30435);
and and18321(N30445,N30447,N30448);
and and18322(N30446,N30449,N30450);
and and18330(N30460,N30462,N30463);
and and18331(N30461,N30464,N30465);
and and18339(N30475,N30477,N30478);
and and18340(N30476,N30479,N30480);
and and18348(N30489,N30491,N30492);
and and18349(N30490,N30493,N30494);
and and18357(N30503,N30505,N30506);
and and18358(N30504,N30507,N30508);
and and18366(N30517,N30519,N30520);
and and18367(N30518,N30521,N30522);
and and18375(N30531,N30533,N30534);
and and18376(N30532,N30535,N30536);
and and18384(N30545,N30547,N30548);
and and18385(N30546,N30549,N30550);
and and18393(N30559,N30561,N30562);
and and18394(N30560,N30563,N30564);
and and18402(N30573,N30575,N30576);
and and18403(N30574,N30577,N30578);
and and18411(N30587,N30589,N30590);
and and18412(N30588,N30591,N30592);
and and18420(N30601,N30603,N30604);
and and18421(N30602,N30605,N30606);
and and18429(N30615,N30617,N30618);
and and18430(N30616,N30619,N30620);
and and18438(N30629,N30631,N30632);
and and18439(N30630,N30633,N30634);
and and18447(N30643,N30645,N30646);
and and18448(N30644,N30647,N30648);
and and18456(N30657,N30659,N30660);
and and18457(N30658,N30661,N30662);
and and18465(N30671,N30673,N30674);
and and18466(N30672,N30675,N30676);
and and18474(N30685,N30687,N30688);
and and18475(N30686,N30689,N30690);
and and18483(N30699,N30701,N30702);
and and18484(N30700,N30703,N30704);
and and18492(N30713,N30715,N30716);
and and18493(N30714,N30717,N30718);
and and18501(N30727,N30729,N30730);
and and18502(N30728,N30731,N30732);
and and18510(N30741,N30743,N30744);
and and18511(N30742,N30745,N30746);
and and18519(N30755,N30757,N30758);
and and18520(N30756,N30759,N30760);
and and18528(N30769,N30771,N30772);
and and18529(N30770,N30773,N30774);
and and18537(N30783,N30785,N30786);
and and18538(N30784,N30787,N30788);
and and18546(N30797,N30799,N30800);
and and18547(N30798,N30801,N30802);
and and18555(N30811,N30813,N30814);
and and18556(N30812,N30815,N30816);
and and18564(N30825,N30827,N30828);
and and18565(N30826,N30829,N30830);
and and18573(N30839,N30841,N30842);
and and18574(N30840,N30843,N30844);
and and18582(N30853,N30855,N30856);
and and18583(N30854,N30857,N30858);
and and18591(N30867,N30869,N30870);
and and18592(N30868,N30871,N30872);
and and18600(N30881,N30883,N30884);
and and18601(N30882,N30885,N30886);
and and18609(N30895,N30897,N30898);
and and18610(N30896,N30899,N30900);
and and18618(N30909,N30911,N30912);
and and18619(N30910,N30913,N30914);
and and18627(N30923,N30925,N30926);
and and18628(N30924,N30927,N30928);
and and18636(N30937,N30939,N30940);
and and18637(N30938,N30941,N30942);
and and18645(N30951,N30953,N30954);
and and18646(N30952,N30955,N30956);
and and18654(N30965,N30967,N30968);
and and18655(N30966,N30969,N30970);
and and18663(N30978,N30980,N30981);
and and18664(N30979,N30982,N30983);
and and18672(N30991,N30993,N30994);
and and18673(N30992,N30995,N30996);
and and18681(N31004,N31006,N31007);
and and18682(N31005,N31008,N31009);
and and18690(N31017,N31019,N31020);
and and18691(N31018,N31021,N31022);
and and18699(N31030,N31032,N31033);
and and18700(N31031,N31034,N31035);
and and18708(N31043,N31045,N31046);
and and18709(N31044,N31047,N31048);
and and18717(N31056,N31058,N31059);
and and18718(N31057,N31060,N31061);
and and18726(N31069,N31071,N31072);
and and18727(N31070,N31073,N31074);
and and18735(N31082,N31084,N31085);
and and18736(N31083,N31086,N31087);
and and18744(N31095,N31097,N31098);
and and18745(N31096,N31099,N31100);
and and18753(N31108,N31110,N31111);
and and18754(N31109,N31112,N31113);
and and18762(N31121,N31123,N31124);
and and18763(N31122,N31125,N31126);
and and18771(N31134,N31136,N31137);
and and18772(N31135,N31138,N31139);
and and18780(N31147,N31149,N31150);
and and18781(N31148,N31151,N31152);
and and18789(N31160,N31162,N31163);
and and18790(N31161,N31164,N31165);
and and18798(N31173,N31175,N31176);
and and18799(N31174,N31177,N31178);
and and18807(N31186,N31188,N31189);
and and18808(N31187,N31190,N31191);
and and18816(N31199,N31201,N31202);
and and18817(N31200,N31203,N31204);
and and18825(N31212,N31214,N31215);
and and18826(N31213,N31216,N31217);
and and18834(N31225,N31227,N31228);
and and18835(N31226,N31229,N31230);
and and18843(N31238,N31240,N31241);
and and18844(N31239,N31242,N31243);
and and18852(N31250,N31252,N31253);
and and18853(N31251,N31254,N31255);
and and18861(N31262,N31264,N31265);
and and18862(N31263,N31266,N31267);
and and18870(N31274,N31276,N31277);
and and18871(N31275,N31278,N31279);
and and18879(N31286,N31288,N31289);
and and18880(N31287,N31290,N31291);
and and18888(N31298,N31300,N31301);
and and18889(N31299,N31302,N31303);
and and18897(N31310,N31312,N31313);
and and18898(N31311,N31314,N31315);
and and18906(N31322,N31324,N31325);
and and18907(N31323,N31326,N31327);
and and18915(N31334,N31336,N31337);
and and18916(N31335,N31338,N31339);
and and18924(N31346,N31348,N31349);
and and18925(N31347,N31350,N31351);
and and18933(N31358,N31360,N31361);
and and18934(N31359,N31362,N31363);
and and18942(N31368,N31370,N31371);
and and18943(N31369,N31372,N31373);
and and18951(N31378,N31380,N31381);
and and18952(N31379,N31382,N31383);
and and18960(N31388,N31390,N31391);
and and18961(N31389,N31392,N31393);
and and18969(N31398,N31400,N31401);
and and18970(N31399,N31402,N31403);
and and18978(N31408,N31410,N31411);
and and18979(N31409,N31412,N31413);
and and18986(N31424,N31426,N31427);
and and18987(N31425,N31428,N31429);
and and18994(N31440,N31442,N31443);
and and18995(N31441,N31444,N31445);
and and19002(N31456,N31458,N31459);
and and19003(N31457,N31460,N31461);
and and19010(N31471,N31473,N31474);
and and19011(N31472,N31475,N31476);
and and19018(N31486,N31488,N31489);
and and19019(N31487,N31490,N31491);
and and19026(N31501,N31503,N31504);
and and19027(N31502,N31505,N31506);
and and19034(N31515,N31517,N31518);
and and19035(N31516,N31519,N31520);
and and19042(N31529,N31531,N31532);
and and19043(N31530,N31533,N31534);
and and19050(N31543,N31545,N31546);
and and19051(N31544,N31547,N31548);
and and19058(N31557,N31559,N31560);
and and19059(N31558,N31561,N31562);
and and19066(N31571,N31573,N31574);
and and19067(N31572,N31575,N31576);
and and19074(N31585,N31587,N31588);
and and19075(N31586,N31589,N31590);
and and19082(N31598,N31600,N31601);
and and19083(N31599,N31602,N31603);
and and19090(N31611,N31613,N31614);
and and19091(N31612,N31615,N31616);
and and19098(N31624,N31626,N31627);
and and19099(N31625,N31628,N31629);
and and19106(N31636,N31638,N31639);
and and19107(N31637,N31640,N31641);
and and19114(N31648,N31650,N31651);
and and19115(N31649,N31652,N31653);
and and19122(N31660,N31662,N31663);
and and19123(N31661,N31664,N31665);
and and19130(N31672,N31674,N31675);
and and19131(N31673,N31676,N31677);
and and19138(N31684,N31686,N31687);
and and19139(N31685,N31688,N31689);
and and19146(N31695,N31697,N31698);
and and19147(N31696,N31699,N31700);
and and19154(N31706,N31708,N31709);
and and19155(N31707,N31710,N31711);
and and19162(N31717,N31719,N31720);
and and19163(N31718,N31721,N31722);
and and19170(N31727,N31729,N31730);
and and19171(N31728,N31731,N31732);
and and17740(N29437,N29441,N29442);
and and17741(N29438,N29443,N29444);
and and17742(N29439,in1,N29445);
and and17743(N29440,N29446,N29447);
and and17750(N29455,N29459,N29460);
and and17751(N29456,N29461,N29462);
and and17752(N29457,in1,N29463);
and and17753(N29458,R0,N29464);
and and17760(N29473,N29477,N29478);
and and17761(N29474,N29479,N29480);
and and17762(N29475,N29481,N29482);
and and17763(N29476,R0,R1);
and and17770(N29490,N29494,N29495);
and and17771(N29491,N29496,N29497);
and and17772(N29492,N29498,in2);
and and17773(N29493,N29499,R1);
and and17780(N29507,N29511,N29512);
and and17781(N29508,N29513,N29514);
and and17782(N29509,in1,N29515);
and and17783(N29510,N29516,N29517);
and and17790(N29523,N29527,N29528);
and and17791(N29524,N29529,N29530);
and and17792(N29525,in1,N29531);
and and17793(N29526,N29532,N29533);
and and17800(N29539,N29543,N29544);
and and17801(N29540,N29545,N29546);
and and17802(N29541,N29547,in2);
and and17803(N29542,R0,N29548);
and and17810(N29553,N29557,N29558);
and and17811(N29554,N29559,N29560);
and and17812(N29555,N29561,N29562);
and and17813(N29556,N29563,N29564);
and and17819(N29571,N29575,N29576);
and and17820(N29572,N29577,N29578);
and and17821(N29573,N29579,R0);
and and17822(N29574,N29580,N29581);
and and17828(N29589,N29593,N29594);
and and17829(N29590,N29595,N29596);
and and17830(N29591,N29597,R0);
and and17831(N29592,N29598,N29599);
and and17837(N29607,N29611,N29612);
and and17838(N29608,N29613,N29614);
and and17839(N29609,in2,N29615);
and and17840(N29610,R1,N29616);
and and17846(N29624,N29628,N29629);
and and17847(N29625,N29630,in2);
and and17848(N29626,N29631,N29632);
and and17849(N29627,N29633,N29634);
and and17855(N29641,N29645,N29646);
and and17856(N29642,N29647,N29648);
and and17857(N29643,N29649,N29650);
and and17858(N29644,N29651,R2);
and and17864(N29658,N29662,N29663);
and and17865(N29659,N29664,in1);
and and17866(N29660,in2,N29665);
and and17867(N29661,N29666,N29667);
and and17873(N29675,N29679,N29680);
and and17874(N29676,N29681,in2);
and and17875(N29677,N29682,N29683);
and and17876(N29678,N29684,N29685);
and and17882(N29692,N29696,N29697);
and and17883(N29693,N29698,in1);
and and17884(N29694,N29699,N29700);
and and17885(N29695,N29701,N29702);
and and17891(N29709,N29713,N29714);
and and17892(N29710,N29715,N29716);
and and17893(N29711,in2,N29717);
and and17894(N29712,N29718,N29719);
and and17900(N29725,N29729,N29730);
and and17901(N29726,N29731,N29732);
and and17902(N29727,R0,N29733);
and and17903(N29728,N29734,R3);
and and17909(N29741,N29745,N29746);
and and17910(N29742,N29747,N29748);
and and17911(N29743,in2,N29749);
and and17912(N29744,R2,N29750);
and and17918(N29757,N29761,N29762);
and and17919(N29758,N29763,N29764);
and and17920(N29759,N29765,N29766);
and and17921(N29760,R2,N29767);
and and17927(N29773,N29777,N29778);
and and17928(N29774,N29779,in1);
and and17929(N29775,N29780,N29781);
and and17930(N29776,R2,N29782);
and and17936(N29789,N29793,N29794);
and and17937(N29790,N29795,N29796);
and and17938(N29791,in2,R0);
and and17939(N29792,N29797,R3);
and and17945(N29805,N29809,N29810);
and and17946(N29806,N29811,N29812);
and and17947(N29807,N29813,N29814);
and and17948(N29808,R2,N29815);
and and17954(N29821,N29825,N29826);
and and17955(N29822,N29827,N29828);
and and17956(N29823,N29829,N29830);
and and17957(N29824,N29831,R3);
and and17963(N29837,N29841,N29842);
and and17964(N29838,N29843,N29844);
and and17965(N29839,in2,N29845);
and and17966(N29840,N29846,R3);
and and17972(N29853,N29857,N29858);
and and17973(N29854,N29859,in1);
and and17974(N29855,N29860,R1);
and and17975(N29856,N29861,N29862);
and and17981(N29869,N29873,N29874);
and and17982(N29870,N29875,N29876);
and and17983(N29871,N29877,N29878);
and and17984(N29872,N29879,R3);
and and17990(N29885,N29889,N29890);
and and17991(N29886,N29891,N29892);
and and17992(N29887,N29893,N29894);
and and17993(N29888,R1,N29895);
and and17999(N29901,N29905,N29906);
and and18000(N29902,N29907,in1);
and and18001(N29903,N29908,R0);
and and18002(N29904,N29909,N29910);
and and18008(N29917,N29921,N29922);
and and18009(N29918,N29923,N29924);
and and18010(N29919,in2,N29925);
and and18011(N29920,R1,N29926);
and and18017(N29933,N29937,N29938);
and and18018(N29934,N29939,N29940);
and and18019(N29935,N29941,N29942);
and and18020(N29936,R2,N29943);
and and18026(N29949,N29953,N29954);
and and18027(N29950,N29955,N29956);
and and18028(N29951,N29957,N29958);
and and18029(N29952,R1,R2);
and and18035(N29965,N29969,N29970);
and and18036(N29966,N29971,in1);
and and18037(N29967,in2,N29972);
and and18038(N29968,N29973,N29974);
and and18044(N29981,N29985,N29986);
and and18045(N29982,N29987,in1);
and and18046(N29983,in2,N29988);
and and18047(N29984,N29989,N29990);
and and18053(N29997,N30001,N30002);
and and18054(N29998,N30003,N30004);
and and18055(N29999,N30005,R1);
and and18056(N30000,N30006,R3);
and and18062(N30012,N30016,N30017);
and and18063(N30013,N30018,in1);
and and18064(N30014,N30019,R0);
and and18065(N30015,R1,N30020);
and and18071(N30027,N30031,N30032);
and and18072(N30028,N30033,N30034);
and and18073(N30029,in2,R0);
and and18074(N30030,R1,N30035);
and and18080(N30042,N30046,N30047);
and and18081(N30043,N30048,in1);
and and18082(N30044,in2,N30049);
and and18083(N30045,R2,N30050);
and and18089(N30057,N30061,N30062);
and and18090(N30058,N30063,in1);
and and18091(N30059,in2,N30064);
and and18092(N30060,N30065,R3);
and and18098(N30072,N30076,N30077);
and and18099(N30073,N30078,N30079);
and and18100(N30074,R0,N30080);
and and18101(N30075,R2,R3);
and and18107(N30087,N30091,N30092);
and and18108(N30088,N30093,N30094);
and and18109(N30089,N30095,R0);
and and18110(N30090,N30096,N30097);
and and18116(N30102,N30106,N30107);
and and18117(N30103,N30108,in1);
and and18118(N30104,N30109,N30110);
and and18119(N30105,R1,N30111);
and and18125(N30117,N30121,N30122);
and and18126(N30118,N30123,in1);
and and18127(N30119,in2,N30124);
and and18128(N30120,N30125,R3);
and and18134(N30132,N30136,N30137);
and and18135(N30133,N30138,in1);
and and18136(N30134,in2,R1);
and and18137(N30135,R2,N30139);
and and18143(N30147,N30151,N30152);
and and18144(N30148,N30153,in1);
and and18145(N30149,in2,N30154);
and and18146(N30150,N30155,R2);
and and18152(N30162,N30166,N30167);
and and18153(N30163,N30168,N30169);
and and18154(N30164,in2,R0);
and and18155(N30165,R1,N30170);
and and18161(N30177,N30181,N30182);
and and18162(N30178,N30183,in1);
and and18163(N30179,N30184,N30185);
and and18164(N30180,R1,R2);
and and18170(N30192,N30196,N30197);
and and18171(N30193,N30198,N30199);
and and18172(N30194,R0,R1);
and and18173(N30195,R2,N30200);
and and18179(N30207,N30211,N30212);
and and18180(N30208,N30213,in1);
and and18181(N30209,in2,R0);
and and18182(N30210,N30214,N30215);
and and18188(N30222,N30226,N30227);
and and18189(N30223,N30228,in1);
and and18190(N30224,N30229,N30230);
and and18191(N30225,R1,N30231);
and and18197(N30237,N30241,N30242);
and and18198(N30238,N30243,in1);
and and18199(N30239,in2,N30244);
and and18200(N30240,R1,N30245);
and and18206(N30252,N30256,N30257);
and and18207(N30253,N30258,in1);
and and18208(N30254,in2,N30259);
and and18209(N30255,R1,N30260);
and and18215(N30267,N30271,N30272);
and and18216(N30268,N30273,in2);
and and18217(N30269,R0,N30274);
and and18218(N30270,N30275,R3);
and and18224(N30282,N30286,N30287);
and and18225(N30283,N30288,N30289);
and and18226(N30284,in2,N30290);
and and18227(N30285,R1,N30291);
and and18233(N30297,N30301,N30302);
and and18234(N30298,N30303,in1);
and and18235(N30299,N30304,N30305);
and and18236(N30300,R1,N30306);
and and18242(N30312,N30316,N30317);
and and18243(N30313,N30318,N30319);
and and18244(N30314,N30320,R0);
and and18245(N30315,R1,N30321);
and and18251(N30327,N30331,N30332);
and and18252(N30328,N30333,N30334);
and and18253(N30329,in2,R1);
and and18254(N30330,R2,N30335);
and and18260(N30342,N30346,N30347);
and and18261(N30343,N30348,in1);
and and18262(N30344,in2,N30349);
and and18263(N30345,R1,N30350);
and and18269(N30357,N30361,N30362);
and and18270(N30358,N30363,N30364);
and and18271(N30359,N30365,R0);
and and18272(N30360,R1,N30366);
and and18278(N30372,N30376,N30377);
and and18279(N30373,N30378,in2);
and and18280(N30374,R0,R1);
and and18281(N30375,N30379,N30380);
and and18287(N30387,N30391,N30392);
and and18288(N30388,N30393,N30394);
and and18289(N30389,N30395,R1);
and and18290(N30390,R2,N30396);
and and18296(N30402,N30406,N30407);
and and18297(N30403,N30408,N30409);
and and18298(N30404,in2,R1);
and and18299(N30405,R2,N30410);
and and18305(N30417,N30421,N30422);
and and18306(N30418,N30423,in1);
and and18307(N30419,R0,N30424);
and and18308(N30420,R2,N30425);
and and18314(N30432,N30436,N30437);
and and18315(N30433,N30438,in1);
and and18316(N30434,N30439,R0);
and and18317(N30435,R1,N30440);
and and18323(N30447,N30451,N30452);
and and18324(N30448,N30453,in1);
and and18325(N30449,N30454,R0);
and and18326(N30450,R1,N30455);
and and18332(N30462,N30466,N30467);
and and18333(N30463,N30468,N30469);
and and18334(N30464,in2,N30470);
and and18335(N30465,N30471,R2);
and and18341(N30477,N30481,N30482);
and and18342(N30478,N30483,in1);
and and18343(N30479,R0,R1);
and and18344(N30480,N30484,R3);
and and18350(N30491,N30495,N30496);
and and18351(N30492,N30497,in1);
and and18352(N30493,N30498,R1);
and and18353(N30494,R2,N30499);
and and18359(N30505,N30509,N30510);
and and18360(N30506,N30511,N30512);
and and18361(N30507,in2,R0);
and and18362(N30508,R2,N30513);
and and18368(N30519,N30523,N30524);
and and18369(N30520,N30525,in1);
and and18370(N30521,in2,R0);
and and18371(N30522,N30526,N30527);
and and18377(N30533,N30537,N30538);
and and18378(N30534,N30539,in1);
and and18379(N30535,in2,N30540);
and and18380(N30536,N30541,R3);
and and18386(N30547,N30551,N30552);
and and18387(N30548,N30553,N30554);
and and18388(N30549,N30555,N30556);
and and18389(N30550,R2,R3);
and and18395(N30561,N30565,N30566);
and and18396(N30562,N30567,N30568);
and and18397(N30563,R0,N30569);
and and18398(N30564,N30570,R3);
and and18404(N30575,N30579,N30580);
and and18405(N30576,N30581,in2);
and and18406(N30577,N30582,N30583);
and and18407(N30578,R2,R3);
and and18413(N30589,N30593,N30594);
and and18414(N30590,N30595,N30596);
and and18415(N30591,N30597,R1);
and and18416(N30592,R2,R3);
and and18422(N30603,N30607,N30608);
and and18423(N30604,N30609,in2);
and and18424(N30605,R0,N30610);
and and18425(N30606,R2,N30611);
and and18431(N30617,N30621,N30622);
and and18432(N30618,N30623,N30624);
and and18433(N30619,in2,R0);
and and18434(N30620,R2,N30625);
and and18440(N30631,N30635,N30636);
and and18441(N30632,N30637,in1);
and and18442(N30633,R0,N30638);
and and18443(N30634,N30639,R3);
and and18449(N30645,N30649,N30650);
and and18450(N30646,N30651,N30652);
and and18451(N30647,in2,R1);
and and18452(N30648,N30653,R3);
and and18458(N30659,N30663,N30664);
and and18459(N30660,N30665,in1);
and and18460(N30661,N30666,N30667);
and and18461(N30662,R2,N30668);
and and18467(N30673,N30677,N30678);
and and18468(N30674,N30679,in1);
and and18469(N30675,in2,R0);
and and18470(N30676,N30680,N30681);
and and18476(N30687,N30691,N30692);
and and18477(N30688,N30693,N30694);
and and18478(N30689,R0,R1);
and and18479(N30690,R2,R3);
and and18485(N30701,N30705,N30706);
and and18486(N30702,N30707,in1);
and and18487(N30703,N30708,R0);
and and18488(N30704,N30709,R2);
and and18494(N30715,N30719,N30720);
and and18495(N30716,N30721,N30722);
and and18496(N30717,in2,N30723);
and and18497(N30718,R1,N30724);
and and18503(N30729,N30733,N30734);
and and18504(N30730,N30735,in1);
and and18505(N30731,in2,N30736);
and and18506(N30732,N30737,R3);
and and18512(N30743,N30747,N30748);
and and18513(N30744,N30749,N30750);
and and18514(N30745,in2,N30751);
and and18515(N30746,R2,N30752);
and and18521(N30757,N30761,N30762);
and and18522(N30758,N30763,in1);
and and18523(N30759,N30764,N30765);
and and18524(N30760,R2,N30766);
and and18530(N30771,N30775,N30776);
and and18531(N30772,N30777,in1);
and and18532(N30773,in2,N30778);
and and18533(N30774,R1,N30779);
and and18539(N30785,N30789,N30790);
and and18540(N30786,N30791,N30792);
and and18541(N30787,N30793,N30794);
and and18542(N30788,R1,R2);
and and18548(N30799,N30803,N30804);
and and18549(N30800,N30805,in1);
and and18550(N30801,N30806,R0);
and and18551(N30802,N30807,R2);
and and18557(N30813,N30817,N30818);
and and18558(N30814,N30819,N30820);
and and18559(N30815,in2,R0);
and and18560(N30816,N30821,R2);
and and18566(N30827,N30831,N30832);
and and18567(N30828,N30833,in1);
and and18568(N30829,N30834,R0);
and and18569(N30830,R1,R2);
and and18575(N30841,N30845,N30846);
and and18576(N30842,N30847,in1);
and and18577(N30843,in2,N30848);
and and18578(N30844,N30849,R2);
and and18584(N30855,N30859,N30860);
and and18585(N30856,N30861,N30862);
and and18586(N30857,N30863,R0);
and and18587(N30858,N30864,R2);
and and18593(N30869,N30873,N30874);
and and18594(N30870,N30875,in1);
and and18595(N30871,N30876,R0);
and and18596(N30872,N30877,N30878);
and and18602(N30883,N30887,N30888);
and and18603(N30884,N30889,N30890);
and and18604(N30885,in2,R0);
and and18605(N30886,N30891,N30892);
and and18611(N30897,N30901,N30902);
and and18612(N30898,N30903,N30904);
and and18613(N30899,in2,N30905);
and and18614(N30900,R2,R3);
and and18620(N30911,N30915,N30916);
and and18621(N30912,N30917,in1);
and and18622(N30913,N30918,N30919);
and and18623(N30914,R2,R3);
and and18629(N30925,N30929,N30930);
and and18630(N30926,N30931,in1);
and and18631(N30927,in2,N30932);
and and18632(N30928,R1,N30933);
and and18638(N30939,N30943,N30944);
and and18639(N30940,N30945,in1);
and and18640(N30941,N30946,R0);
and and18641(N30942,R1,N30947);
and and18647(N30953,N30957,N30958);
and and18648(N30954,N30959,in2);
and and18649(N30955,R0,N30960);
and and18650(N30956,R2,N30961);
and and18656(N30967,N30971,N30972);
and and18657(N30968,N30973,in1);
and and18658(N30969,N30974,R1);
and and18659(N30970,N30975,R3);
and and18665(N30980,N30984,N30985);
and and18666(N30981,N30986,in1);
and and18667(N30982,in2,R0);
and and18668(N30983,R1,R3);
and and18674(N30993,N30997,N30998);
and and18675(N30994,N30999,in2);
and and18676(N30995,R0,N31000);
and and18677(N30996,N31001,R3);
and and18683(N31006,N31010,N31011);
and and18684(N31007,N31012,in1);
and and18685(N31008,in2,N31013);
and and18686(N31009,R1,R2);
and and18692(N31019,N31023,N31024);
and and18693(N31020,N31025,in2);
and and18694(N31021,R0,R1);
and and18695(N31022,R2,R3);
and and18701(N31032,N31036,N31037);
and and18702(N31033,N31038,in1);
and and18703(N31034,in2,R0);
and and18704(N31035,R1,N31039);
and and18710(N31045,N31049,N31050);
and and18711(N31046,N31051,in1);
and and18712(N31047,in2,N31052);
and and18713(N31048,R1,R2);
and and18719(N31058,N31062,N31063);
and and18720(N31059,N31064,in2);
and and18721(N31060,N31065,R1);
and and18722(N31061,N31066,R3);
and and18728(N31071,N31075,N31076);
and and18729(N31072,N31077,in1);
and and18730(N31073,N31078,R1);
and and18731(N31074,R2,N31079);
and and18737(N31084,N31088,N31089);
and and18738(N31085,N31090,in1);
and and18739(N31086,in2,N31091);
and and18740(N31087,N31092,R3);
and and18746(N31097,N31101,N31102);
and and18747(N31098,N31103,in1);
and and18748(N31099,in2,N31104);
and and18749(N31100,R1,N31105);
and and18755(N31110,N31114,N31115);
and and18756(N31111,N31116,in1);
and and18757(N31112,in2,R0);
and and18758(N31113,R1,N31117);
and and18764(N31123,N31127,N31128);
and and18765(N31124,N31129,N31130);
and and18766(N31125,R0,N31131);
and and18767(N31126,R2,R3);
and and18773(N31136,N31140,N31141);
and and18774(N31137,N31142,in1);
and and18775(N31138,in2,N31143);
and and18776(N31139,R1,R2);
and and18782(N31149,N31153,N31154);
and and18783(N31150,N31155,N31156);
and and18784(N31151,in2,R0);
and and18785(N31152,R1,R2);
and and18791(N31162,N31166,N31167);
and and18792(N31163,N31168,N31169);
and and18793(N31164,in2,R0);
and and18794(N31165,R1,N31170);
and and18800(N31175,N31179,N31180);
and and18801(N31176,N31181,N31182);
and and18802(N31177,R0,R1);
and and18803(N31178,R2,N31183);
and and18809(N31188,N31192,N31193);
and and18810(N31189,N31194,in1);
and and18811(N31190,R0,N31195);
and and18812(N31191,R2,R3);
and and18818(N31201,N31205,N31206);
and and18819(N31202,N31207,in1);
and and18820(N31203,in2,N31208);
and and18821(N31204,N31209,R2);
and and18827(N31214,N31218,N31219);
and and18828(N31215,N31220,in1);
and and18829(N31216,in2,R0);
and and18830(N31217,N31221,R2);
and and18836(N31227,N31231,N31232);
and and18837(N31228,N31233,N31234);
and and18838(N31229,in2,R0);
and and18839(N31230,R1,N31235);
and and18845(N31240,N31244,N31245);
and and18846(N31241,N31246,N31247);
and and18847(N31242,N31248,R0);
and and18848(N31243,R1,R3);
and and18854(N31252,N31256,N31257);
and and18855(N31253,N31258,in1);
and and18856(N31254,N31259,R0);
and and18857(N31255,R1,R2);
and and18863(N31264,N31268,N31269);
and and18864(N31265,N31270,in1);
and and18865(N31266,in2,R1);
and and18866(N31267,R2,R3);
and and18872(N31276,N31280,N31281);
and and18873(N31277,N31282,in1);
and and18874(N31278,in2,R0);
and and18875(N31279,N31283,R3);
and and18881(N31288,N31292,N31293);
and and18882(N31289,N31294,in1);
and and18883(N31290,in2,R0);
and and18884(N31291,R1,R2);
and and18890(N31300,N31304,N31305);
and and18891(N31301,N31306,N31307);
and and18892(N31302,N31308,R0);
and and18893(N31303,R1,R2);
and and18899(N31312,N31316,N31317);
and and18900(N31313,N31318,in1);
and and18901(N31314,in2,N31319);
and and18902(N31315,R1,R2);
and and18908(N31324,N31328,N31329);
and and18909(N31325,N31330,N31331);
and and18910(N31326,in2,R0);
and and18911(N31327,R1,R3);
and and18917(N31336,N31340,N31341);
and and18918(N31337,N31342,in1);
and and18919(N31338,N31343,R0);
and and18920(N31339,R1,R3);
and and18926(N31348,N31352,N31353);
and and18927(N31349,N31354,in1);
and and18928(N31350,R0,R1);
and and18929(N31351,R2,N31355);
and and18935(N31360,N31364,N31365);
and and18936(N31361,N31366,in1);
and and18937(N31362,in2,R0);
and and18938(N31363,R1,R3);
and and18944(N31370,N31374,N31375);
and and18945(N31371,N31376,in1);
and and18946(N31372,in2,R0);
and and18947(N31373,R2,R3);
and and18953(N31380,N31384,N31385);
and and18954(N31381,N31386,in1);
and and18955(N31382,in2,R0);
and and18956(N31383,R1,R2);
and and18962(N31390,N31394,N31395);
and and18963(N31391,N31396,in1);
and and18964(N31392,in2,R0);
and and18965(N31393,R1,R2);
and and18971(N31400,N31404,N31405);
and and18972(N31401,N31406,in1);
and and18973(N31402,in2,R1);
and and18974(N31403,R2,R3);
and and18980(N31410,N31414,N31415);
and and18981(N31411,in1,N31416);
and and18982(N31412,N31417,N31418);
and and18983(N31413,N31419,N31420);
and and18988(N31426,N31430,N31431);
and and18989(N31427,N31432,N31433);
and and18990(N31428,N31434,N31435);
and and18991(N31429,N31436,N31437);
and and18996(N31442,N31446,N31447);
and and18997(N31443,N31448,N31449);
and and18998(N31444,N31450,R2);
and and18999(N31445,N31451,N31452);
and and19004(N31458,N31462,N31463);
and and19005(N31459,in1,N31464);
and and19006(N31460,N31465,R3);
and and19007(N31461,N31466,N31467);
and and19012(N31473,N31477,N31478);
and and19013(N31474,N31479,N31480);
and and19014(N31475,N31481,R1);
and and19015(N31476,N31482,R4);
and and19020(N31488,N31492,N31493);
and and19021(N31489,N31494,N31495);
and and19022(N31490,R1,N31496);
and and19023(N31491,R4,N31497);
and and19028(N31503,N31507,N31508);
and and19029(N31504,N31509,R0);
and and19030(N31505,R1,N31510);
and and19031(N31506,R3,N31511);
and and19036(N31517,N31521,N31522);
and and19037(N31518,N31523,N31524);
and and19038(N31519,R0,N31525);
and and19039(N31520,R2,N31526);
and and19044(N31531,N31535,N31536);
and and19045(N31532,N31537,R0);
and and19046(N31533,R1,R2);
and and19047(N31534,N31538,N31539);
and and19052(N31545,N31549,N31550);
and and19053(N31546,in1,N31551);
and and19054(N31547,N31552,R1);
and and19055(N31548,N31553,N31554);
and and19060(N31559,N31563,N31564);
and and19061(N31560,N31565,N31566);
and and19062(N31561,N31567,R3);
and and19063(N31562,N31568,R5);
and and19068(N31573,N31577,N31578);
and and19069(N31574,N31579,in2);
and and19070(N31575,R0,N31580);
and and19071(N31576,N31581,R4);
and and19076(N31587,N31591,N31592);
and and19077(N31588,N31593,in2);
and and19078(N31589,N31594,R2);
and and19079(N31590,R3,N31595);
and and19084(N31600,N31604,N31605);
and and19085(N31601,N31606,in2);
and and19086(N31602,N31607,R3);
and and19087(N31603,N31608,N31609);
and and19092(N31613,N31617,N31618);
and and19093(N31614,N31619,N31620);
and and19094(N31615,N31621,R1);
and and19095(N31616,R3,R5);
and and19100(N31626,N31630,N31631);
and and19101(N31627,N31632,N31633);
and and19102(N31628,R1,R2);
and and19103(N31629,R3,N31634);
and and19108(N31638,N31642,N31643);
and and19109(N31639,in1,N31644);
and and19110(N31640,R2,R3);
and and19111(N31641,N31645,R5);
and and19116(N31650,N31654,N31655);
and and19117(N31651,N31656,R0);
and and19118(N31652,R1,R2);
and and19119(N31653,R3,N31657);
and and19124(N31662,N31666,N31667);
and and19125(N31663,N31668,in2);
and and19126(N31664,R0,R1);
and and19127(N31665,N31669,R4);
and and19132(N31674,N31678,N31679);
and and19133(N31675,N31680,N31681);
and and19134(N31676,R1,R2);
and and19135(N31677,R3,R5);
and and19140(N31686,N31690,N31691);
and and19141(N31687,N31692,N31693);
and and19142(N31688,R2,R3);
and and19143(N31689,R4,R5);
and and19148(N31697,N31701,N31702);
and and19149(N31698,in1,in2);
and and19150(N31699,R0,R3);
and and19151(N31700,R4,R5);
and and19156(N31708,N31712,N31713);
and and19157(N31709,in1,R0);
and and19158(N31710,R1,R2);
and and19159(N31711,R4,R5);
and and19164(N31719,N31723,N31724);
and and19165(N31720,R0,R1);
and and19166(N31721,R2,R3);
and and19167(N31722,R4,R5);
and and19172(N31729,N31733,N31734);
and and19173(N31730,N31735,N31736);
and and19174(N31731,R4,N31737);
and and19175(N31732,N31738,N31739);
and and17744(N29441,N29448,N29449);
and and17745(N29442,R4,R5);
and and17746(N29443,N29450,N29451);
and and17754(N29459,N29465,N29466);
and and17755(N29460,N29467,R5);
and and17756(N29461,N29468,N29469);
and and17764(N29477,N29483,N29484);
and and17765(N29478,N29485,R5);
and and17766(N29479,R6,N29486);
and and17774(N29494,N29500,N29501);
and and17775(N29495,N29502,R5);
and and17776(N29496,R6,N29503);
and and17784(N29511,R2,R3);
and and17785(N29512,N29518,N29519);
and and17786(N29513,R6,R7);
and and17794(N29527,R2,R3);
and and17795(N29528,R4,N29534);
and and17796(N29529,R6,N29535);
and and17804(N29543,R2,R3);
and and17805(N29544,N29549,R5);
and and17806(N29545,R6,R7);
and and17814(N29557,R3,N29565);
and and17815(N29558,N29566,N29567);
and and17823(N29575,N29582,N29583);
and and17824(N29576,N29584,N29585);
and and17832(N29593,N29600,N29601);
and and17833(N29594,N29602,N29603);
and and17841(N29611,N29617,N29618);
and and17842(N29612,N29619,N29620);
and and17850(N29628,N29635,N29636);
and and17851(N29629,N29637,R7);
and and17859(N29645,R3,N29652);
and and17860(N29646,N29653,N29654);
and and17868(N29662,N29668,N29669);
and and17869(N29663,N29670,N29671);
and and17877(N29679,N29686,N29687);
and and17878(N29680,R6,N29688);
and and17886(N29696,N29703,N29704);
and and17887(N29697,R6,N29705);
and and17895(N29713,R4,R5);
and and17896(N29714,N29720,N29721);
and and17904(N29729,N29735,R5);
and and17905(N29730,N29736,N29737);
and and17913(N29745,R4,N29751);
and and17914(N29746,N29752,N29753);
and and17922(N29761,R4,R5);
and and17923(N29762,N29768,N29769);
and and17931(N29777,N29783,N29784);
and and17932(N29778,N29785,R7);
and and17940(N29793,N29798,N29799);
and and17941(N29794,N29800,N29801);
and and17949(N29809,N29816,R5);
and and17950(N29810,N29817,R7);
and and17958(N29825,R4,N29832);
and and17959(N29826,N29833,R7);
and and17967(N29841,N29847,R5);
and and17968(N29842,N29848,N29849);
and and17976(N29857,R4,N29863);
and and17977(N29858,N29864,N29865);
and and17985(N29873,N29880,R5);
and and17986(N29874,R6,N29881);
and and17994(N29889,N29896,R4);
and and17995(N29890,R6,N29897);
and and18003(N29905,R4,N29911);
and and18004(N29906,N29912,N29913);
and and18012(N29921,N29927,N29928);
and and18013(N29922,N29929,R7);
and and18021(N29937,R4,N29944);
and and18022(N29938,N29945,R7);
and and18030(N29953,N29959,R5);
and and18031(N29954,N29960,N29961);
and and18039(N29969,N29975,N29976);
and and18040(N29970,R6,N29977);
and and18048(N29985,N29991,N29992);
and and18049(N29986,N29993,R7);
and and18057(N30001,N30007,N30008);
and and18058(N30002,R6,R7);
and and18066(N30016,N30021,N30022);
and and18067(N30017,N30023,R7);
and and18075(N30031,R3,N30036);
and and18076(N30032,N30037,N30038);
and and18084(N30046,N30051,R5);
and and18085(N30047,N30052,N30053);
and and18093(N30061,N30066,N30067);
and and18094(N30062,N30068,R7);
and and18102(N30076,R4,N30081);
and and18103(N30077,N30082,N30083);
and and18111(N30091,R3,R4);
and and18112(N30092,N30098,R6);
and and18120(N30106,R3,R5);
and and18121(N30107,N30112,N30113);
and and18129(N30121,R4,N30126);
and and18130(N30122,N30127,N30128);
and and18138(N30136,N30140,N30141);
and and18139(N30137,N30142,N30143);
and and18147(N30151,R3,N30156);
and and18148(N30152,N30157,N30158);
and and18156(N30166,N30171,N30172);
and and18157(N30167,R5,N30173);
and and18165(N30181,N30186,R4);
and and18166(N30182,N30187,N30188);
and and18174(N30196,N30201,N30202);
and and18175(N30197,R6,N30203);
and and18183(N30211,R3,N30216);
and and18184(N30212,N30217,N30218);
and and18192(N30226,N30232,R5);
and and18193(N30227,R6,N30233);
and and18201(N30241,N30246,R5);
and and18202(N30242,N30247,N30248);
and and18210(N30256,R4,N30261);
and and18211(N30257,N30262,N30263);
and and18219(N30271,R4,N30276);
and and18220(N30272,N30277,N30278);
and and18228(N30286,R4,N30292);
and and18229(N30287,N30293,R7);
and and18237(N30301,R4,N30307);
and and18238(N30302,N30308,R7);
and and18246(N30316,N30322,N30323);
and and18247(N30317,R6,R7);
and and18255(N30331,N30336,N30337);
and and18256(N30332,R6,N30338);
and and18264(N30346,N30351,N30352);
and and18265(N30347,N30353,R7);
and and18273(N30361,R3,R5);
and and18274(N30362,N30367,N30368);
and and18282(N30376,N30381,N30382);
and and18283(N30377,R6,N30383);
and and18291(N30391,R4,N30397);
and and18292(N30392,R6,N30398);
and and18300(N30406,N30411,R5);
and and18301(N30407,N30412,N30413);
and and18309(N30421,R4,N30426);
and and18310(N30422,N30427,N30428);
and and18318(N30436,R3,N30441);
and and18319(N30437,N30442,N30443);
and and18327(N30451,N30456,N30457);
and and18328(N30452,N30458,R7);
and and18336(N30466,R3,N30472);
and and18337(N30467,R6,N30473);
and and18345(N30481,R4,N30485);
and and18346(N30482,N30486,N30487);
and and18354(N30495,R4,R5);
and and18355(N30496,N30500,N30501);
and and18363(N30509,R4,N30514);
and and18364(N30510,R6,N30515);
and and18372(N30523,R3,N30528);
and and18373(N30524,N30529,R6);
and and18381(N30537,R4,R5);
and and18382(N30538,N30542,N30543);
and and18390(N30551,R4,R5);
and and18391(N30552,N30557,R7);
and and18399(N30565,R4,R5);
and and18400(N30566,N30571,R7);
and and18408(N30579,N30584,R5);
and and18409(N30580,R6,N30585);
and and18417(N30593,R4,R5);
and and18418(N30594,N30598,N30599);
and and18426(N30607,N30612,R5);
and and18427(N30608,N30613,R7);
and and18435(N30621,N30626,N30627);
and and18436(N30622,R6,R7);
and and18444(N30635,N30640,N30641);
and and18445(N30636,R6,R7);
and and18453(N30649,N30654,R5);
and and18454(N30650,N30655,R7);
and and18462(N30663,R4,R5);
and and18463(N30664,N30669,R7);
and and18471(N30677,R4,N30682);
and and18472(N30678,R6,N30683);
and and18480(N30691,N30695,R5);
and and18481(N30692,N30696,N30697);
and and18489(N30705,R3,N30710);
and and18490(N30706,R5,N30711);
and and18498(N30719,R3,R4);
and and18499(N30720,N30725,R7);
and and18507(N30733,N30738,R5);
and and18508(N30734,R6,N30739);
and and18516(N30747,R4,N30753);
and and18517(N30748,R6,R7);
and and18525(N30761,R4,N30767);
and and18526(N30762,R6,R7);
and and18534(N30775,R4,N30780);
and and18535(N30776,R6,N30781);
and and18543(N30789,N30795,R4);
and and18544(N30790,R5,R7);
and and18552(N30803,R4,N30808);
and and18553(N30804,N30809,R7);
and and18561(N30817,R4,N30822);
and and18562(N30818,N30823,R7);
and and18570(N30831,N30835,N30836);
and and18571(N30832,R5,N30837);
and and18579(N30845,R4,N30850);
and and18580(N30846,N30851,R7);
and and18588(N30859,R3,R4);
and and18589(N30860,R5,N30865);
and and18597(N30873,R3,R4);
and and18598(N30874,N30879,R7);
and and18606(N30887,R3,R4);
and and18607(N30888,N30893,R7);
and and18615(N30901,R4,N30906);
and and18616(N30902,N30907,R7);
and and18624(N30915,R4,N30920);
and and18625(N30916,N30921,R7);
and and18633(N30929,N30934,R4);
and and18634(N30930,N30935,R6);
and and18642(N30943,N30948,R4);
and and18643(N30944,N30949,R7);
and and18651(N30957,N30962,N30963);
and and18652(N30958,R6,R7);
and and18660(N30971,R4,N30976);
and and18661(N30972,R6,R7);
and and18669(N30984,N30987,N30988);
and and18670(N30985,N30989,R7);
and and18678(N30997,R4,R5);
and and18679(N30998,R6,N31002);
and and18687(N31010,R3,R5);
and and18688(N31011,N31014,N31015);
and and18696(N31023,N31026,N31027);
and and18697(N31024,N31028,R7);
and and18705(N31036,N31040,R5);
and and18706(N31037,N31041,R7);
and and18714(N31049,N31053,R5);
and and18715(N31050,R6,N31054);
and and18723(N31062,N31067,R5);
and and18724(N31063,R6,R7);
and and18732(N31075,R4,R5);
and and18733(N31076,R6,N31080);
and and18741(N31088,R4,N31093);
and and18742(N31089,R6,R7);
and and18750(N31101,R3,R4);
and and18751(N31102,N31106,R7);
and and18759(N31114,N31118,N31119);
and and18760(N31115,R6,R7);
and and18768(N31127,R4,N31132);
and and18769(N31128,R6,R7);
and and18777(N31140,N31144,R4);
and and18778(N31141,R6,N31145);
and and18786(N31153,N31157,R4);
and and18787(N31154,R5,N31158);
and and18795(N31166,R3,N31171);
and and18796(N31167,R6,R7);
and and18804(N31179,R4,N31184);
and and18805(N31180,R6,R7);
and and18813(N31192,R4,N31196);
and and18814(N31193,N31197,R7);
and and18822(N31205,R3,R5);
and and18823(N31206,R6,N31210);
and and18831(N31218,N31222,R5);
and and18832(N31219,N31223,R7);
and and18840(N31231,R3,N31236);
and and18841(N31232,R5,R7);
and and18849(N31244,R4,R5);
and and18850(N31245,R6,R7);
and and18858(N31256,R3,N31260);
and and18859(N31257,R5,R7);
and and18867(N31268,N31271,N31272);
and and18868(N31269,R6,R7);
and and18876(N31280,R4,N31284);
and and18877(N31281,R6,R7);
and and18885(N31292,R3,N31295);
and and18886(N31293,N31296,R6);
and and18894(N31304,R3,R4);
and and18895(N31305,R5,R7);
and and18903(N31316,R4,R5);
and and18904(N31317,N31320,R7);
and and18912(N31328,R4,N31332);
and and18913(N31329,R6,R7);
and and18921(N31340,R4,N31344);
and and18922(N31341,R6,R7);
and and18930(N31352,R4,N31356);
and and18931(N31353,R6,R7);
and and18939(N31364,R4,R5);
and and18940(N31365,R6,R7);
and and18948(N31374,R4,R5);
and and18949(N31375,R6,R7);
and and18957(N31384,R3,R5);
and and18958(N31385,R6,R7);
and and18966(N31394,R3,R4);
and and18967(N31395,R5,R7);
and and18975(N31404,R4,R5);
and and18976(N31405,R6,R7);
and and18984(N31414,N31421,N31422);
and and18992(N31430,R6,N31438);
and and19000(N31446,N31453,N31454);
and and19008(N31462,N31468,N31469);
and and19016(N31477,N31483,N31484);
and and19024(N31492,N31498,N31499);
and and19032(N31507,N31512,N31513);
and and19040(N31521,N31527,R6);
and and19048(N31535,N31540,N31541);
and and19056(N31549,R6,N31555);
and and19064(N31563,N31569,R7);
and and19072(N31577,N31582,N31583);
and and19080(N31591,N31596,R6);
and and19088(N31604,R6,R7);
and and19096(N31617,N31622,R7);
and and19104(N31630,R6,R7);
and and19112(N31642,R6,N31646);
and and19120(N31654,R6,N31658);
and and19128(N31666,R5,N31670);
and and19136(N31678,R6,N31682);
and and19144(N31690,R6,R7);
and and19152(N31701,N31703,N31704);
and and19160(N31712,N31714,N31715);
and and19168(N31723,R6,N31725);
and and19176(N31912,N31913,N31914);
and and19186(N31929,N31930,N31931);
and and19196(N31945,N31946,N31947);
and and19206(N31960,N31961,N31962);
and and19216(N31975,N31976,N31977);
and and19225(N31993,N31994,N31995);
and and19234(N32011,N32012,N32013);
and and19243(N32029,N32030,N32031);
and and19252(N32046,N32047,N32048);
and and19261(N32063,N32064,N32065);
and and19270(N32080,N32081,N32082);
and and19279(N32097,N32098,N32099);
and and19288(N32114,N32115,N32116);
and and19297(N32131,N32132,N32133);
and and19306(N32148,N32149,N32150);
and and19315(N32165,N32166,N32167);
and and19324(N32182,N32183,N32184);
and and19333(N32199,N32200,N32201);
and and19342(N32216,N32217,N32218);
and and19351(N32233,N32234,N32235);
and and19360(N32250,N32251,N32252);
and and19369(N32266,N32267,N32268);
and and19378(N32282,N32283,N32284);
and and19387(N32298,N32299,N32300);
and and19396(N32314,N32315,N32316);
and and19405(N32330,N32331,N32332);
and and19414(N32346,N32347,N32348);
and and19423(N32362,N32363,N32364);
and and19432(N32378,N32379,N32380);
and and19441(N32394,N32395,N32396);
and and19450(N32410,N32411,N32412);
and and19459(N32426,N32427,N32428);
and and19468(N32442,N32443,N32444);
and and19477(N32458,N32459,N32460);
and and19486(N32474,N32475,N32476);
and and19495(N32490,N32491,N32492);
and and19504(N32506,N32507,N32508);
and and19513(N32522,N32523,N32524);
and and19522(N32538,N32539,N32540);
and and19531(N32554,N32555,N32556);
and and19540(N32570,N32571,N32572);
and and19549(N32586,N32587,N32588);
and and19558(N32602,N32603,N32604);
and and19567(N32617,N32618,N32619);
and and19576(N32632,N32633,N32634);
and and19585(N32647,N32648,N32649);
and and19594(N32662,N32663,N32664);
and and19603(N32677,N32678,N32679);
and and19612(N32692,N32693,N32694);
and and19621(N32707,N32708,N32709);
and and19630(N32722,N32723,N32724);
and and19639(N32737,N32738,N32739);
and and19648(N32752,N32753,N32754);
and and19657(N32767,N32768,N32769);
and and19666(N32782,N32783,N32784);
and and19675(N32797,N32798,N32799);
and and19684(N32812,N32813,N32814);
and and19693(N32827,N32828,N32829);
and and19702(N32842,N32843,N32844);
and and19711(N32857,N32858,N32859);
and and19720(N32872,N32873,N32874);
and and19729(N32887,N32888,N32889);
and and19738(N32902,N32903,N32904);
and and19747(N32917,N32918,N32919);
and and19756(N32932,N32933,N32934);
and and19765(N32947,N32948,N32949);
and and19774(N32962,N32963,N32964);
and and19783(N32977,N32978,N32979);
and and19792(N32992,N32993,N32994);
and and19801(N33007,N33008,N33009);
and and19810(N33022,N33023,N33024);
and and19819(N33037,N33038,N33039);
and and19828(N33052,N33053,N33054);
and and19837(N33067,N33068,N33069);
and and19846(N33082,N33083,N33084);
and and19855(N33097,N33098,N33099);
and and19864(N33112,N33113,N33114);
and and19873(N33127,N33128,N33129);
and and19882(N33141,N33142,N33143);
and and19891(N33155,N33156,N33157);
and and19900(N33169,N33170,N33171);
and and19909(N33183,N33184,N33185);
and and19918(N33197,N33198,N33199);
and and19927(N33211,N33212,N33213);
and and19936(N33225,N33226,N33227);
and and19945(N33239,N33240,N33241);
and and19954(N33253,N33254,N33255);
and and19963(N33267,N33268,N33269);
and and19972(N33281,N33282,N33283);
and and19981(N33295,N33296,N33297);
and and19990(N33309,N33310,N33311);
and and19999(N33323,N33324,N33325);
and and20008(N33337,N33338,N33339);
and and20017(N33351,N33352,N33353);
and and20026(N33365,N33366,N33367);
and and20035(N33379,N33380,N33381);
and and20044(N33393,N33394,N33395);
and and20053(N33407,N33408,N33409);
and and20062(N33421,N33422,N33423);
and and20071(N33435,N33436,N33437);
and and20080(N33449,N33450,N33451);
and and20089(N33463,N33464,N33465);
and and20098(N33477,N33478,N33479);
and and20107(N33491,N33492,N33493);
and and20116(N33505,N33506,N33507);
and and20125(N33519,N33520,N33521);
and and20134(N33533,N33534,N33535);
and and20143(N33547,N33548,N33549);
and and20152(N33561,N33562,N33563);
and and20161(N33575,N33576,N33577);
and and20170(N33589,N33590,N33591);
and and20179(N33602,N33603,N33604);
and and20188(N33615,N33616,N33617);
and and20197(N33628,N33629,N33630);
and and20206(N33641,N33642,N33643);
and and20215(N33654,N33655,N33656);
and and20224(N33667,N33668,N33669);
and and20233(N33680,N33681,N33682);
and and20242(N33693,N33694,N33695);
and and20251(N33706,N33707,N33708);
and and20260(N33719,N33720,N33721);
and and20269(N33732,N33733,N33734);
and and20278(N33745,N33746,N33747);
and and20287(N33758,N33759,N33760);
and and20296(N33771,N33772,N33773);
and and20305(N33784,N33785,N33786);
and and20314(N33797,N33798,N33799);
and and20323(N33810,N33811,N33812);
and and20332(N33823,N33824,N33825);
and and20341(N33836,N33837,N33838);
and and20350(N33849,N33850,N33851);
and and20359(N33862,N33863,N33864);
and and20368(N33874,N33875,N33876);
and and20377(N33886,N33887,N33888);
and and20386(N33898,N33899,N33900);
and and20395(N33910,N33911,N33912);
and and20404(N33922,N33923,N33924);
and and20413(N33934,N33935,N33936);
and and20422(N33946,N33947,N33948);
and and20431(N33958,N33959,N33960);
and and20440(N33970,N33971,N33972);
and and20449(N33982,N33983,N33984);
and and20458(N33994,N33995,N33996);
and and20467(N34006,N34007,N34008);
and and20476(N34018,N34019,N34020);
and and20485(N34030,N34031,N34032);
and and20494(N34042,N34043,N34044);
and and20503(N34053,N34054,N34055);
and and20512(N34064,N34065,N34066);
and and20520(N34080,N34081,N34082);
and and20528(N34095,N34096,N34097);
and and20536(N34110,N34111,N34112);
and and20544(N34125,N34126,N34127);
and and20552(N34140,N34141,N34142);
and and20560(N34154,N34155,N34156);
and and20568(N34168,N34169,N34170);
and and20576(N34182,N34183,N34184);
and and20584(N34196,N34197,N34198);
and and20592(N34210,N34211,N34212);
and and20600(N34224,N34225,N34226);
and and20608(N34238,N34239,N34240);
and and20616(N34251,N34252,N34253);
and and20624(N34264,N34265,N34266);
and and20632(N34277,N34278,N34279);
and and20640(N34290,N34291,N34292);
and and20648(N34302,N34303,N34304);
and and20656(N34314,N34315,N34316);
and and20664(N34326,N34327,N34328);
and and20672(N34337,N34338,N34339);
and and20680(N34348,N34349,N34350);
and and20688(N34359,N34360,N34361);
and and20696(N34370,N34371,N34372);
and and20704(N34381,N34382,N34383);
and and19177(N31913,N31915,N31916);
and and19178(N31914,N31917,N31918);
and and19187(N31930,N31932,N31933);
and and19188(N31931,N31934,N31935);
and and19197(N31946,N31948,N31949);
and and19198(N31947,N31950,N31951);
and and19207(N31961,N31963,N31964);
and and19208(N31962,N31965,N31966);
and and19217(N31976,N31978,N31979);
and and19218(N31977,N31980,N31981);
and and19226(N31994,N31996,N31997);
and and19227(N31995,N31998,N31999);
and and19235(N32012,N32014,N32015);
and and19236(N32013,N32016,N32017);
and and19244(N32030,N32032,N32033);
and and19245(N32031,N32034,N32035);
and and19253(N32047,N32049,N32050);
and and19254(N32048,N32051,N32052);
and and19262(N32064,N32066,N32067);
and and19263(N32065,N32068,N32069);
and and19271(N32081,N32083,N32084);
and and19272(N32082,N32085,N32086);
and and19280(N32098,N32100,N32101);
and and19281(N32099,N32102,N32103);
and and19289(N32115,N32117,N32118);
and and19290(N32116,N32119,N32120);
and and19298(N32132,N32134,N32135);
and and19299(N32133,N32136,N32137);
and and19307(N32149,N32151,N32152);
and and19308(N32150,N32153,N32154);
and and19316(N32166,N32168,N32169);
and and19317(N32167,N32170,N32171);
and and19325(N32183,N32185,N32186);
and and19326(N32184,N32187,N32188);
and and19334(N32200,N32202,N32203);
and and19335(N32201,N32204,N32205);
and and19343(N32217,N32219,N32220);
and and19344(N32218,N32221,N32222);
and and19352(N32234,N32236,N32237);
and and19353(N32235,N32238,N32239);
and and19361(N32251,N32253,N32254);
and and19362(N32252,N32255,N32256);
and and19370(N32267,N32269,N32270);
and and19371(N32268,N32271,N32272);
and and19379(N32283,N32285,N32286);
and and19380(N32284,N32287,N32288);
and and19388(N32299,N32301,N32302);
and and19389(N32300,N32303,N32304);
and and19397(N32315,N32317,N32318);
and and19398(N32316,N32319,N32320);
and and19406(N32331,N32333,N32334);
and and19407(N32332,N32335,N32336);
and and19415(N32347,N32349,N32350);
and and19416(N32348,N32351,N32352);
and and19424(N32363,N32365,N32366);
and and19425(N32364,N32367,N32368);
and and19433(N32379,N32381,N32382);
and and19434(N32380,N32383,N32384);
and and19442(N32395,N32397,N32398);
and and19443(N32396,N32399,N32400);
and and19451(N32411,N32413,N32414);
and and19452(N32412,N32415,N32416);
and and19460(N32427,N32429,N32430);
and and19461(N32428,N32431,N32432);
and and19469(N32443,N32445,N32446);
and and19470(N32444,N32447,N32448);
and and19478(N32459,N32461,N32462);
and and19479(N32460,N32463,N32464);
and and19487(N32475,N32477,N32478);
and and19488(N32476,N32479,N32480);
and and19496(N32491,N32493,N32494);
and and19497(N32492,N32495,N32496);
and and19505(N32507,N32509,N32510);
and and19506(N32508,N32511,N32512);
and and19514(N32523,N32525,N32526);
and and19515(N32524,N32527,N32528);
and and19523(N32539,N32541,N32542);
and and19524(N32540,N32543,N32544);
and and19532(N32555,N32557,N32558);
and and19533(N32556,N32559,N32560);
and and19541(N32571,N32573,N32574);
and and19542(N32572,N32575,N32576);
and and19550(N32587,N32589,N32590);
and and19551(N32588,N32591,N32592);
and and19559(N32603,N32605,N32606);
and and19560(N32604,N32607,N32608);
and and19568(N32618,N32620,N32621);
and and19569(N32619,N32622,N32623);
and and19577(N32633,N32635,N32636);
and and19578(N32634,N32637,N32638);
and and19586(N32648,N32650,N32651);
and and19587(N32649,N32652,N32653);
and and19595(N32663,N32665,N32666);
and and19596(N32664,N32667,N32668);
and and19604(N32678,N32680,N32681);
and and19605(N32679,N32682,N32683);
and and19613(N32693,N32695,N32696);
and and19614(N32694,N32697,N32698);
and and19622(N32708,N32710,N32711);
and and19623(N32709,N32712,N32713);
and and19631(N32723,N32725,N32726);
and and19632(N32724,N32727,N32728);
and and19640(N32738,N32740,N32741);
and and19641(N32739,N32742,N32743);
and and19649(N32753,N32755,N32756);
and and19650(N32754,N32757,N32758);
and and19658(N32768,N32770,N32771);
and and19659(N32769,N32772,N32773);
and and19667(N32783,N32785,N32786);
and and19668(N32784,N32787,N32788);
and and19676(N32798,N32800,N32801);
and and19677(N32799,N32802,N32803);
and and19685(N32813,N32815,N32816);
and and19686(N32814,N32817,N32818);
and and19694(N32828,N32830,N32831);
and and19695(N32829,N32832,N32833);
and and19703(N32843,N32845,N32846);
and and19704(N32844,N32847,N32848);
and and19712(N32858,N32860,N32861);
and and19713(N32859,N32862,N32863);
and and19721(N32873,N32875,N32876);
and and19722(N32874,N32877,N32878);
and and19730(N32888,N32890,N32891);
and and19731(N32889,N32892,N32893);
and and19739(N32903,N32905,N32906);
and and19740(N32904,N32907,N32908);
and and19748(N32918,N32920,N32921);
and and19749(N32919,N32922,N32923);
and and19757(N32933,N32935,N32936);
and and19758(N32934,N32937,N32938);
and and19766(N32948,N32950,N32951);
and and19767(N32949,N32952,N32953);
and and19775(N32963,N32965,N32966);
and and19776(N32964,N32967,N32968);
and and19784(N32978,N32980,N32981);
and and19785(N32979,N32982,N32983);
and and19793(N32993,N32995,N32996);
and and19794(N32994,N32997,N32998);
and and19802(N33008,N33010,N33011);
and and19803(N33009,N33012,N33013);
and and19811(N33023,N33025,N33026);
and and19812(N33024,N33027,N33028);
and and19820(N33038,N33040,N33041);
and and19821(N33039,N33042,N33043);
and and19829(N33053,N33055,N33056);
and and19830(N33054,N33057,N33058);
and and19838(N33068,N33070,N33071);
and and19839(N33069,N33072,N33073);
and and19847(N33083,N33085,N33086);
and and19848(N33084,N33087,N33088);
and and19856(N33098,N33100,N33101);
and and19857(N33099,N33102,N33103);
and and19865(N33113,N33115,N33116);
and and19866(N33114,N33117,N33118);
and and19874(N33128,N33130,N33131);
and and19875(N33129,N33132,N33133);
and and19883(N33142,N33144,N33145);
and and19884(N33143,N33146,N33147);
and and19892(N33156,N33158,N33159);
and and19893(N33157,N33160,N33161);
and and19901(N33170,N33172,N33173);
and and19902(N33171,N33174,N33175);
and and19910(N33184,N33186,N33187);
and and19911(N33185,N33188,N33189);
and and19919(N33198,N33200,N33201);
and and19920(N33199,N33202,N33203);
and and19928(N33212,N33214,N33215);
and and19929(N33213,N33216,N33217);
and and19937(N33226,N33228,N33229);
and and19938(N33227,N33230,N33231);
and and19946(N33240,N33242,N33243);
and and19947(N33241,N33244,N33245);
and and19955(N33254,N33256,N33257);
and and19956(N33255,N33258,N33259);
and and19964(N33268,N33270,N33271);
and and19965(N33269,N33272,N33273);
and and19973(N33282,N33284,N33285);
and and19974(N33283,N33286,N33287);
and and19982(N33296,N33298,N33299);
and and19983(N33297,N33300,N33301);
and and19991(N33310,N33312,N33313);
and and19992(N33311,N33314,N33315);
and and20000(N33324,N33326,N33327);
and and20001(N33325,N33328,N33329);
and and20009(N33338,N33340,N33341);
and and20010(N33339,N33342,N33343);
and and20018(N33352,N33354,N33355);
and and20019(N33353,N33356,N33357);
and and20027(N33366,N33368,N33369);
and and20028(N33367,N33370,N33371);
and and20036(N33380,N33382,N33383);
and and20037(N33381,N33384,N33385);
and and20045(N33394,N33396,N33397);
and and20046(N33395,N33398,N33399);
and and20054(N33408,N33410,N33411);
and and20055(N33409,N33412,N33413);
and and20063(N33422,N33424,N33425);
and and20064(N33423,N33426,N33427);
and and20072(N33436,N33438,N33439);
and and20073(N33437,N33440,N33441);
and and20081(N33450,N33452,N33453);
and and20082(N33451,N33454,N33455);
and and20090(N33464,N33466,N33467);
and and20091(N33465,N33468,N33469);
and and20099(N33478,N33480,N33481);
and and20100(N33479,N33482,N33483);
and and20108(N33492,N33494,N33495);
and and20109(N33493,N33496,N33497);
and and20117(N33506,N33508,N33509);
and and20118(N33507,N33510,N33511);
and and20126(N33520,N33522,N33523);
and and20127(N33521,N33524,N33525);
and and20135(N33534,N33536,N33537);
and and20136(N33535,N33538,N33539);
and and20144(N33548,N33550,N33551);
and and20145(N33549,N33552,N33553);
and and20153(N33562,N33564,N33565);
and and20154(N33563,N33566,N33567);
and and20162(N33576,N33578,N33579);
and and20163(N33577,N33580,N33581);
and and20171(N33590,N33592,N33593);
and and20172(N33591,N33594,N33595);
and and20180(N33603,N33605,N33606);
and and20181(N33604,N33607,N33608);
and and20189(N33616,N33618,N33619);
and and20190(N33617,N33620,N33621);
and and20198(N33629,N33631,N33632);
and and20199(N33630,N33633,N33634);
and and20207(N33642,N33644,N33645);
and and20208(N33643,N33646,N33647);
and and20216(N33655,N33657,N33658);
and and20217(N33656,N33659,N33660);
and and20225(N33668,N33670,N33671);
and and20226(N33669,N33672,N33673);
and and20234(N33681,N33683,N33684);
and and20235(N33682,N33685,N33686);
and and20243(N33694,N33696,N33697);
and and20244(N33695,N33698,N33699);
and and20252(N33707,N33709,N33710);
and and20253(N33708,N33711,N33712);
and and20261(N33720,N33722,N33723);
and and20262(N33721,N33724,N33725);
and and20270(N33733,N33735,N33736);
and and20271(N33734,N33737,N33738);
and and20279(N33746,N33748,N33749);
and and20280(N33747,N33750,N33751);
and and20288(N33759,N33761,N33762);
and and20289(N33760,N33763,N33764);
and and20297(N33772,N33774,N33775);
and and20298(N33773,N33776,N33777);
and and20306(N33785,N33787,N33788);
and and20307(N33786,N33789,N33790);
and and20315(N33798,N33800,N33801);
and and20316(N33799,N33802,N33803);
and and20324(N33811,N33813,N33814);
and and20325(N33812,N33815,N33816);
and and20333(N33824,N33826,N33827);
and and20334(N33825,N33828,N33829);
and and20342(N33837,N33839,N33840);
and and20343(N33838,N33841,N33842);
and and20351(N33850,N33852,N33853);
and and20352(N33851,N33854,N33855);
and and20360(N33863,N33865,N33866);
and and20361(N33864,N33867,N33868);
and and20369(N33875,N33877,N33878);
and and20370(N33876,N33879,N33880);
and and20378(N33887,N33889,N33890);
and and20379(N33888,N33891,N33892);
and and20387(N33899,N33901,N33902);
and and20388(N33900,N33903,N33904);
and and20396(N33911,N33913,N33914);
and and20397(N33912,N33915,N33916);
and and20405(N33923,N33925,N33926);
and and20406(N33924,N33927,N33928);
and and20414(N33935,N33937,N33938);
and and20415(N33936,N33939,N33940);
and and20423(N33947,N33949,N33950);
and and20424(N33948,N33951,N33952);
and and20432(N33959,N33961,N33962);
and and20433(N33960,N33963,N33964);
and and20441(N33971,N33973,N33974);
and and20442(N33972,N33975,N33976);
and and20450(N33983,N33985,N33986);
and and20451(N33984,N33987,N33988);
and and20459(N33995,N33997,N33998);
and and20460(N33996,N33999,N34000);
and and20468(N34007,N34009,N34010);
and and20469(N34008,N34011,N34012);
and and20477(N34019,N34021,N34022);
and and20478(N34020,N34023,N34024);
and and20486(N34031,N34033,N34034);
and and20487(N34032,N34035,N34036);
and and20495(N34043,N34045,N34046);
and and20496(N34044,N34047,N34048);
and and20504(N34054,N34056,N34057);
and and20505(N34055,N34058,N34059);
and and20513(N34065,N34067,N34068);
and and20514(N34066,N34069,N34070);
and and20521(N34081,N34083,N34084);
and and20522(N34082,N34085,N34086);
and and20529(N34096,N34098,N34099);
and and20530(N34097,N34100,N34101);
and and20537(N34111,N34113,N34114);
and and20538(N34112,N34115,N34116);
and and20545(N34126,N34128,N34129);
and and20546(N34127,N34130,N34131);
and and20553(N34141,N34143,N34144);
and and20554(N34142,N34145,N34146);
and and20561(N34155,N34157,N34158);
and and20562(N34156,N34159,N34160);
and and20569(N34169,N34171,N34172);
and and20570(N34170,N34173,N34174);
and and20577(N34183,N34185,N34186);
and and20578(N34184,N34187,N34188);
and and20585(N34197,N34199,N34200);
and and20586(N34198,N34201,N34202);
and and20593(N34211,N34213,N34214);
and and20594(N34212,N34215,N34216);
and and20601(N34225,N34227,N34228);
and and20602(N34226,N34229,N34230);
and and20609(N34239,N34241,N34242);
and and20610(N34240,N34243,N34244);
and and20617(N34252,N34254,N34255);
and and20618(N34253,N34256,N34257);
and and20625(N34265,N34267,N34268);
and and20626(N34266,N34269,N34270);
and and20633(N34278,N34280,N34281);
and and20634(N34279,N34282,N34283);
and and20641(N34291,N34293,N34294);
and and20642(N34292,N34295,N34296);
and and20649(N34303,N34305,N34306);
and and20650(N34304,N34307,N34308);
and and20657(N34315,N34317,N34318);
and and20658(N34316,N34319,N34320);
and and20665(N34327,N34329,N34330);
and and20666(N34328,N34331,N34332);
and and20673(N34338,N34340,N34341);
and and20674(N34339,N34342,N34343);
and and20681(N34349,N34351,N34352);
and and20682(N34350,N34353,N34354);
and and20689(N34360,N34362,N34363);
and and20690(N34361,N34364,N34365);
and and20697(N34371,N34373,N34374);
and and20698(N34372,N34375,N34376);
and and20705(N34382,N34384,N34385);
and and20706(N34383,N34386,N34387);
and and19179(N31915,N31919,N31920);
and and19180(N31916,N31921,N31922);
and and19181(N31917,N31923,N31924);
and and19182(N31918,N31925,N31926);
and and19189(N31932,N31936,N31937);
and and19190(N31933,N31938,N31939);
and and19191(N31934,in1,N31940);
and and19192(N31935,R0,N31941);
and and19199(N31948,N31952,N31953);
and and19200(N31949,N31954,N31955);
and and19201(N31950,in1,in2);
and and19202(N31951,N31956,R1);
and and19209(N31963,N31967,N31968);
and and19210(N31964,N31969,N31970);
and and19211(N31965,in1,in2);
and and19212(N31966,N31971,N31972);
and and19219(N31978,N31982,N31983);
and and19220(N31979,N31984,N31985);
and and19221(N31980,N31986,R1);
and and19222(N31981,N31987,N31988);
and and19228(N31996,N32000,N32001);
and and19229(N31997,N32002,N32003);
and and19230(N31998,N32004,N32005);
and and19231(N31999,N32006,N32007);
and and19237(N32014,N32018,N32019);
and and19238(N32015,N32020,N32021);
and and19239(N32016,in2,N32022);
and and19240(N32017,N32023,N32024);
and and19246(N32032,N32036,N32037);
and and19247(N32033,N32038,N32039);
and and19248(N32034,N32040,N32041);
and and19249(N32035,N32042,N32043);
and and19255(N32049,N32053,N32054);
and and19256(N32050,N32055,in1);
and and19257(N32051,N32056,N32057);
and and19258(N32052,N32058,N32059);
and and19264(N32066,N32070,N32071);
and and19265(N32067,N32072,N32073);
and and19266(N32068,N32074,R1);
and and19267(N32069,R2,N32075);
and and19273(N32083,N32087,N32088);
and and19274(N32084,N32089,N32090);
and and19275(N32085,N32091,N32092);
and and19276(N32086,R2,R3);
and and19282(N32100,N32104,N32105);
and and19283(N32101,N32106,N32107);
and and19284(N32102,N32108,N32109);
and and19285(N32103,N32110,R3);
and and19291(N32117,N32121,N32122);
and and19292(N32118,N32123,in1);
and and19293(N32119,in2,N32124);
and and19294(N32120,N32125,N32126);
and and19300(N32134,N32138,N32139);
and and19301(N32135,N32140,N32141);
and and19302(N32136,N32142,N32143);
and and19303(N32137,R1,N32144);
and and19309(N32151,N32155,N32156);
and and19310(N32152,N32157,N32158);
and and19311(N32153,N32159,R0);
and and19312(N32154,N32160,N32161);
and and19318(N32168,N32172,N32173);
and and19319(N32169,N32174,N32175);
and and19320(N32170,N32176,R0);
and and19321(N32171,N32177,N32178);
and and19327(N32185,N32189,N32190);
and and19328(N32186,N32191,N32192);
and and19329(N32187,N32193,N32194);
and and19330(N32188,N32195,N32196);
and and19336(N32202,N32206,N32207);
and and19337(N32203,N32208,N32209);
and and19338(N32204,in2,R0);
and and19339(N32205,N32210,N32211);
and and19345(N32219,N32223,N32224);
and and19346(N32220,N32225,in1);
and and19347(N32221,N32226,R0);
and and19348(N32222,N32227,N32228);
and and19354(N32236,N32240,N32241);
and and19355(N32237,N32242,in1);
and and19356(N32238,N32243,N32244);
and and19357(N32239,R1,N32245);
and and19363(N32253,N32257,N32258);
and and19364(N32254,N32259,N32260);
and and19365(N32255,in2,N32261);
and and19366(N32256,R1,N32262);
and and19372(N32269,N32273,N32274);
and and19373(N32270,N32275,in1);
and and19374(N32271,N32276,N32277);
and and19375(N32272,N32278,R3);
and and19381(N32285,N32289,N32290);
and and19382(N32286,N32291,in1);
and and19383(N32287,N32292,N32293);
and and19384(N32288,N32294,R3);
and and19390(N32301,N32305,N32306);
and and19391(N32302,N32307,N32308);
and and19392(N32303,in2,N32309);
and and19393(N32304,R2,N32310);
and and19399(N32317,N32321,N32322);
and and19400(N32318,N32323,in1);
and and19401(N32319,N32324,N32325);
and and19402(N32320,N32326,R2);
and and19408(N32333,N32337,N32338);
and and19409(N32334,N32339,in1);
and and19410(N32335,N32340,N32341);
and and19411(N32336,R2,R3);
and and19417(N32349,N32353,N32354);
and and19418(N32350,N32355,N32356);
and and19419(N32351,N32357,N32358);
and and19420(N32352,N32359,R3);
and and19426(N32365,N32369,N32370);
and and19427(N32366,N32371,N32372);
and and19428(N32367,N32373,N32374);
and and19429(N32368,N32375,R3);
and and19435(N32381,N32385,N32386);
and and19436(N32382,N32387,in2);
and and19437(N32383,N32388,N32389);
and and19438(N32384,R2,N32390);
and and19444(N32397,N32401,N32402);
and and19445(N32398,N32403,in1);
and and19446(N32399,N32404,N32405);
and and19447(N32400,R2,N32406);
and and19453(N32413,N32417,N32418);
and and19454(N32414,N32419,N32420);
and and19455(N32415,N32421,R0);
and and19456(N32416,N32422,N32423);
and and19462(N32429,N32433,N32434);
and and19463(N32430,N32435,N32436);
and and19464(N32431,N32437,N32438);
and and19465(N32432,R1,N32439);
and and19471(N32445,N32449,N32450);
and and19472(N32446,N32451,in2);
and and19473(N32447,R0,N32452);
and and19474(N32448,N32453,N32454);
and and19480(N32461,N32465,N32466);
and and19481(N32462,N32467,N32468);
and and19482(N32463,in2,R0);
and and19483(N32464,N32469,N32470);
and and19489(N32477,N32481,N32482);
and and19490(N32478,N32483,N32484);
and and19491(N32479,N32485,R1);
and and19492(N32480,R2,N32486);
and and19498(N32493,N32497,N32498);
and and19499(N32494,N32499,in1);
and and19500(N32495,in2,N32500);
and and19501(N32496,N32501,N32502);
and and19507(N32509,N32513,N32514);
and and19508(N32510,N32515,in1);
and and19509(N32511,N32516,N32517);
and and19510(N32512,R1,N32518);
and and19516(N32525,N32529,N32530);
and and19517(N32526,N32531,N32532);
and and19518(N32527,N32533,R0);
and and19519(N32528,R1,N32534);
and and19525(N32541,N32545,N32546);
and and19526(N32542,N32547,in1);
and and19527(N32543,in2,R0);
and and19528(N32544,N32548,N32549);
and and19534(N32557,N32561,N32562);
and and19535(N32558,N32563,N32564);
and and19536(N32559,N32565,N32566);
and and19537(N32560,R2,N32567);
and and19543(N32573,N32577,N32578);
and and19544(N32574,N32579,in1);
and and19545(N32575,N32580,N32581);
and and19546(N32576,N32582,N32583);
and and19552(N32589,N32593,N32594);
and and19553(N32590,N32595,N32596);
and and19554(N32591,in2,N32597);
and and19555(N32592,N32598,R2);
and and19561(N32605,N32609,N32610);
and and19562(N32606,N32611,in1);
and and19563(N32607,in2,N32612);
and and19564(N32608,N32613,N32614);
and and19570(N32620,N32624,N32625);
and and19571(N32621,N32626,in2);
and and19572(N32622,R0,N32627);
and and19573(N32623,N32628,R3);
and and19579(N32635,N32639,N32640);
and and19580(N32636,N32641,in1);
and and19581(N32637,N32642,R0);
and and19582(N32638,N32643,N32644);
and and19588(N32650,N32654,N32655);
and and19589(N32651,N32656,N32657);
and and19590(N32652,N32658,R1);
and and19591(N32653,N32659,R3);
and and19597(N32665,N32669,N32670);
and and19598(N32666,N32671,N32672);
and and19599(N32667,R0,N32673);
and and19600(N32668,R2,R3);
and and19606(N32680,N32684,N32685);
and and19607(N32681,N32686,N32687);
and and19608(N32682,in2,N32688);
and and19609(N32683,N32689,R3);
and and19615(N32695,N32699,N32700);
and and19616(N32696,N32701,in1);
and and19617(N32697,N32702,N32703);
and and19618(N32698,N32704,R3);
and and19624(N32710,N32714,N32715);
and and19625(N32711,N32716,in1);
and and19626(N32712,N32717,N32718);
and and19627(N32713,R1,N32719);
and and19633(N32725,N32729,N32730);
and and19634(N32726,N32731,N32732);
and and19635(N32727,R0,R1);
and and19636(N32728,N32733,R3);
and and19642(N32740,N32744,N32745);
and and19643(N32741,N32746,N32747);
and and19644(N32742,in2,N32748);
and and19645(N32743,R2,N32749);
and and19651(N32755,N32759,N32760);
and and19652(N32756,N32761,in1);
and and19653(N32757,in2,N32762);
and and19654(N32758,N32763,R3);
and and19660(N32770,N32774,N32775);
and and19661(N32771,N32776,in1);
and and19662(N32772,N32777,R0);
and and19663(N32773,R1,N32778);
and and19669(N32785,N32789,N32790);
and and19670(N32786,N32791,N32792);
and and19671(N32787,in2,N32793);
and and19672(N32788,R1,R2);
and and19678(N32800,N32804,N32805);
and and19679(N32801,N32806,N32807);
and and19680(N32802,N32808,R0);
and and19681(N32803,R1,N32809);
and and19687(N32815,N32819,N32820);
and and19688(N32816,N32821,N32822);
and and19689(N32817,N32823,R1);
and and19690(N32818,R2,N32824);
and and19696(N32830,N32834,N32835);
and and19697(N32831,N32836,N32837);
and and19698(N32832,N32838,R1);
and and19699(N32833,N32839,N32840);
and and19705(N32845,N32849,N32850);
and and19706(N32846,N32851,in1);
and and19707(N32847,in2,R0);
and and19708(N32848,N32852,N32853);
and and19714(N32860,N32864,N32865);
and and19715(N32861,N32866,N32867);
and and19716(N32862,in2,N32868);
and and19717(N32863,N32869,R3);
and and19723(N32875,N32879,N32880);
and and19724(N32876,N32881,N32882);
and and19725(N32877,N32883,N32884);
and and19726(N32878,R2,R3);
and and19732(N32890,N32894,N32895);
and and19733(N32891,N32896,in1);
and and19734(N32892,N32897,R0);
and and19735(N32893,N32898,N32899);
and and19741(N32905,N32909,N32910);
and and19742(N32906,N32911,N32912);
and and19743(N32907,N32913,R0);
and and19744(N32908,N32914,R2);
and and19750(N32920,N32924,N32925);
and and19751(N32921,N32926,in1);
and and19752(N32922,in2,N32927);
and and19753(N32923,R1,N32928);
and and19759(N32935,N32939,N32940);
and and19760(N32936,N32941,in1);
and and19761(N32937,N32942,R0);
and and19762(N32938,N32943,N32944);
and and19768(N32950,N32954,N32955);
and and19769(N32951,N32956,N32957);
and and19770(N32952,in2,R1);
and and19771(N32953,N32958,N32959);
and and19777(N32965,N32969,N32970);
and and19778(N32966,N32971,N32972);
and and19779(N32967,N32973,R0);
and and19780(N32968,R1,N32974);
and and19786(N32980,N32984,N32985);
and and19787(N32981,N32986,N32987);
and and19788(N32982,N32988,R1);
and and19789(N32983,N32989,N32990);
and and19795(N32995,N32999,N33000);
and and19796(N32996,N33001,N33002);
and and19797(N32997,N33003,R0);
and and19798(N32998,R2,R3);
and and19804(N33010,N33014,N33015);
and and19805(N33011,N33016,N33017);
and and19806(N33012,N33018,R0);
and and19807(N33013,R1,R2);
and and19813(N33025,N33029,N33030);
and and19814(N33026,N33031,N33032);
and and19815(N33027,N33033,R0);
and and19816(N33028,N33034,R3);
and and19822(N33040,N33044,N33045);
and and19823(N33041,N33046,N33047);
and and19824(N33042,N33048,R0);
and and19825(N33043,R1,N33049);
and and19831(N33055,N33059,N33060);
and and19832(N33056,N33061,N33062);
and and19833(N33057,N33063,R1);
and and19834(N33058,R2,R3);
and and19840(N33070,N33074,N33075);
and and19841(N33071,N33076,N33077);
and and19842(N33072,R0,R1);
and and19843(N33073,N33078,N33079);
and and19849(N33085,N33089,N33090);
and and19850(N33086,N33091,in1);
and and19851(N33087,N33092,N33093);
and and19852(N33088,N33094,R3);
and and19858(N33100,N33104,N33105);
and and19859(N33101,N33106,in1);
and and19860(N33102,in2,N33107);
and and19861(N33103,N33108,N33109);
and and19867(N33115,N33119,N33120);
and and19868(N33116,N33121,N33122);
and and19869(N33117,R0,R1);
and and19870(N33118,N33123,N33124);
and and19876(N33130,N33134,N33135);
and and19877(N33131,N33136,in2);
and and19878(N33132,R0,R1);
and and19879(N33133,N33137,N33138);
and and19885(N33144,N33148,N33149);
and and19886(N33145,N33150,in1);
and and19887(N33146,in2,R0);
and and19888(N33147,R1,N33151);
and and19894(N33158,N33162,N33163);
and and19895(N33159,N33164,N33165);
and and19896(N33160,in2,R0);
and and19897(N33161,R1,N33166);
and and19903(N33172,N33176,N33177);
and and19904(N33173,N33178,N33179);
and and19905(N33174,in2,R0);
and and19906(N33175,N33180,N33181);
and and19912(N33186,N33190,N33191);
and and19913(N33187,N33192,N33193);
and and19914(N33188,N33194,R1);
and and19915(N33189,N33195,R3);
and and19921(N33200,N33204,N33205);
and and19922(N33201,N33206,in1);
and and19923(N33202,N33207,N33208);
and and19924(N33203,R1,R3);
and and19930(N33214,N33218,N33219);
and and19931(N33215,N33220,N33221);
and and19932(N33216,in2,R0);
and and19933(N33217,R1,N33222);
and and19939(N33228,N33232,N33233);
and and19940(N33229,N33234,in1);
and and19941(N33230,R0,R1);
and and19942(N33231,N33235,R3);
and and19948(N33242,N33246,N33247);
and and19949(N33243,N33248,in1);
and and19950(N33244,in2,N33249);
and and19951(N33245,R1,N33250);
and and19957(N33256,N33260,N33261);
and and19958(N33257,N33262,in1);
and and19959(N33258,N33263,N33264);
and and19960(N33259,R1,N33265);
and and19966(N33270,N33274,N33275);
and and19967(N33271,N33276,N33277);
and and19968(N33272,R0,N33278);
and and19969(N33273,N33279,R3);
and and19975(N33284,N33288,N33289);
and and19976(N33285,N33290,in2);
and and19977(N33286,N33291,R1);
and and19978(N33287,R2,R3);
and and19984(N33298,N33302,N33303);
and and19985(N33299,N33304,N33305);
and and19986(N33300,N33306,R0);
and and19987(N33301,N33307,R3);
and and19993(N33312,N33316,N33317);
and and19994(N33313,N33318,N33319);
and and19995(N33314,N33320,R0);
and and19996(N33315,R1,R2);
and and20002(N33326,N33330,N33331);
and and20003(N33327,N33332,N33333);
and and20004(N33328,in2,N33334);
and and20005(N33329,R1,R2);
and and20011(N33340,N33344,N33345);
and and20012(N33341,N33346,in1);
and and20013(N33342,in2,R1);
and and20014(N33343,N33347,N33348);
and and20020(N33354,N33358,N33359);
and and20021(N33355,N33360,in1);
and and20022(N33356,in2,R0);
and and20023(N33357,N33361,N33362);
and and20029(N33368,N33372,N33373);
and and20030(N33369,N33374,in1);
and and20031(N33370,N33375,N33376);
and and20032(N33371,N33377,R3);
and and20038(N33382,N33386,N33387);
and and20039(N33383,N33388,N33389);
and and20040(N33384,in2,R0);
and and20041(N33385,R2,R3);
and and20047(N33396,N33400,N33401);
and and20048(N33397,N33402,N33403);
and and20049(N33398,in2,R0);
and and20050(N33399,R1,N33404);
and and20056(N33410,N33414,N33415);
and and20057(N33411,N33416,N33417);
and and20058(N33412,N33418,R0);
and and20059(N33413,R1,N33419);
and and20065(N33424,N33428,N33429);
and and20066(N33425,N33430,N33431);
and and20067(N33426,R0,N33432);
and and20068(N33427,R2,N33433);
and and20074(N33438,N33442,N33443);
and and20075(N33439,N33444,N33445);
and and20076(N33440,in2,N33446);
and and20077(N33441,N33447,R2);
and and20083(N33452,N33456,N33457);
and and20084(N33453,N33458,in2);
and and20085(N33454,N33459,N33460);
and and20086(N33455,R2,R3);
and and20092(N33466,N33470,N33471);
and and20093(N33467,N33472,in1);
and and20094(N33468,in2,N33473);
and and20095(N33469,R1,R2);
and and20101(N33480,N33484,N33485);
and and20102(N33481,N33486,N33487);
and and20103(N33482,in2,R0);
and and20104(N33483,N33488,R2);
and and20110(N33494,N33498,N33499);
and and20111(N33495,N33500,in1);
and and20112(N33496,in2,N33501);
and and20113(N33497,N33502,R2);
and and20119(N33508,N33512,N33513);
and and20120(N33509,N33514,N33515);
and and20121(N33510,in2,R0);
and and20122(N33511,R1,N33516);
and and20128(N33522,N33526,N33527);
and and20129(N33523,N33528,N33529);
and and20130(N33524,in2,R0);
and and20131(N33525,R1,R2);
and and20137(N33536,N33540,N33541);
and and20138(N33537,N33542,N33543);
and and20139(N33538,in2,R0);
and and20140(N33539,N33544,N33545);
and and20146(N33550,N33554,N33555);
and and20147(N33551,N33556,N33557);
and and20148(N33552,N33558,N33559);
and and20149(N33553,R1,R2);
and and20155(N33564,N33568,N33569);
and and20156(N33565,N33570,in1);
and and20157(N33566,N33571,N33572);
and and20158(N33567,R2,R3);
and and20164(N33578,N33582,N33583);
and and20165(N33579,N33584,in2);
and and20166(N33580,N33585,N33586);
and and20167(N33581,R2,N33587);
and and20173(N33592,N33596,N33597);
and and20174(N33593,N33598,N33599);
and and20175(N33594,N33600,R0);
and and20176(N33595,R1,N33601);
and and20182(N33605,N33609,N33610);
and and20183(N33606,N33611,N33612);
and and20184(N33607,N33613,R0);
and and20185(N33608,R1,R2);
and and20191(N33618,N33622,N33623);
and and20192(N33619,N33624,in1);
and and20193(N33620,N33625,R1);
and and20194(N33621,R2,R3);
and and20200(N33631,N33635,N33636);
and and20201(N33632,N33637,in1);
and and20202(N33633,in2,R0);
and and20203(N33634,R1,N33638);
and and20209(N33644,N33648,N33649);
and and20210(N33645,N33650,in1);
and and20211(N33646,in2,R0);
and and20212(N33647,N33651,R2);
and and20218(N33657,N33661,N33662);
and and20219(N33658,N33663,in1);
and and20220(N33659,in2,R0);
and and20221(N33660,R1,N33664);
and and20227(N33670,N33674,N33675);
and and20228(N33671,N33676,in1);
and and20229(N33672,in2,R0);
and and20230(N33673,N33677,R3);
and and20236(N33683,N33687,N33688);
and and20237(N33684,N33689,N33690);
and and20238(N33685,in2,N33691);
and and20239(N33686,R2,R3);
and and20245(N33696,N33700,N33701);
and and20246(N33697,N33702,in1);
and and20247(N33698,N33703,R0);
and and20248(N33699,R1,R2);
and and20254(N33709,N33713,N33714);
and and20255(N33710,N33715,N33716);
and and20256(N33711,N33717,R0);
and and20257(N33712,N33718,R2);
and and20263(N33722,N33726,N33727);
and and20264(N33723,N33728,N33729);
and and20265(N33724,N33730,R0);
and and20266(N33725,R1,N33731);
and and20272(N33735,N33739,N33740);
and and20273(N33736,N33741,in1);
and and20274(N33737,R0,N33742);
and and20275(N33738,R2,N33743);
and and20281(N33748,N33752,N33753);
and and20282(N33749,N33754,N33755);
and and20283(N33750,N33756,R1);
and and20284(N33751,R2,R3);
and and20290(N33761,N33765,N33766);
and and20291(N33762,N33767,in1);
and and20292(N33763,N33768,R1);
and and20293(N33764,N33769,R3);
and and20299(N33774,N33778,N33779);
and and20300(N33775,N33780,in1);
and and20301(N33776,N33781,R1);
and and20302(N33777,R2,N33782);
and and20308(N33787,N33791,N33792);
and and20309(N33788,N33793,in1);
and and20310(N33789,in2,R0);
and and20311(N33790,R1,R2);
and and20317(N33800,N33804,N33805);
and and20318(N33801,N33806,in1);
and and20319(N33802,in2,R0);
and and20320(N33803,N33807,R3);
and and20326(N33813,N33817,N33818);
and and20327(N33814,N33819,in1);
and and20328(N33815,in2,N33820);
and and20329(N33816,R1,N33821);
and and20335(N33826,N33830,N33831);
and and20336(N33827,N33832,N33833);
and and20337(N33828,R0,R1);
and and20338(N33829,R2,R3);
and and20344(N33839,N33843,N33844);
and and20345(N33840,N33845,in1);
and and20346(N33841,in2,R0);
and and20347(N33842,R1,N33846);
and and20353(N33852,N33856,N33857);
and and20354(N33853,N33858,in1);
and and20355(N33854,in2,R0);
and and20356(N33855,R1,N33859);
and and20362(N33865,N33869,N33870);
and and20363(N33866,N33871,N33872);
and and20364(N33867,in2,R0);
and and20365(N33868,R1,R2);
and and20371(N33877,N33881,N33882);
and and20372(N33878,N33883,N33884);
and and20373(N33879,R0,R1);
and and20374(N33880,R2,R3);
and and20380(N33889,N33893,N33894);
and and20381(N33890,N33895,N33896);
and and20382(N33891,in2,R1);
and and20383(N33892,R2,N33897);
and and20389(N33901,N33905,N33906);
and and20390(N33902,N33907,in1);
and and20391(N33903,N33908,N33909);
and and20392(N33904,R1,R2);
and and20398(N33913,N33917,N33918);
and and20399(N33914,N33919,in1);
and and20400(N33915,in2,N33920);
and and20401(N33916,R1,R2);
and and20407(N33925,N33929,N33930);
and and20408(N33926,N33931,in1);
and and20409(N33927,in2,R0);
and and20410(N33928,R1,R2);
and and20416(N33937,N33941,N33942);
and and20417(N33938,N33943,in1);
and and20418(N33939,N33944,N33945);
and and20419(N33940,R2,R3);
and and20425(N33949,N33953,N33954);
and and20426(N33950,N33955,in1);
and and20427(N33951,in2,R0);
and and20428(N33952,R1,R2);
and and20434(N33961,N33965,N33966);
and and20435(N33962,N33967,in2);
and and20436(N33963,R0,R1);
and and20437(N33964,R2,R3);
and and20443(N33973,N33977,N33978);
and and20444(N33974,N33979,in1);
and and20445(N33975,in2,R0);
and and20446(N33976,N33980,R2);
and and20452(N33985,N33989,N33990);
and and20453(N33986,N33991,in2);
and and20454(N33987,N33992,R1);
and and20455(N33988,R2,R3);
and and20461(N33997,N34001,N34002);
and and20462(N33998,N34003,in1);
and and20463(N33999,R0,R1);
and and20464(N34000,R2,N34004);
and and20470(N34009,N34013,N34014);
and and20471(N34010,N34015,in2);
and and20472(N34011,R0,N34016);
and and20473(N34012,R2,R3);
and and20479(N34021,N34025,N34026);
and and20480(N34022,N34027,in1);
and and20481(N34023,in2,R0);
and and20482(N34024,R1,R2);
and and20488(N34033,N34037,N34038);
and and20489(N34034,N34039,in1);
and and20490(N34035,in2,R0);
and and20491(N34036,R1,R2);
and and20497(N34045,N34049,N34050);
and and20498(N34046,N34051,in1);
and and20499(N34047,in2,R0);
and and20500(N34048,R1,R3);
and and20506(N34056,N34060,N34061);
and and20507(N34057,N34062,in1);
and and20508(N34058,in2,R0);
and and20509(N34059,N34063,R2);
and and20515(N34067,N34071,N34072);
and and20516(N34068,N34073,N34074);
and and20517(N34069,N34075,R2);
and and20518(N34070,N34076,N34077);
and and20523(N34083,N34087,N34088);
and and20524(N34084,N34089,N34090);
and and20525(N34085,R2,N34091);
and and20526(N34086,R4,N34092);
and and20531(N34098,N34102,N34103);
and and20532(N34099,N34104,in2);
and and20533(N34100,N34105,N34106);
and and20534(N34101,N34107,N34108);
and and20539(N34113,N34117,N34118);
and and20540(N34114,N34119,R0);
and and20541(N34115,N34120,R2);
and and20542(N34116,N34121,N34122);
and and20547(N34128,N34132,N34133);
and and20548(N34129,N34134,in2);
and and20549(N34130,N34135,N34136);
and and20550(N34131,R4,N34137);
and and20555(N34143,N34147,N34148);
and and20556(N34144,N34149,N34150);
and and20557(N34145,N34151,R1);
and and20558(N34146,N34152,R3);
and and20563(N34157,N34161,N34162);
and and20564(N34158,N34163,N34164);
and and20565(N34159,R0,R1);
and and20566(N34160,N34165,R4);
and and20571(N34171,N34175,N34176);
and and20572(N34172,N34177,in2);
and and20573(N34173,N34178,R1);
and and20574(N34174,N34179,N34180);
and and20579(N34185,N34189,N34190);
and and20580(N34186,N34191,N34192);
and and20581(N34187,N34193,R3);
and and20582(N34188,R4,N34194);
and and20587(N34199,N34203,N34204);
and and20588(N34200,N34205,N34206);
and and20589(N34201,N34207,R3);
and and20590(N34202,N34208,R5);
and and20595(N34213,N34217,N34218);
and and20596(N34214,N34219,N34220);
and and20597(N34215,R1,R2);
and and20598(N34216,N34221,R5);
and and20603(N34227,N34231,N34232);
and and20604(N34228,N34233,in2);
and and20605(N34229,N34234,N34235);
and and20606(N34230,R4,N34236);
and and20611(N34241,N34245,N34246);
and and20612(N34242,in2,R0);
and and20613(N34243,R1,R2);
and and20614(N34244,N34247,N34248);
and and20619(N34254,N34258,N34259);
and and20620(N34255,in1,R0);
and and20621(N34256,N34260,R2);
and and20622(N34257,N34261,N34262);
and and20627(N34267,N34271,N34272);
and and20628(N34268,N34273,in2);
and and20629(N34269,R0,R1);
and and20630(N34270,R2,N34274);
and and20635(N34280,N34284,N34285);
and and20636(N34281,N34286,R0);
and and20637(N34282,R1,R2);
and and20638(N34283,N34287,R5);
and and20643(N34293,N34297,N34298);
and and20644(N34294,N34299,N34300);
and and20645(N34295,R1,R2);
and and20646(N34296,R3,R4);
and and20651(N34305,N34309,N34310);
and and20652(N34306,in1,N34311);
and and20653(N34307,R0,R2);
and and20654(N34308,R4,N34312);
and and20659(N34317,N34321,N34322);
and and20660(N34318,in1,in2);
and and20661(N34319,R0,N34323);
and and20662(N34320,R2,R4);
and and20667(N34329,N34333,N34334);
and and20668(N34330,in1,in2);
and and20669(N34331,R1,R3);
and and20670(N34332,R4,R5);
and and20675(N34340,N34344,N34345);
and and20676(N34341,in1,N34346);
and and20677(N34342,R2,R3);
and and20678(N34343,R4,R5);
and and20683(N34351,N34355,N34356);
and and20684(N34352,N34357,in2);
and and20685(N34353,R1,R2);
and and20686(N34354,R3,R4);
and and20691(N34362,N34366,N34367);
and and20692(N34363,N34368,R1);
and and20693(N34364,N34369,R3);
and and20694(N34365,R4,R5);
and and20699(N34373,N34377,N34378);
and and20700(N34374,in1,R0);
and and20701(N34375,R2,R3);
and and20702(N34376,R4,R5);
and and20707(N34384,N34388,N34389);
and and20708(N34385,in1,N34390);
and and20709(N34386,R0,R2);
and and20710(N34387,R3,R4);
and and19183(N31919,R2,R3);
and and19184(N31920,R4,N31927);
and and19185(N31921,R6,N31928);
and and19193(N31936,R2,N31942);
and and19194(N31937,N31943,N31944);
and and19195(N31938,R6,R7);
and and19203(N31952,R2,N31957);
and and19204(N31953,R4,N31958);
and and19205(N31954,N31959,R7);
and and19213(N31967,R2,N31973);
and and19214(N31968,R4,R5);
and and19215(N31969,N31974,R7);
and and19223(N31982,N31989,N31990);
and and19224(N31983,N31991,N31992);
and and19232(N32000,N32008,N32009);
and and19233(N32001,N32010,R7);
and and19241(N32018,N32025,N32026);
and and19242(N32019,N32027,N32028);
and and19250(N32036,R4,R5);
and and19251(N32037,N32044,N32045);
and and19259(N32053,N32060,N32061);
and and19260(N32054,N32062,R7);
and and19268(N32070,N32076,N32077);
and and19269(N32071,N32078,N32079);
and and19277(N32087,N32093,N32094);
and and19278(N32088,N32095,N32096);
and and19286(N32104,N32111,N32112);
and and19287(N32105,R6,N32113);
and and19295(N32121,N32127,N32128);
and and19296(N32122,N32129,N32130);
and and19304(N32138,N32145,N32146);
and and19305(N32139,N32147,R6);
and and19313(N32155,R3,N32162);
and and19314(N32156,N32163,N32164);
and and19322(N32172,N32179,N32180);
and and19323(N32173,R6,N32181);
and and19331(N32189,R3,R5);
and and19332(N32190,N32197,N32198);
and and19340(N32206,N32212,N32213);
and and19341(N32207,N32214,N32215);
and and19349(N32223,N32229,N32230);
and and19350(N32224,N32231,N32232);
and and19358(N32240,N32246,N32247);
and and19359(N32241,N32248,N32249);
and and19367(N32257,R3,N32263);
and and19368(N32258,N32264,N32265);
and and19376(N32273,N32279,N32280);
and and19377(N32274,N32281,R7);
and and19385(N32289,R4,N32295);
and and19386(N32290,N32296,N32297);
and and19394(N32305,N32311,N32312);
and and19395(N32306,N32313,R7);
and and19403(N32321,N32327,N32328);
and and19404(N32322,N32329,R7);
and and19412(N32337,N32342,N32343);
and and19413(N32338,N32344,N32345);
and and19421(N32353,N32360,R5);
and and19422(N32354,N32361,R7);
and and19430(N32369,N32376,N32377);
and and19431(N32370,R6,R7);
and and19439(N32385,N32391,N32392);
and and19440(N32386,R6,N32393);
and and19448(N32401,N32407,N32408);
and and19449(N32402,R6,N32409);
and and19457(N32417,R4,N32424);
and and19458(N32418,N32425,R7);
and and19466(N32433,R4,N32440);
and and19467(N32434,N32441,R7);
and and19475(N32449,N32455,N32456);
and and19476(N32450,N32457,R7);
and and19484(N32465,R4,N32471);
and and19485(N32466,N32472,N32473);
and and19493(N32481,N32487,N32488);
and and19494(N32482,N32489,R7);
and and19502(N32497,R3,N32503);
and and19503(N32498,N32504,N32505);
and and19511(N32513,N32519,N32520);
and and19512(N32514,N32521,R7);
and and19520(N32529,N32535,N32536);
and and19521(N32530,R6,N32537);
and and19529(N32545,N32550,N32551);
and and19530(N32546,N32552,N32553);
and and19538(N32561,R4,N32568);
and and19539(N32562,N32569,R7);
and and19547(N32577,R4,R5);
and and19548(N32578,N32584,N32585);
and and19556(N32593,N32599,N32600);
and and19557(N32594,R5,N32601);
and and19565(N32609,R4,N32615);
and and19566(N32610,N32616,R7);
and and19574(N32624,N32629,R5);
and and19575(N32625,N32630,N32631);
and and19583(N32639,R3,R5);
and and19584(N32640,N32645,N32646);
and and19592(N32654,R4,R5);
and and19593(N32655,N32660,N32661);
and and19601(N32669,N32674,N32675);
and and19602(N32670,R6,N32676);
and and19610(N32684,R4,R5);
and and19611(N32685,N32690,N32691);
and and19619(N32699,R4,R5);
and and19620(N32700,N32705,N32706);
and and19628(N32714,R3,N32720);
and and19629(N32715,N32721,R6);
and and19637(N32729,N32734,N32735);
and and19638(N32730,N32736,R7);
and and19646(N32744,R4,R5);
and and19647(N32745,N32750,N32751);
and and19655(N32759,N32764,N32765);
and and19656(N32760,R6,N32766);
and and19664(N32774,N32779,R4);
and and19665(N32775,N32780,N32781);
and and19673(N32789,N32794,R4);
and and19674(N32790,N32795,N32796);
and and19682(N32804,N32810,R5);
and and19683(N32805,N32811,R7);
and and19691(N32819,N32825,R5);
and and19692(N32820,R6,N32826);
and and19700(N32834,R4,R5);
and and19701(N32835,R6,N32841);
and and19709(N32849,N32854,N32855);
and and19710(N32850,R6,N32856);
and and19718(N32864,N32870,N32871);
and and19719(N32865,R6,R7);
and and19727(N32879,R4,R5);
and and19728(N32880,N32885,N32886);
and and19736(N32894,R4,N32900);
and and19737(N32895,R6,N32901);
and and19745(N32909,R3,N32915);
and and19746(N32910,R5,N32916);
and and19754(N32924,N32929,R4);
and and19755(N32925,N32930,N32931);
and and19763(N32939,R3,R4);
and and19764(N32940,N32945,N32946);
and and19772(N32954,R4,N32960);
and and19773(N32955,N32961,R7);
and and19781(N32969,N32975,N32976);
and and19782(N32970,R6,R7);
and and19790(N32984,R4,R5);
and and19791(N32985,N32991,R7);
and and19799(N32999,N33004,N33005);
and and19800(N33000,N33006,R7);
and and19808(N33014,N33019,N33020);
and and19809(N33015,N33021,R7);
and and19817(N33029,R4,R5);
and and19818(N33030,N33035,N33036);
and and19826(N33044,R4,R5);
and and19827(N33045,N33050,N33051);
and and19835(N33059,N33064,R5);
and and19836(N33060,N33065,N33066);
and and19844(N33074,N33080,R5);
and and19845(N33075,N33081,R7);
and and19853(N33089,N33095,N33096);
and and19854(N33090,R6,R7);
and and19862(N33104,R3,R4);
and and19863(N33105,N33110,N33111);
and and19871(N33119,N33125,N33126);
and and19872(N33120,R6,R7);
and and19880(N33134,N33139,R5);
and and19881(N33135,R6,N33140);
and and19889(N33148,R3,N33152);
and and19890(N33149,N33153,N33154);
and and19898(N33162,R3,R4);
and and19899(N33163,N33167,N33168);
and and19907(N33176,R3,R5);
and and19908(N33177,N33182,R7);
and and19916(N33190,R4,N33196);
and and19917(N33191,R6,R7);
and and19925(N33204,R4,N33209);
and and19926(N33205,R6,N33210);
and and19934(N33218,R3,N33223);
and and19935(N33219,N33224,R6);
and and19943(N33232,N33236,N33237);
and and19944(N33233,R6,N33238);
and and19952(N33246,R3,N33251);
and and19953(N33247,N33252,R7);
and and19961(N33260,R4,N33266);
and and19962(N33261,R6,R7);
and and19970(N33274,R4,R5);
and and19971(N33275,R6,N33280);
and and19979(N33288,N33292,N33293);
and and19980(N33289,R6,N33294);
and and19988(N33302,R4,N33308);
and and19989(N33303,R6,R7);
and and19997(N33316,R3,N33321);
and and19998(N33317,R6,N33322);
and and20006(N33330,N33335,R5);
and and20007(N33331,R6,N33336);
and and20015(N33344,N33349,R5);
and and20016(N33345,R6,N33350);
and and20024(N33358,R4,R5);
and and20025(N33359,N33363,N33364);
and and20033(N33372,R4,N33378);
and and20034(N33373,R6,R7);
and and20042(N33386,N33390,R5);
and and20043(N33387,N33391,N33392);
and and20051(N33400,N33405,R4);
and and20052(N33401,N33406,R6);
and and20060(N33414,R4,N33420);
and and20061(N33415,R6,R7);
and and20069(N33428,R4,N33434);
and and20070(N33429,R6,R7);
and and20078(N33442,R4,N33448);
and and20079(N33443,R6,R7);
and and20087(N33456,N33461,N33462);
and and20088(N33457,R6,R7);
and and20096(N33470,N33474,N33475);
and and20097(N33471,R6,N33476);
and and20105(N33484,R3,N33489);
and and20106(N33485,N33490,R7);
and and20114(N33498,R3,N33503);
and and20115(N33499,N33504,R7);
and and20123(N33512,R3,R5);
and and20124(N33513,N33517,N33518);
and and20132(N33526,N33530,N33531);
and and20133(N33527,N33532,R7);
and and20141(N33540,R3,R4);
and and20142(N33541,R5,N33546);
and and20150(N33554,R3,R5);
and and20151(N33555,R6,N33560);
and and20159(N33568,R4,N33573);
and and20160(N33569,N33574,R7);
and and20168(N33582,R4,N33588);
and and20169(N33583,R6,R7);
and and20177(N33596,R3,R4);
and and20178(N33597,R5,R7);
and and20186(N33609,R3,N33614);
and and20187(N33610,R5,R7);
and and20195(N33622,N33626,N33627);
and and20196(N33623,R6,R7);
and and20204(N33635,R4,N33639);
and and20205(N33636,N33640,R7);
and and20213(N33648,R3,N33652);
and and20214(N33649,R6,N33653);
and and20222(N33661,R3,N33665);
and and20223(N33662,N33666,R7);
and and20231(N33674,N33678,R5);
and and20232(N33675,R6,N33679);
and and20240(N33687,R4,R5);
and and20241(N33688,R6,N33692);
and and20249(N33700,R3,N33704);
and and20250(N33701,N33705,R7);
and and20258(N33713,R3,R5);
and and20259(N33714,R6,R7);
and and20267(N33726,R3,R5);
and and20268(N33727,R6,R7);
and and20276(N33739,R4,R5);
and and20277(N33740,R6,N33744);
and and20285(N33752,N33757,R5);
and and20286(N33753,R6,R7);
and and20294(N33765,R4,R5);
and and20295(N33766,N33770,R7);
and and20303(N33778,R4,R5);
and and20304(N33779,N33783,R7);
and and20312(N33791,N33794,N33795);
and and20313(N33792,N33796,R7);
and and20321(N33804,R4,N33808);
and and20322(N33805,N33809,R7);
and and20330(N33817,R3,N33822);
and and20331(N33818,R6,R7);
and and20339(N33830,N33834,R5);
and and20340(N33831,R6,N33835);
and and20348(N33843,N33847,R5);
and and20349(N33844,R6,N33848);
and and20357(N33856,R3,N33860);
and and20358(N33857,R6,N33861);
and and20366(N33869,N33873,R4);
and and20367(N33870,R5,R7);
and and20375(N33881,R4,N33885);
and and20376(N33882,R6,R7);
and and20384(N33893,R4,R5);
and and20385(N33894,R6,R7);
and and20393(N33905,R4,R5);
and and20394(N33906,R6,R7);
and and20402(N33917,R3,N33921);
and and20403(N33918,R5,R7);
and and20411(N33929,N33932,N33933);
and and20412(N33930,R5,R6);
and and20420(N33941,R4,R5);
and and20421(N33942,R6,R7);
and and20429(N33953,R3,R5);
and and20430(N33954,N33956,N33957);
and and20438(N33965,N33968,N33969);
and and20439(N33966,R6,R7);
and and20447(N33977,R3,R4);
and and20448(N33978,N33981,R6);
and and20456(N33989,R4,R5);
and and20457(N33990,R6,N33993);
and and20465(N34001,N34005,R5);
and and20466(N34002,R6,R7);
and and20474(N34013,R4,N34017);
and and20475(N34014,R6,R7);
and and20483(N34025,R4,R5);
and and20484(N34026,N34028,N34029);
and and20492(N34037,N34040,N34041);
and and20493(N34038,R6,R7);
and and20501(N34049,R4,R5);
and and20502(N34050,N34052,R7);
and and20510(N34060,R3,R5);
and and20511(N34061,R6,R7);
and and20519(N34071,N34078,N34079);
and and20527(N34087,N34093,N34094);
and and20535(N34102,R6,N34109);
and and20543(N34117,N34123,N34124);
and and20551(N34132,N34138,N34139);
and and20559(N34147,N34153,R7);
and and20567(N34161,N34166,N34167);
and and20575(N34175,R6,N34181);
and and20583(N34189,N34195,R7);
and and20591(N34203,R6,N34209);
and and20599(N34217,N34222,N34223);
and and20607(N34231,R6,N34237);
and and20615(N34245,N34249,N34250);
and and20623(N34258,R5,N34263);
and and20631(N34271,N34275,N34276);
and and20639(N34284,N34288,N34289);
and and20647(N34297,N34301,R7);
and and20655(N34309,R6,N34313);
and and20663(N34321,N34324,N34325);
and and20671(N34333,N34335,N34336);
and and20679(N34344,R6,N34347);
and and20687(N34355,R5,N34358);
and and20695(N34366,R6,R7);
and and20703(N34377,N34379,N34380);
and and20711(N34388,N34391,R6);
and and20712(N34582,N34583,N34584);
and and20722(N34602,N34603,N34604);
and and20732(N34620,N34621,N34622);
and and20742(N34637,N34638,N34639);
and and20751(N34655,N34656,N34657);
and and20760(N34673,N34674,N34675);
and and20769(N34691,N34692,N34693);
and and20778(N34709,N34710,N34711);
and and20787(N34727,N34728,N34729);
and and20796(N34744,N34745,N34746);
and and20805(N34761,N34762,N34763);
and and20814(N34778,N34779,N34780);
and and20823(N34794,N34795,N34796);
and and20832(N34810,N34811,N34812);
and and20841(N34826,N34827,N34828);
and and20850(N34842,N34843,N34844);
and and20859(N34858,N34859,N34860);
and and20868(N34874,N34875,N34876);
and and20877(N34890,N34891,N34892);
and and20886(N34906,N34907,N34908);
and and20895(N34922,N34923,N34924);
and and20904(N34938,N34939,N34940);
and and20913(N34954,N34955,N34956);
and and20922(N34970,N34971,N34972);
and and20931(N34986,N34987,N34988);
and and20940(N35002,N35003,N35004);
and and20949(N35018,N35019,N35020);
and and20958(N35034,N35035,N35036);
and and20967(N35050,N35051,N35052);
and and20976(N35066,N35067,N35068);
and and20985(N35082,N35083,N35084);
and and20994(N35098,N35099,N35100);
and and21003(N35114,N35115,N35116);
and and21012(N35130,N35131,N35132);
and and21021(N35146,N35147,N35148);
and and21030(N35161,N35162,N35163);
and and21039(N35176,N35177,N35178);
and and21048(N35191,N35192,N35193);
and and21057(N35206,N35207,N35208);
and and21066(N35221,N35222,N35223);
and and21075(N35236,N35237,N35238);
and and21084(N35251,N35252,N35253);
and and21093(N35266,N35267,N35268);
and and21102(N35281,N35282,N35283);
and and21111(N35296,N35297,N35298);
and and21120(N35311,N35312,N35313);
and and21129(N35326,N35327,N35328);
and and21138(N35341,N35342,N35343);
and and21147(N35356,N35357,N35358);
and and21156(N35371,N35372,N35373);
and and21165(N35386,N35387,N35388);
and and21174(N35401,N35402,N35403);
and and21183(N35416,N35417,N35418);
and and21192(N35431,N35432,N35433);
and and21201(N35446,N35447,N35448);
and and21210(N35461,N35462,N35463);
and and21219(N35476,N35477,N35478);
and and21228(N35491,N35492,N35493);
and and21237(N35506,N35507,N35508);
and and21246(N35521,N35522,N35523);
and and21255(N35536,N35537,N35538);
and and21264(N35551,N35552,N35553);
and and21273(N35566,N35567,N35568);
and and21282(N35581,N35582,N35583);
and and21291(N35596,N35597,N35598);
and and21300(N35610,N35611,N35612);
and and21309(N35624,N35625,N35626);
and and21318(N35638,N35639,N35640);
and and21327(N35652,N35653,N35654);
and and21336(N35666,N35667,N35668);
and and21345(N35680,N35681,N35682);
and and21354(N35694,N35695,N35696);
and and21363(N35708,N35709,N35710);
and and21372(N35722,N35723,N35724);
and and21381(N35736,N35737,N35738);
and and21390(N35750,N35751,N35752);
and and21399(N35764,N35765,N35766);
and and21408(N35778,N35779,N35780);
and and21417(N35792,N35793,N35794);
and and21426(N35806,N35807,N35808);
and and21435(N35820,N35821,N35822);
and and21444(N35834,N35835,N35836);
and and21453(N35848,N35849,N35850);
and and21462(N35862,N35863,N35864);
and and21471(N35876,N35877,N35878);
and and21480(N35890,N35891,N35892);
and and21489(N35904,N35905,N35906);
and and21498(N35918,N35919,N35920);
and and21507(N35932,N35933,N35934);
and and21516(N35946,N35947,N35948);
and and21525(N35960,N35961,N35962);
and and21534(N35974,N35975,N35976);
and and21543(N35988,N35989,N35990);
and and21552(N36002,N36003,N36004);
and and21561(N36016,N36017,N36018);
and and21570(N36030,N36031,N36032);
and and21579(N36044,N36045,N36046);
and and21588(N36058,N36059,N36060);
and and21597(N36072,N36073,N36074);
and and21606(N36086,N36087,N36088);
and and21615(N36100,N36101,N36102);
and and21624(N36114,N36115,N36116);
and and21633(N36128,N36129,N36130);
and and21642(N36142,N36143,N36144);
and and21651(N36156,N36157,N36158);
and and21660(N36170,N36171,N36172);
and and21669(N36184,N36185,N36186);
and and21678(N36197,N36198,N36199);
and and21687(N36210,N36211,N36212);
and and21696(N36223,N36224,N36225);
and and21705(N36236,N36237,N36238);
and and21714(N36249,N36250,N36251);
and and21723(N36262,N36263,N36264);
and and21732(N36275,N36276,N36277);
and and21741(N36288,N36289,N36290);
and and21750(N36301,N36302,N36303);
and and21759(N36314,N36315,N36316);
and and21768(N36327,N36328,N36329);
and and21777(N36340,N36341,N36342);
and and21786(N36353,N36354,N36355);
and and21795(N36366,N36367,N36368);
and and21804(N36379,N36380,N36381);
and and21813(N36392,N36393,N36394);
and and21822(N36405,N36406,N36407);
and and21831(N36418,N36419,N36420);
and and21840(N36431,N36432,N36433);
and and21849(N36444,N36445,N36446);
and and21858(N36457,N36458,N36459);
and and21867(N36470,N36471,N36472);
and and21876(N36483,N36484,N36485);
and and21885(N36496,N36497,N36498);
and and21894(N36509,N36510,N36511);
and and21903(N36522,N36523,N36524);
and and21912(N36535,N36536,N36537);
and and21921(N36548,N36549,N36550);
and and21930(N36561,N36562,N36563);
and and21939(N36574,N36575,N36576);
and and21948(N36587,N36588,N36589);
and and21957(N36600,N36601,N36602);
and and21966(N36613,N36614,N36615);
and and21975(N36626,N36627,N36628);
and and21984(N36639,N36640,N36641);
and and21993(N36651,N36652,N36653);
and and22002(N36663,N36664,N36665);
and and22011(N36675,N36676,N36677);
and and22020(N36687,N36688,N36689);
and and22029(N36699,N36700,N36701);
and and22038(N36711,N36712,N36713);
and and22047(N36723,N36724,N36725);
and and22056(N36735,N36736,N36737);
and and22065(N36747,N36748,N36749);
and and22074(N36758,N36759,N36760);
and and22083(N36769,N36770,N36771);
and and22092(N36780,N36781,N36782);
and and22101(N36791,N36792,N36793);
and and22110(N36802,N36803,N36804);
and and22119(N36813,N36814,N36815);
and and22127(N36828,N36829,N36830);
and and22135(N36843,N36844,N36845);
and and22143(N36858,N36859,N36860);
and and22151(N36873,N36874,N36875);
and and22159(N36888,N36889,N36890);
and and22167(N36902,N36903,N36904);
and and22175(N36916,N36917,N36918);
and and22183(N36930,N36931,N36932);
and and22191(N36944,N36945,N36946);
and and22199(N36958,N36959,N36960);
and and22207(N36972,N36973,N36974);
and and22215(N36986,N36987,N36988);
and and22223(N37000,N37001,N37002);
and and22231(N37014,N37015,N37016);
and and22239(N37028,N37029,N37030);
and and22247(N37042,N37043,N37044);
and and22255(N37055,N37056,N37057);
and and22263(N37068,N37069,N37070);
and and22271(N37081,N37082,N37083);
and and22279(N37094,N37095,N37096);
and and22287(N37107,N37108,N37109);
and and22295(N37119,N37120,N37121);
and and22303(N37131,N37132,N37133);
and and22311(N37143,N37144,N37145);
and and22319(N37155,N37156,N37157);
and and22327(N37167,N37168,N37169);
and and22335(N37179,N37180,N37181);
and and22343(N37190,N37191,N37192);
and and22351(N37201,N37202,N37203);
and and22359(N37212,N37213,N37214);
and and22367(N37222,N37223,N37224);
and and22375(N37232,N37233,N37234);
and and22383(N37242,N37243,N37244);
and and22390(N37253,N37254,N37255);
and and20713(N34583,N34585,N34586);
and and20714(N34584,N34587,N34588);
and and20723(N34603,N34605,N34606);
and and20724(N34604,N34607,N34608);
and and20733(N34621,N34623,N34624);
and and20734(N34622,N34625,N34626);
and and20743(N34638,N34640,N34641);
and and20744(N34639,N34642,N34643);
and and20752(N34656,N34658,N34659);
and and20753(N34657,N34660,N34661);
and and20761(N34674,N34676,N34677);
and and20762(N34675,N34678,N34679);
and and20770(N34692,N34694,N34695);
and and20771(N34693,N34696,N34697);
and and20779(N34710,N34712,N34713);
and and20780(N34711,N34714,N34715);
and and20788(N34728,N34730,N34731);
and and20789(N34729,N34732,N34733);
and and20797(N34745,N34747,N34748);
and and20798(N34746,N34749,N34750);
and and20806(N34762,N34764,N34765);
and and20807(N34763,N34766,N34767);
and and20815(N34779,N34781,N34782);
and and20816(N34780,N34783,N34784);
and and20824(N34795,N34797,N34798);
and and20825(N34796,N34799,N34800);
and and20833(N34811,N34813,N34814);
and and20834(N34812,N34815,N34816);
and and20842(N34827,N34829,N34830);
and and20843(N34828,N34831,N34832);
and and20851(N34843,N34845,N34846);
and and20852(N34844,N34847,N34848);
and and20860(N34859,N34861,N34862);
and and20861(N34860,N34863,N34864);
and and20869(N34875,N34877,N34878);
and and20870(N34876,N34879,N34880);
and and20878(N34891,N34893,N34894);
and and20879(N34892,N34895,N34896);
and and20887(N34907,N34909,N34910);
and and20888(N34908,N34911,N34912);
and and20896(N34923,N34925,N34926);
and and20897(N34924,N34927,N34928);
and and20905(N34939,N34941,N34942);
and and20906(N34940,N34943,N34944);
and and20914(N34955,N34957,N34958);
and and20915(N34956,N34959,N34960);
and and20923(N34971,N34973,N34974);
and and20924(N34972,N34975,N34976);
and and20932(N34987,N34989,N34990);
and and20933(N34988,N34991,N34992);
and and20941(N35003,N35005,N35006);
and and20942(N35004,N35007,N35008);
and and20950(N35019,N35021,N35022);
and and20951(N35020,N35023,N35024);
and and20959(N35035,N35037,N35038);
and and20960(N35036,N35039,N35040);
and and20968(N35051,N35053,N35054);
and and20969(N35052,N35055,N35056);
and and20977(N35067,N35069,N35070);
and and20978(N35068,N35071,N35072);
and and20986(N35083,N35085,N35086);
and and20987(N35084,N35087,N35088);
and and20995(N35099,N35101,N35102);
and and20996(N35100,N35103,N35104);
and and21004(N35115,N35117,N35118);
and and21005(N35116,N35119,N35120);
and and21013(N35131,N35133,N35134);
and and21014(N35132,N35135,N35136);
and and21022(N35147,N35149,N35150);
and and21023(N35148,N35151,N35152);
and and21031(N35162,N35164,N35165);
and and21032(N35163,N35166,N35167);
and and21040(N35177,N35179,N35180);
and and21041(N35178,N35181,N35182);
and and21049(N35192,N35194,N35195);
and and21050(N35193,N35196,N35197);
and and21058(N35207,N35209,N35210);
and and21059(N35208,N35211,N35212);
and and21067(N35222,N35224,N35225);
and and21068(N35223,N35226,N35227);
and and21076(N35237,N35239,N35240);
and and21077(N35238,N35241,N35242);
and and21085(N35252,N35254,N35255);
and and21086(N35253,N35256,N35257);
and and21094(N35267,N35269,N35270);
and and21095(N35268,N35271,N35272);
and and21103(N35282,N35284,N35285);
and and21104(N35283,N35286,N35287);
and and21112(N35297,N35299,N35300);
and and21113(N35298,N35301,N35302);
and and21121(N35312,N35314,N35315);
and and21122(N35313,N35316,N35317);
and and21130(N35327,N35329,N35330);
and and21131(N35328,N35331,N35332);
and and21139(N35342,N35344,N35345);
and and21140(N35343,N35346,N35347);
and and21148(N35357,N35359,N35360);
and and21149(N35358,N35361,N35362);
and and21157(N35372,N35374,N35375);
and and21158(N35373,N35376,N35377);
and and21166(N35387,N35389,N35390);
and and21167(N35388,N35391,N35392);
and and21175(N35402,N35404,N35405);
and and21176(N35403,N35406,N35407);
and and21184(N35417,N35419,N35420);
and and21185(N35418,N35421,N35422);
and and21193(N35432,N35434,N35435);
and and21194(N35433,N35436,N35437);
and and21202(N35447,N35449,N35450);
and and21203(N35448,N35451,N35452);
and and21211(N35462,N35464,N35465);
and and21212(N35463,N35466,N35467);
and and21220(N35477,N35479,N35480);
and and21221(N35478,N35481,N35482);
and and21229(N35492,N35494,N35495);
and and21230(N35493,N35496,N35497);
and and21238(N35507,N35509,N35510);
and and21239(N35508,N35511,N35512);
and and21247(N35522,N35524,N35525);
and and21248(N35523,N35526,N35527);
and and21256(N35537,N35539,N35540);
and and21257(N35538,N35541,N35542);
and and21265(N35552,N35554,N35555);
and and21266(N35553,N35556,N35557);
and and21274(N35567,N35569,N35570);
and and21275(N35568,N35571,N35572);
and and21283(N35582,N35584,N35585);
and and21284(N35583,N35586,N35587);
and and21292(N35597,N35599,N35600);
and and21293(N35598,N35601,N35602);
and and21301(N35611,N35613,N35614);
and and21302(N35612,N35615,N35616);
and and21310(N35625,N35627,N35628);
and and21311(N35626,N35629,N35630);
and and21319(N35639,N35641,N35642);
and and21320(N35640,N35643,N35644);
and and21328(N35653,N35655,N35656);
and and21329(N35654,N35657,N35658);
and and21337(N35667,N35669,N35670);
and and21338(N35668,N35671,N35672);
and and21346(N35681,N35683,N35684);
and and21347(N35682,N35685,N35686);
and and21355(N35695,N35697,N35698);
and and21356(N35696,N35699,N35700);
and and21364(N35709,N35711,N35712);
and and21365(N35710,N35713,N35714);
and and21373(N35723,N35725,N35726);
and and21374(N35724,N35727,N35728);
and and21382(N35737,N35739,N35740);
and and21383(N35738,N35741,N35742);
and and21391(N35751,N35753,N35754);
and and21392(N35752,N35755,N35756);
and and21400(N35765,N35767,N35768);
and and21401(N35766,N35769,N35770);
and and21409(N35779,N35781,N35782);
and and21410(N35780,N35783,N35784);
and and21418(N35793,N35795,N35796);
and and21419(N35794,N35797,N35798);
and and21427(N35807,N35809,N35810);
and and21428(N35808,N35811,N35812);
and and21436(N35821,N35823,N35824);
and and21437(N35822,N35825,N35826);
and and21445(N35835,N35837,N35838);
and and21446(N35836,N35839,N35840);
and and21454(N35849,N35851,N35852);
and and21455(N35850,N35853,N35854);
and and21463(N35863,N35865,N35866);
and and21464(N35864,N35867,N35868);
and and21472(N35877,N35879,N35880);
and and21473(N35878,N35881,N35882);
and and21481(N35891,N35893,N35894);
and and21482(N35892,N35895,N35896);
and and21490(N35905,N35907,N35908);
and and21491(N35906,N35909,N35910);
and and21499(N35919,N35921,N35922);
and and21500(N35920,N35923,N35924);
and and21508(N35933,N35935,N35936);
and and21509(N35934,N35937,N35938);
and and21517(N35947,N35949,N35950);
and and21518(N35948,N35951,N35952);
and and21526(N35961,N35963,N35964);
and and21527(N35962,N35965,N35966);
and and21535(N35975,N35977,N35978);
and and21536(N35976,N35979,N35980);
and and21544(N35989,N35991,N35992);
and and21545(N35990,N35993,N35994);
and and21553(N36003,N36005,N36006);
and and21554(N36004,N36007,N36008);
and and21562(N36017,N36019,N36020);
and and21563(N36018,N36021,N36022);
and and21571(N36031,N36033,N36034);
and and21572(N36032,N36035,N36036);
and and21580(N36045,N36047,N36048);
and and21581(N36046,N36049,N36050);
and and21589(N36059,N36061,N36062);
and and21590(N36060,N36063,N36064);
and and21598(N36073,N36075,N36076);
and and21599(N36074,N36077,N36078);
and and21607(N36087,N36089,N36090);
and and21608(N36088,N36091,N36092);
and and21616(N36101,N36103,N36104);
and and21617(N36102,N36105,N36106);
and and21625(N36115,N36117,N36118);
and and21626(N36116,N36119,N36120);
and and21634(N36129,N36131,N36132);
and and21635(N36130,N36133,N36134);
and and21643(N36143,N36145,N36146);
and and21644(N36144,N36147,N36148);
and and21652(N36157,N36159,N36160);
and and21653(N36158,N36161,N36162);
and and21661(N36171,N36173,N36174);
and and21662(N36172,N36175,N36176);
and and21670(N36185,N36187,N36188);
and and21671(N36186,N36189,N36190);
and and21679(N36198,N36200,N36201);
and and21680(N36199,N36202,N36203);
and and21688(N36211,N36213,N36214);
and and21689(N36212,N36215,N36216);
and and21697(N36224,N36226,N36227);
and and21698(N36225,N36228,N36229);
and and21706(N36237,N36239,N36240);
and and21707(N36238,N36241,N36242);
and and21715(N36250,N36252,N36253);
and and21716(N36251,N36254,N36255);
and and21724(N36263,N36265,N36266);
and and21725(N36264,N36267,N36268);
and and21733(N36276,N36278,N36279);
and and21734(N36277,N36280,N36281);
and and21742(N36289,N36291,N36292);
and and21743(N36290,N36293,N36294);
and and21751(N36302,N36304,N36305);
and and21752(N36303,N36306,N36307);
and and21760(N36315,N36317,N36318);
and and21761(N36316,N36319,N36320);
and and21769(N36328,N36330,N36331);
and and21770(N36329,N36332,N36333);
and and21778(N36341,N36343,N36344);
and and21779(N36342,N36345,N36346);
and and21787(N36354,N36356,N36357);
and and21788(N36355,N36358,N36359);
and and21796(N36367,N36369,N36370);
and and21797(N36368,N36371,N36372);
and and21805(N36380,N36382,N36383);
and and21806(N36381,N36384,N36385);
and and21814(N36393,N36395,N36396);
and and21815(N36394,N36397,N36398);
and and21823(N36406,N36408,N36409);
and and21824(N36407,N36410,N36411);
and and21832(N36419,N36421,N36422);
and and21833(N36420,N36423,N36424);
and and21841(N36432,N36434,N36435);
and and21842(N36433,N36436,N36437);
and and21850(N36445,N36447,N36448);
and and21851(N36446,N36449,N36450);
and and21859(N36458,N36460,N36461);
and and21860(N36459,N36462,N36463);
and and21868(N36471,N36473,N36474);
and and21869(N36472,N36475,N36476);
and and21877(N36484,N36486,N36487);
and and21878(N36485,N36488,N36489);
and and21886(N36497,N36499,N36500);
and and21887(N36498,N36501,N36502);
and and21895(N36510,N36512,N36513);
and and21896(N36511,N36514,N36515);
and and21904(N36523,N36525,N36526);
and and21905(N36524,N36527,N36528);
and and21913(N36536,N36538,N36539);
and and21914(N36537,N36540,N36541);
and and21922(N36549,N36551,N36552);
and and21923(N36550,N36553,N36554);
and and21931(N36562,N36564,N36565);
and and21932(N36563,N36566,N36567);
and and21940(N36575,N36577,N36578);
and and21941(N36576,N36579,N36580);
and and21949(N36588,N36590,N36591);
and and21950(N36589,N36592,N36593);
and and21958(N36601,N36603,N36604);
and and21959(N36602,N36605,N36606);
and and21967(N36614,N36616,N36617);
and and21968(N36615,N36618,N36619);
and and21976(N36627,N36629,N36630);
and and21977(N36628,N36631,N36632);
and and21985(N36640,N36642,N36643);
and and21986(N36641,N36644,N36645);
and and21994(N36652,N36654,N36655);
and and21995(N36653,N36656,N36657);
and and22003(N36664,N36666,N36667);
and and22004(N36665,N36668,N36669);
and and22012(N36676,N36678,N36679);
and and22013(N36677,N36680,N36681);
and and22021(N36688,N36690,N36691);
and and22022(N36689,N36692,N36693);
and and22030(N36700,N36702,N36703);
and and22031(N36701,N36704,N36705);
and and22039(N36712,N36714,N36715);
and and22040(N36713,N36716,N36717);
and and22048(N36724,N36726,N36727);
and and22049(N36725,N36728,N36729);
and and22057(N36736,N36738,N36739);
and and22058(N36737,N36740,N36741);
and and22066(N36748,N36750,N36751);
and and22067(N36749,N36752,N36753);
and and22075(N36759,N36761,N36762);
and and22076(N36760,N36763,N36764);
and and22084(N36770,N36772,N36773);
and and22085(N36771,N36774,N36775);
and and22093(N36781,N36783,N36784);
and and22094(N36782,N36785,N36786);
and and22102(N36792,N36794,N36795);
and and22103(N36793,N36796,N36797);
and and22111(N36803,N36805,N36806);
and and22112(N36804,N36807,N36808);
and and22120(N36814,N36816,N36817);
and and22121(N36815,N36818,N36819);
and and22128(N36829,N36831,N36832);
and and22129(N36830,N36833,N36834);
and and22136(N36844,N36846,N36847);
and and22137(N36845,N36848,N36849);
and and22144(N36859,N36861,N36862);
and and22145(N36860,N36863,N36864);
and and22152(N36874,N36876,N36877);
and and22153(N36875,N36878,N36879);
and and22160(N36889,N36891,N36892);
and and22161(N36890,N36893,N36894);
and and22168(N36903,N36905,N36906);
and and22169(N36904,N36907,N36908);
and and22176(N36917,N36919,N36920);
and and22177(N36918,N36921,N36922);
and and22184(N36931,N36933,N36934);
and and22185(N36932,N36935,N36936);
and and22192(N36945,N36947,N36948);
and and22193(N36946,N36949,N36950);
and and22200(N36959,N36961,N36962);
and and22201(N36960,N36963,N36964);
and and22208(N36973,N36975,N36976);
and and22209(N36974,N36977,N36978);
and and22216(N36987,N36989,N36990);
and and22217(N36988,N36991,N36992);
and and22224(N37001,N37003,N37004);
and and22225(N37002,N37005,N37006);
and and22232(N37015,N37017,N37018);
and and22233(N37016,N37019,N37020);
and and22240(N37029,N37031,N37032);
and and22241(N37030,N37033,N37034);
and and22248(N37043,N37045,N37046);
and and22249(N37044,N37047,N37048);
and and22256(N37056,N37058,N37059);
and and22257(N37057,N37060,N37061);
and and22264(N37069,N37071,N37072);
and and22265(N37070,N37073,N37074);
and and22272(N37082,N37084,N37085);
and and22273(N37083,N37086,N37087);
and and22280(N37095,N37097,N37098);
and and22281(N37096,N37099,N37100);
and and22288(N37108,N37110,N37111);
and and22289(N37109,N37112,N37113);
and and22296(N37120,N37122,N37123);
and and22297(N37121,N37124,N37125);
and and22304(N37132,N37134,N37135);
and and22305(N37133,N37136,N37137);
and and22312(N37144,N37146,N37147);
and and22313(N37145,N37148,N37149);
and and22320(N37156,N37158,N37159);
and and22321(N37157,N37160,N37161);
and and22328(N37168,N37170,N37171);
and and22329(N37169,N37172,N37173);
and and22336(N37180,N37182,N37183);
and and22337(N37181,N37184,N37185);
and and22344(N37191,N37193,N37194);
and and22345(N37192,N37195,N37196);
and and22352(N37202,N37204,N37205);
and and22353(N37203,N37206,N37207);
and and22360(N37213,N37215,N37216);
and and22361(N37214,N37217,N37218);
and and22368(N37223,N37225,N37226);
and and22369(N37224,N37227,N37228);
and and22376(N37233,N37235,N37236);
and and22377(N37234,N37237,N37238);
and and22384(N37243,N37245,N37246);
and and22385(N37244,N37247,N37248);
and and22391(N37254,N37256,N37257);
and and22392(N37255,N37258,N37259);
and and20715(N34585,N34589,N34590);
and and20716(N34586,N34591,N34592);
and and20717(N34587,N34593,N34594);
and and20718(N34588,N34595,R1);
and and20725(N34605,N34609,N34610);
and and20726(N34606,N34611,N34612);
and and20727(N34607,N34613,in2);
and and20728(N34608,N34614,R1);
and and20735(N34623,N34627,N34628);
and and20736(N34624,N34629,N34630);
and and20737(N34625,N34631,N34632);
and and20738(N34626,N34633,N34634);
and and20745(N34640,N34644,N34645);
and and20746(N34641,N34646,N34647);
and and20747(N34642,N34648,N34649);
and and20748(N34643,N34650,N34651);
and and20754(N34658,N34662,N34663);
and and20755(N34659,N34664,N34665);
and and20756(N34660,in2,N34666);
and and20757(N34661,N34667,N34668);
and and20763(N34676,N34680,N34681);
and and20764(N34677,N34682,in1);
and and20765(N34678,N34683,N34684);
and and20766(N34679,N34685,N34686);
and and20772(N34694,N34698,N34699);
and and20773(N34695,N34700,N34701);
and and20774(N34696,N34702,N34703);
and and20775(N34697,N34704,N34705);
and and20781(N34712,N34716,N34717);
and and20782(N34713,N34718,N34719);
and and20783(N34714,N34720,N34721);
and and20784(N34715,N34722,R2);
and and20790(N34730,N34734,N34735);
and and20791(N34731,N34736,N34737);
and and20792(N34732,N34738,R0);
and and20793(N34733,N34739,N34740);
and and20799(N34747,N34751,N34752);
and and20800(N34748,N34753,N34754);
and and20801(N34749,R0,N34755);
and and20802(N34750,N34756,N34757);
and and20808(N34764,N34768,N34769);
and and20809(N34765,N34770,N34771);
and and20810(N34766,in2,R0);
and and20811(N34767,N34772,N34773);
and and20817(N34781,N34785,N34786);
and and20818(N34782,N34787,N34788);
and and20819(N34783,in2,N34789);
and and20820(N34784,N34790,N34791);
and and20826(N34797,N34801,N34802);
and and20827(N34798,N34803,in1);
and and20828(N34799,N34804,R1);
and and20829(N34800,N34805,R3);
and and20835(N34813,N34817,N34818);
and and20836(N34814,N34819,N34820);
and and20837(N34815,in2,N34821);
and and20838(N34816,R2,N34822);
and and20844(N34829,N34833,N34834);
and and20845(N34830,N34835,in1);
and and20846(N34831,N34836,N34837);
and and20847(N34832,R2,N34838);
and and20853(N34845,N34849,N34850);
and and20854(N34846,N34851,N34852);
and and20855(N34847,R0,N34853);
and and20856(N34848,R2,N34854);
and and20862(N34861,N34865,N34866);
and and20863(N34862,N34867,N34868);
and and20864(N34863,in2,N34869);
and and20865(N34864,N34870,R3);
and and20871(N34877,N34881,N34882);
and and20872(N34878,N34883,in1);
and and20873(N34879,N34884,N34885);
and and20874(N34880,N34886,R3);
and and20880(N34893,N34897,N34898);
and and20881(N34894,N34899,in1);
and and20882(N34895,in2,N34900);
and and20883(N34896,N34901,N34902);
and and20889(N34909,N34913,N34914);
and and20890(N34910,N34915,N34916);
and and20891(N34911,R0,N34917);
and and20892(N34912,N34918,R3);
and and20898(N34925,N34929,N34930);
and and20899(N34926,N34931,N34932);
and and20900(N34927,N34933,N34934);
and and20901(N34928,R1,N34935);
and and20907(N34941,N34945,N34946);
and and20908(N34942,N34947,N34948);
and and20909(N34943,N34949,N34950);
and and20910(N34944,R2,N34951);
and and20916(N34957,N34961,N34962);
and and20917(N34958,N34963,in1);
and and20918(N34959,N34964,N34965);
and and20919(N34960,N34966,R3);
and and20925(N34973,N34977,N34978);
and and20926(N34974,N34979,N34980);
and and20927(N34975,in2,R0);
and and20928(N34976,N34981,N34982);
and and20934(N34989,N34993,N34994);
and and20935(N34990,N34995,in1);
and and20936(N34991,R0,N34996);
and and20937(N34992,N34997,N34998);
and and20943(N35005,N35009,N35010);
and and20944(N35006,N35011,N35012);
and and20945(N35007,N35013,N35014);
and and20946(N35008,N35015,R3);
and and20952(N35021,N35025,N35026);
and and20953(N35022,N35027,N35028);
and and20954(N35023,N35029,N35030);
and and20955(N35024,N35031,R3);
and and20961(N35037,N35041,N35042);
and and20962(N35038,N35043,in1);
and and20963(N35039,N35044,N35045);
and and20964(N35040,N35046,N35047);
and and20970(N35053,N35057,N35058);
and and20971(N35054,N35059,N35060);
and and20972(N35055,N35061,N35062);
and and20973(N35056,N35063,R3);
and and20979(N35069,N35073,N35074);
and and20980(N35070,N35075,in2);
and and20981(N35071,R0,N35076);
and and20982(N35072,R2,N35077);
and and20988(N35085,N35089,N35090);
and and20989(N35086,N35091,in1);
and and20990(N35087,in2,N35092);
and and20991(N35088,N35093,R2);
and and20997(N35101,N35105,N35106);
and and20998(N35102,N35107,N35108);
and and20999(N35103,in2,R0);
and and21000(N35104,N35109,N35110);
and and21006(N35117,N35121,N35122);
and and21007(N35118,N35123,N35124);
and and21008(N35119,N35125,N35126);
and and21009(N35120,N35127,R2);
and and21015(N35133,N35137,N35138);
and and21016(N35134,N35139,N35140);
and and21017(N35135,N35141,R1);
and and21018(N35136,R2,N35142);
and and21024(N35149,N35153,N35154);
and and21025(N35150,N35155,in1);
and and21026(N35151,R0,N35156);
and and21027(N35152,R2,R3);
and and21033(N35164,N35168,N35169);
and and21034(N35165,N35170,N35171);
and and21035(N35166,R0,R1);
and and21036(N35167,N35172,N35173);
and and21042(N35179,N35183,N35184);
and and21043(N35180,N35185,N35186);
and and21044(N35181,in2,R0);
and and21045(N35182,R1,N35187);
and and21051(N35194,N35198,N35199);
and and21052(N35195,N35200,N35201);
and and21053(N35196,in2,R0);
and and21054(N35197,N35202,N35203);
and and21060(N35209,N35213,N35214);
and and21061(N35210,N35215,in1);
and and21062(N35211,N35216,R0);
and and21063(N35212,N35217,N35218);
and and21069(N35224,N35228,N35229);
and and21070(N35225,N35230,in1);
and and21071(N35226,N35231,N35232);
and and21072(N35227,R1,N35233);
and and21078(N35239,N35243,N35244);
and and21079(N35240,N35245,N35246);
and and21080(N35241,R0,N35247);
and and21081(N35242,R2,N35248);
and and21087(N35254,N35258,N35259);
and and21088(N35255,N35260,N35261);
and and21089(N35256,N35262,R0);
and and21090(N35257,N35263,R3);
and and21096(N35269,N35273,N35274);
and and21097(N35270,N35275,N35276);
and and21098(N35271,in2,N35277);
and and21099(N35272,R2,N35278);
and and21105(N35284,N35288,N35289);
and and21106(N35285,N35290,in1);
and and21107(N35286,N35291,R0);
and and21108(N35287,R1,N35292);
and and21114(N35299,N35303,N35304);
and and21115(N35300,N35305,in1);
and and21116(N35301,N35306,R0);
and and21117(N35302,N35307,N35308);
and and21123(N35314,N35318,N35319);
and and21124(N35315,N35320,N35321);
and and21125(N35316,N35322,R0);
and and21126(N35317,R1,R2);
and and21132(N35329,N35333,N35334);
and and21133(N35330,N35335,in1);
and and21134(N35331,in2,R0);
and and21135(N35332,N35336,N35337);
and and21141(N35344,N35348,N35349);
and and21142(N35345,N35350,N35351);
and and21143(N35346,N35352,R0);
and and21144(N35347,R2,N35353);
and and21150(N35359,N35363,N35364);
and and21151(N35360,N35365,N35366);
and and21152(N35361,R0,N35367);
and and21153(N35362,N35368,R3);
and and21159(N35374,N35378,N35379);
and and21160(N35375,N35380,in1);
and and21161(N35376,in2,R0);
and and21162(N35377,R1,N35381);
and and21168(N35389,N35393,N35394);
and and21169(N35390,N35395,in1);
and and21170(N35391,N35396,N35397);
and and21171(N35392,R1,N35398);
and and21177(N35404,N35408,N35409);
and and21178(N35405,N35410,N35411);
and and21179(N35406,N35412,N35413);
and and21180(N35407,N35414,R3);
and and21186(N35419,N35423,N35424);
and and21187(N35420,N35425,in1);
and and21188(N35421,N35426,R0);
and and21189(N35422,N35427,N35428);
and and21195(N35434,N35438,N35439);
and and21196(N35435,N35440,in1);
and and21197(N35436,N35441,N35442);
and and21198(N35437,N35443,R3);
and and21204(N35449,N35453,N35454);
and and21205(N35450,N35455,in1);
and and21206(N35451,N35456,N35457);
and and21207(N35452,R1,N35458);
and and21213(N35464,N35468,N35469);
and and21214(N35465,N35470,N35471);
and and21215(N35466,in2,N35472);
and and21216(N35467,R1,N35473);
and and21222(N35479,N35483,N35484);
and and21223(N35480,N35485,in1);
and and21224(N35481,N35486,N35487);
and and21225(N35482,R1,R2);
and and21231(N35494,N35498,N35499);
and and21232(N35495,N35500,N35501);
and and21233(N35496,N35502,R0);
and and21234(N35497,N35503,R2);
and and21240(N35509,N35513,N35514);
and and21241(N35510,N35515,N35516);
and and21242(N35511,R0,N35517);
and and21243(N35512,R2,N35518);
and and21249(N35524,N35528,N35529);
and and21250(N35525,N35530,N35531);
and and21251(N35526,N35532,R0);
and and21252(N35527,R1,N35533);
and and21258(N35539,N35543,N35544);
and and21259(N35540,N35545,N35546);
and and21260(N35541,in2,N35547);
and and21261(N35542,N35548,R2);
and and21267(N35554,N35558,N35559);
and and21268(N35555,N35560,in1);
and and21269(N35556,in2,N35561);
and and21270(N35557,N35562,N35563);
and and21276(N35569,N35573,N35574);
and and21277(N35570,N35575,N35576);
and and21278(N35571,in2,R0);
and and21279(N35572,N35577,R2);
and and21285(N35584,N35588,N35589);
and and21286(N35585,N35590,in1);
and and21287(N35586,N35591,N35592);
and and21288(N35587,R1,R2);
and and21294(N35599,N35603,N35604);
and and21295(N35600,N35605,in2);
and and21296(N35601,N35606,R1);
and and21297(N35602,N35607,R3);
and and21303(N35613,N35617,N35618);
and and21304(N35614,N35619,N35620);
and and21305(N35615,in2,R0);
and and21306(N35616,R1,N35621);
and and21312(N35627,N35631,N35632);
and and21313(N35628,N35633,in1);
and and21314(N35629,in2,R0);
and and21315(N35630,N35634,R2);
and and21321(N35641,N35645,N35646);
and and21322(N35642,N35647,in2);
and and21323(N35643,R0,N35648);
and and21324(N35644,N35649,R3);
and and21330(N35655,N35659,N35660);
and and21331(N35656,N35661,N35662);
and and21332(N35657,R0,R1);
and and21333(N35658,N35663,R3);
and and21339(N35669,N35673,N35674);
and and21340(N35670,N35675,N35676);
and and21341(N35671,N35677,N35678);
and and21342(N35672,R1,R2);
and and21348(N35683,N35687,N35688);
and and21349(N35684,N35689,in1);
and and21350(N35685,in2,N35690);
and and21351(N35686,R1,N35691);
and and21357(N35697,N35701,N35702);
and and21358(N35698,N35703,N35704);
and and21359(N35699,in2,R0);
and and21360(N35700,R1,N35705);
and and21366(N35711,N35715,N35716);
and and21367(N35712,N35717,N35718);
and and21368(N35713,in2,N35719);
and and21369(N35714,R1,R2);
and and21375(N35725,N35729,N35730);
and and21376(N35726,N35731,in1);
and and21377(N35727,N35732,R0);
and and21378(N35728,N35733,R2);
and and21384(N35739,N35743,N35744);
and and21385(N35740,N35745,in1);
and and21386(N35741,N35746,R0);
and and21387(N35742,N35747,R2);
and and21393(N35753,N35757,N35758);
and and21394(N35754,N35759,N35760);
and and21395(N35755,in2,R0);
and and21396(N35756,R2,R3);
and and21402(N35767,N35771,N35772);
and and21403(N35768,N35773,N35774);
and and21404(N35769,N35775,R0);
and and21405(N35770,R1,N35776);
and and21411(N35781,N35785,N35786);
and and21412(N35782,N35787,in1);
and and21413(N35783,in2,N35788);
and and21414(N35784,R1,R3);
and and21420(N35795,N35799,N35800);
and and21421(N35796,N35801,N35802);
and and21422(N35797,in2,N35803);
and and21423(N35798,R1,N35804);
and and21429(N35809,N35813,N35814);
and and21430(N35810,N35815,N35816);
and and21431(N35811,in2,N35817);
and and21432(N35812,R1,R2);
and and21438(N35823,N35827,N35828);
and and21439(N35824,N35829,N35830);
and and21440(N35825,N35831,R0);
and and21441(N35826,N35832,R3);
and and21447(N35837,N35841,N35842);
and and21448(N35838,N35843,in1);
and and21449(N35839,in2,N35844);
and and21450(N35840,N35845,R2);
and and21456(N35851,N35855,N35856);
and and21457(N35852,N35857,in1);
and and21458(N35853,in2,N35858);
and and21459(N35854,R1,R2);
and and21465(N35865,N35869,N35870);
and and21466(N35866,N35871,in1);
and and21467(N35867,N35872,R1);
and and21468(N35868,R2,R3);
and and21474(N35879,N35883,N35884);
and and21475(N35880,N35885,in1);
and and21476(N35881,in2,N35886);
and and21477(N35882,N35887,R3);
and and21483(N35893,N35897,N35898);
and and21484(N35894,N35899,in1);
and and21485(N35895,in2,N35900);
and and21486(N35896,N35901,R3);
and and21492(N35907,N35911,N35912);
and and21493(N35908,in0,N35913);
and and21494(N35909,R0,N35914);
and and21495(N35910,R2,N35915);
and and21501(N35921,N35925,N35926);
and and21502(N35922,in1,N35927);
and and21503(N35923,R0,N35928);
and and21504(N35924,R2,N35929);
and and21510(N35935,N35939,N35940);
and and21511(N35936,N35941,N35942);
and and21512(N35937,in2,R0);
and and21513(N35938,N35943,R2);
and and21519(N35949,N35953,N35954);
and and21520(N35950,in0,N35955);
and and21521(N35951,N35956,R1);
and and21522(N35952,N35957,R3);
and and21528(N35963,N35967,N35968);
and and21529(N35964,in1,N35969);
and and21530(N35965,N35970,R1);
and and21531(N35966,N35971,R3);
and and21537(N35977,N35981,N35982);
and and21538(N35978,N35983,in1);
and and21539(N35979,in2,N35984);
and and21540(N35980,N35985,R2);
and and21546(N35991,N35995,N35996);
and and21547(N35992,N35997,N35998);
and and21548(N35993,N35999,R0);
and and21549(N35994,R1,R2);
and and21555(N36005,N36009,N36010);
and and21556(N36006,N36011,in1);
and and21557(N36007,in2,N36012);
and and21558(N36008,R1,N36013);
and and21564(N36019,N36023,N36024);
and and21565(N36020,N36025,N36026);
and and21566(N36021,N36027,R0);
and and21567(N36022,R1,N36028);
and and21573(N36033,N36037,N36038);
and and21574(N36034,N36039,in1);
and and21575(N36035,in2,R0);
and and21576(N36036,N36040,R3);
and and21582(N36047,N36051,N36052);
and and21583(N36048,N36053,N36054);
and and21584(N36049,N36055,R1);
and and21585(N36050,R2,R3);
and and21591(N36061,N36065,N36066);
and and21592(N36062,N36067,in1);
and and21593(N36063,R0,R1);
and and21594(N36064,N36068,N36069);
and and21600(N36075,N36079,N36080);
and and21601(N36076,N36081,in1);
and and21602(N36077,N36082,N36083);
and and21603(N36078,N36084,R2);
and and21609(N36089,N36093,N36094);
and and21610(N36090,N36095,in1);
and and21611(N36091,in2,N36096);
and and21612(N36092,R1,R2);
and and21618(N36103,N36107,N36108);
and and21619(N36104,N36109,in1);
and and21620(N36105,N36110,R0);
and and21621(N36106,N36111,R3);
and and21627(N36117,N36121,N36122);
and and21628(N36118,N36123,N36124);
and and21629(N36119,N36125,R0);
and and21630(N36120,R1,R3);
and and21636(N36131,N36135,N36136);
and and21637(N36132,N36137,in1);
and and21638(N36133,N36138,R0);
and and21639(N36134,R1,R2);
and and21645(N36145,N36149,N36150);
and and21646(N36146,N36151,N36152);
and and21647(N36147,N36153,R0);
and and21648(N36148,R1,R2);
and and21654(N36159,N36163,N36164);
and and21655(N36160,N36165,in1);
and and21656(N36161,N36166,N36167);
and and21657(N36162,R2,N36168);
and and21663(N36173,N36177,N36178);
and and21664(N36174,N36179,in1);
and and21665(N36175,in2,R0);
and and21666(N36176,N36180,R2);
and and21672(N36187,N36191,N36192);
and and21673(N36188,N36193,N36194);
and and21674(N36189,in2,N36195);
and and21675(N36190,R2,R3);
and and21681(N36200,N36204,N36205);
and and21682(N36201,N36206,in1);
and and21683(N36202,N36207,R1);
and and21684(N36203,R2,R3);
and and21690(N36213,N36217,N36218);
and and21691(N36214,N36219,in1);
and and21692(N36215,N36220,R1);
and and21693(N36216,N36221,R3);
and and21699(N36226,N36230,N36231);
and and21700(N36227,N36232,N36233);
and and21701(N36228,in2,R1);
and and21702(N36229,N36234,R3);
and and21708(N36239,N36243,N36244);
and and21709(N36240,N36245,in1);
and and21710(N36241,N36246,R0);
and and21711(N36242,N36247,R2);
and and21717(N36252,N36256,N36257);
and and21718(N36253,N36258,N36259);
and and21719(N36254,in2,R0);
and and21720(N36255,N36260,R2);
and and21726(N36265,N36269,N36270);
and and21727(N36266,N36271,in1);
and and21728(N36267,N36272,R0);
and and21729(N36268,R1,N36273);
and and21735(N36278,N36282,N36283);
and and21736(N36279,N36284,in1);
and and21737(N36280,N36285,R0);
and and21738(N36281,N36286,R3);
and and21744(N36291,N36295,N36296);
and and21745(N36292,N36297,N36298);
and and21746(N36293,in2,R0);
and and21747(N36294,N36299,R3);
and and21753(N36304,N36308,N36309);
and and21754(N36305,N36310,in1);
and and21755(N36306,in2,R0);
and and21756(N36307,R1,N36311);
and and21762(N36317,N36321,N36322);
and and21763(N36318,N36323,in1);
and and21764(N36319,in2,R0);
and and21765(N36320,R1,R2);
and and21771(N36330,N36334,N36335);
and and21772(N36331,N36336,N36337);
and and21773(N36332,N36338,N36339);
and and21774(N36333,R2,R3);
and and21780(N36343,N36347,N36348);
and and21781(N36344,in0,in2);
and and21782(N36345,R0,N36349);
and and21783(N36346,N36350,R3);
and and21789(N36356,N36360,N36361);
and and21790(N36357,in0,in1);
and and21791(N36358,R0,N36362);
and and21792(N36359,N36363,R3);
and and21798(N36369,N36373,N36374);
and and21799(N36370,N36375,N36376);
and and21800(N36371,in2,R0);
and and21801(N36372,R1,R2);
and and21807(N36382,N36386,N36387);
and and21808(N36383,N36388,in1);
and and21809(N36384,in2,N36389);
and and21810(N36385,R1,R2);
and and21816(N36395,N36399,N36400);
and and21817(N36396,N36401,N36402);
and and21818(N36397,in2,R0);
and and21819(N36398,N36403,R2);
and and21825(N36408,N36412,N36413);
and and21826(N36409,N36414,N36415);
and and21827(N36410,in2,R0);
and and21828(N36411,R1,N36416);
and and21834(N36421,N36425,N36426);
and and21835(N36422,N36427,N36428);
and and21836(N36423,in2,R0);
and and21837(N36424,N36429,R2);
and and21843(N36434,N36438,N36439);
and and21844(N36435,N36440,in1);
and and21845(N36436,N36441,R0);
and and21846(N36437,N36442,R2);
and and21852(N36447,N36451,N36452);
and and21853(N36448,N36453,in1);
and and21854(N36449,in2,R1);
and and21855(N36450,N36454,N36455);
and and21861(N36460,N36464,N36465);
and and21862(N36461,N36466,N36467);
and and21863(N36462,N36468,R0);
and and21864(N36463,R2,R3);
and and21870(N36473,N36477,N36478);
and and21871(N36474,N36479,in1);
and and21872(N36475,N36480,N36481);
and and21873(N36476,R1,N36482);
and and21879(N36486,N36490,N36491);
and and21880(N36487,N36492,in1);
and and21881(N36488,in2,R0);
and and21882(N36489,R2,R3);
and and21888(N36499,N36503,N36504);
and and21889(N36500,N36505,N36506);
and and21890(N36501,in2,R1);
and and21891(N36502,R2,N36507);
and and21897(N36512,N36516,N36517);
and and21898(N36513,N36518,in1);
and and21899(N36514,in2,N36519);
and and21900(N36515,N36520,R2);
and and21906(N36525,N36529,N36530);
and and21907(N36526,N36531,in1);
and and21908(N36527,N36532,R0);
and and21909(N36528,R1,N36533);
and and21915(N36538,N36542,N36543);
and and21916(N36539,N36544,N36545);
and and21917(N36540,in2,N36546);
and and21918(N36541,R1,R2);
and and21924(N36551,N36555,N36556);
and and21925(N36552,N36557,in1);
and and21926(N36553,N36558,R0);
and and21927(N36554,N36559,R2);
and and21933(N36564,N36568,N36569);
and and21934(N36565,N36570,in1);
and and21935(N36566,in2,R0);
and and21936(N36567,N36571,N36572);
and and21942(N36577,N36581,N36582);
and and21943(N36578,N36583,in1);
and and21944(N36579,in2,R0);
and and21945(N36580,R1,N36584);
and and21951(N36590,N36594,N36595);
and and21952(N36591,N36596,in1);
and and21953(N36592,in2,R0);
and and21954(N36593,N36597,N36598);
and and21960(N36603,N36607,N36608);
and and21961(N36604,in0,in2);
and and21962(N36605,R0,N36609);
and and21963(N36606,R2,N36610);
and and21969(N36616,N36620,N36621);
and and21970(N36617,in0,in2);
and and21971(N36618,N36622,R1);
and and21972(N36619,N36623,R3);
and and21978(N36629,N36633,N36634);
and and21979(N36630,N36635,in1);
and and21980(N36631,in2,R1);
and and21981(N36632,N36636,R3);
and and21987(N36642,N36646,N36647);
and and21988(N36643,N36648,N36649);
and and21989(N36644,R0,R1);
and and21990(N36645,N36650,R3);
and and21996(N36654,N36658,N36659);
and and21997(N36655,N36660,in2);
and and21998(N36656,R0,R1);
and and21999(N36657,R2,R3);
and and22005(N36666,N36670,N36671);
and and22006(N36667,N36672,N36673);
and and22007(N36668,in2,R0);
and and22008(N36669,N36674,R2);
and and22014(N36678,N36682,N36683);
and and22015(N36679,N36684,in1);
and and22016(N36680,in2,R0);
and and22017(N36681,R1,N36685);
and and22023(N36690,N36694,N36695);
and and22024(N36691,N36696,in1);
and and22025(N36692,in2,R0);
and and22026(N36693,R1,R2);
and and22032(N36702,N36706,N36707);
and and22033(N36703,N36708,N36709);
and and22034(N36704,in2,N36710);
and and22035(N36705,R1,R3);
and and22041(N36714,N36718,N36719);
and and22042(N36715,N36720,in1);
and and22043(N36716,in2,N36721);
and and22044(N36717,R1,R3);
and and22050(N36726,N36730,N36731);
and and22051(N36727,N36732,in1);
and and22052(N36728,N36733,R1);
and and22053(N36729,R2,R3);
and and22059(N36738,N36742,N36743);
and and22060(N36739,N36744,in1);
and and22061(N36740,N36745,R0);
and and22062(N36741,R2,R3);
and and22068(N36750,N36754,N36755);
and and22069(N36751,N36756,in1);
and and22070(N36752,in2,R1);
and and22071(N36753,R2,N36757);
and and22077(N36761,N36765,N36766);
and and22078(N36762,N36767,in1);
and and22079(N36763,R0,N36768);
and and22080(N36764,R2,R3);
and and22086(N36772,N36776,N36777);
and and22087(N36773,N36778,in1);
and and22088(N36774,R0,R1);
and and22089(N36775,R2,N36779);
and and22095(N36783,N36787,N36788);
and and22096(N36784,N36789,in1);
and and22097(N36785,in2,R0);
and and22098(N36786,R1,R2);
and and22104(N36794,N36798,N36799);
and and22105(N36795,N36800,in1);
and and22106(N36796,in2,R0);
and and22107(N36797,N36801,R2);
and and22113(N36805,N36809,N36810);
and and22114(N36806,N36811,in1);
and and22115(N36807,in2,R0);
and and22116(N36808,R2,R3);
and and22122(N36816,N36820,N36821);
and and22123(N36817,N36822,N36823);
and and22124(N36818,N36824,N36825);
and and22125(N36819,R4,R5);
and and22130(N36831,N36835,N36836);
and and22131(N36832,N36837,N36838);
and and22132(N36833,N36839,R3);
and and22133(N36834,R4,N36840);
and and22138(N36846,N36850,N36851);
and and22139(N36847,N36852,N36853);
and and22140(N36848,R2,N36854);
and and22141(N36849,N36855,N36856);
and and22146(N36861,N36865,N36866);
and and22147(N36862,N36867,N36868);
and and22148(N36863,R2,R3);
and and22149(N36864,N36869,N36870);
and and22154(N36876,N36880,N36881);
and and22155(N36877,N36882,N36883);
and and22156(N36878,R2,N36884);
and and22157(N36879,N36885,N36886);
and and22162(N36891,N36895,N36896);
and and22163(N36892,in1,in2);
and and22164(N36893,N36897,R1);
and and22165(N36894,N36898,N36899);
and and22170(N36905,N36909,N36910);
and and22171(N36906,N36911,N36912);
and and22172(N36907,R2,R3);
and and22173(N36908,R4,N36913);
and and22178(N36919,N36923,N36924);
and and22179(N36920,in1,N36925);
and and22180(N36921,N36926,N36927);
and and22181(N36922,R3,R4);
and and22186(N36933,N36937,N36938);
and and22187(N36934,in1,N36939);
and and22188(N36935,R1,R2);
and and22189(N36936,N36940,N36941);
and and22194(N36947,N36951,in0);
and and22195(N36948,N36952,N36953);
and and22196(N36949,R2,N36954);
and and22197(N36950,N36955,N36956);
and and22202(N36961,N36965,in0);
and and22203(N36962,N36966,R1);
and and22204(N36963,N36967,N36968);
and and22205(N36964,N36969,R5);
and and22210(N36975,N36979,in0);
and and22211(N36976,N36980,N36981);
and and22212(N36977,N36982,R3);
and and22213(N36978,N36983,R5);
and and22218(N36989,N36993,N36994);
and and22219(N36990,in1,in2);
and and22220(N36991,N36995,N36996);
and and22221(N36992,R4,N36997);
and and22226(N37003,N37007,N37008);
and and22227(N37004,N37009,N37010);
and and22228(N37005,R1,N37011);
and and22229(N37006,N37012,R4);
and and22234(N37017,N37021,N37022);
and and22235(N37018,in1,N37023);
and and22236(N37019,N37024,R1);
and and22237(N37020,R2,N37025);
and and22242(N37031,N37035,N37036);
and and22243(N37032,N37037,N37038);
and and22244(N37033,N37039,R2);
and and22245(N37034,R3,R4);
and and22250(N37045,N37049,N37050);
and and22251(N37046,N37051,N37052);
and and22252(N37047,R0,R1);
and and22253(N37048,N37053,R3);
and and22258(N37058,N37062,N37063);
and and22259(N37059,N37064,N37065);
and and22260(N37060,R1,N37066);
and and22261(N37061,R3,R5);
and and22266(N37071,N37075,in0);
and and22267(N37072,R0,N37076);
and and22268(N37073,N37077,N37078);
and and22269(N37074,R4,N37079);
and and22274(N37084,N37088,in0);
and and22275(N37085,R0,N37089);
and and22276(N37086,N37090,N37091);
and and22277(N37087,R4,N37092);
and and22282(N37097,N37101,in0);
and and22283(N37098,R0,N37102);
and and22284(N37099,N37103,R3);
and and22285(N37100,R4,N37104);
and and22290(N37110,N37114,N37115);
and and22291(N37111,in1,N37116);
and and22292(N37112,R1,R2);
and and22293(N37113,R3,R4);
and and22298(N37122,N37126,N37127);
and and22299(N37123,N37128,N37129);
and and22300(N37124,R1,R2);
and and22301(N37125,R3,N37130);
and and22306(N37134,N37138,N37139);
and and22307(N37135,in1,N37140);
and and22308(N37136,R0,R1);
and and22309(N37137,R4,N37141);
and and22314(N37146,N37150,N37151);
and and22315(N37147,in1,in2);
and and22316(N37148,R0,R2);
and and22317(N37149,N37152,N37153);
and and22322(N37158,N37162,N37163);
and and22323(N37159,N37164,R0);
and and22324(N37160,R1,R2);
and and22325(N37161,N37165,R4);
and and22330(N37170,N37174,N37175);
and and22331(N37171,N37176,R0);
and and22332(N37172,R1,R2);
and and22333(N37173,N37177,R4);
and and22338(N37182,N37186,N37187);
and and22339(N37183,in2,N37188);
and and22340(N37184,R1,R2);
and and22341(N37185,R3,R4);
and and22346(N37193,N37197,N37198);
and and22347(N37194,N37199,N37200);
and and22348(N37195,R1,R2);
and and22349(N37196,R3,R4);
and and22354(N37204,N37208,N37209);
and and22355(N37205,in1,N37210);
and and22356(N37206,R1,R2);
and and22357(N37207,R3,R5);
and and22362(N37215,N37219,N37220);
and and22363(N37216,N37221,in2);
and and22364(N37217,R0,R1);
and and22365(N37218,R3,R4);
and and22370(N37225,N37229,in0);
and and22371(N37226,R0,R1);
and and22372(N37227,R2,R3);
and and22373(N37228,N37230,N37231);
and and22378(N37235,N37239,N37240);
and and22379(N37236,in1,in2);
and and22380(N37237,N37241,R1);
and and22381(N37238,R2,R3);
and and22386(N37245,in0,N37249);
and and22387(N37246,R1,N37250);
and and22388(N37247,N37251,N37252);
and and22389(N37248,R6,R7);
and and22393(N37256,in0,N37260);
and and22394(N37257,N37261,R2);
and and22395(N37258,N37262,R5);
and and22396(N37259,N37263,R7);
and and20719(N34589,N34596,N34597);
and and20720(N34590,N34598,N34599);
and and20721(N34591,N34600,N34601);
and and20729(N34609,R2,N34615);
and and20730(N34610,N34616,N34617);
and and20731(N34611,N34618,N34619);
and and20739(N34627,R2,R3);
and and20740(N34628,N34635,R5);
and and20741(N34629,R6,N34636);
and and20749(N34644,N34652,N34653);
and and20750(N34645,N34654,R7);
and and20758(N34662,N34669,N34670);
and and20759(N34663,N34671,N34672);
and and20767(N34680,N34687,N34688);
and and20768(N34681,N34689,N34690);
and and20776(N34698,N34706,N34707);
and and20777(N34699,R6,N34708);
and and20785(N34716,N34723,N34724);
and and20786(N34717,N34725,N34726);
and and20794(N34734,R3,N34741);
and and20795(N34735,N34742,N34743);
and and20803(N34751,N34758,N34759);
and and20804(N34752,N34760,R7);
and and20812(N34768,N34774,N34775);
and and20813(N34769,N34776,N34777);
and and20821(N34785,R4,N34792);
and and20822(N34786,N34793,R7);
and and20830(N34801,N34806,N34807);
and and20831(N34802,N34808,N34809);
and and20839(N34817,N34823,R5);
and and20840(N34818,N34824,N34825);
and and20848(N34833,N34839,R5);
and and20849(N34834,N34840,N34841);
and and20857(N34849,N34855,N34856);
and and20858(N34850,R6,N34857);
and and20866(N34865,N34871,N34872);
and and20867(N34866,N34873,R7);
and and20875(N34881,N34887,N34888);
and and20876(N34882,N34889,R7);
and and20884(N34897,N34903,N34904);
and and20885(N34898,N34905,R7);
and and20893(N34913,N34919,N34920);
and and20894(N34914,R6,N34921);
and and20902(N34929,R3,N34936);
and and20903(N34930,N34937,R6);
and and20911(N34945,R4,R5);
and and20912(N34946,N34952,N34953);
and and20920(N34961,N34967,N34968);
and and20921(N34962,R6,N34969);
and and20929(N34977,N34983,N34984);
and and20930(N34978,R6,N34985);
and and20938(N34993,N34999,N35000);
and and20939(N34994,R6,N35001);
and and20947(N35009,N35016,R5);
and and20948(N35010,N35017,R7);
and and20956(N35025,N35032,N35033);
and and20957(N35026,R6,R7);
and and20965(N35041,R4,N35048);
and and20966(N35042,R6,N35049);
and and20974(N35057,R4,N35064);
and and20975(N35058,R6,N35065);
and and20983(N35073,N35078,N35079);
and and20984(N35074,N35080,N35081);
and and20992(N35089,N35094,N35095);
and and20993(N35090,N35096,N35097);
and and21001(N35105,R4,N35111);
and and21002(N35106,N35112,N35113);
and and21010(N35121,R3,N35128);
and and21011(N35122,N35129,R7);
and and21019(N35137,N35143,R5);
and and21020(N35138,N35144,N35145);
and and21028(N35153,N35157,N35158);
and and21029(N35154,N35159,N35160);
and and21037(N35168,N35174,R5);
and and21038(N35169,R6,N35175);
and and21046(N35183,R3,N35188);
and and21047(N35184,N35189,N35190);
and and21055(N35198,R3,N35204);
and and21056(N35199,R5,N35205);
and and21064(N35213,R3,N35219);
and and21065(N35214,R5,N35220);
and and21073(N35228,R4,R5);
and and21074(N35229,N35234,N35235);
and and21082(N35243,R4,N35249);
and and21083(N35244,R6,N35250);
and and21091(N35258,N35264,R5);
and and21092(N35259,R6,N35265);
and and21100(N35273,R4,N35279);
and and21101(N35274,R6,N35280);
and and21109(N35288,R4,N35293);
and and21110(N35289,N35294,N35295);
and and21118(N35303,R3,N35309);
and and21119(N35304,N35310,R7);
and and21127(N35318,N35323,N35324);
and and21128(N35319,R6,N35325);
and and21136(N35333,R3,N35338);
and and21137(N35334,N35339,N35340);
and and21145(N35348,N35354,N35355);
and and21146(N35349,R6,R7);
and and21154(N35363,N35369,N35370);
and and21155(N35364,R6,R7);
and and21163(N35378,N35382,N35383);
and and21164(N35379,N35384,N35385);
and and21172(N35393,N35399,R5);
and and21173(N35394,R6,N35400);
and and21181(N35408,R4,N35415);
and and21182(N35409,R6,R7);
and and21190(N35423,R3,R4);
and and21191(N35424,N35429,N35430);
and and21199(N35438,N35444,R5);
and and21200(N35439,R6,N35445);
and and21208(N35453,R4,N35459);
and and21209(N35454,R6,N35460);
and and21217(N35468,R4,N35474);
and and21218(N35469,R6,N35475);
and and21226(N35483,N35488,N35489);
and and21227(N35484,N35490,R7);
and and21235(N35498,R4,N35504);
and and21236(N35499,N35505,R7);
and and21244(N35513,R4,R5);
and and21245(N35514,N35519,N35520);
and and21253(N35528,N35534,R4);
and and21254(N35529,R5,N35535);
and and21262(N35543,N35549,R4);
and and21263(N35544,N35550,R7);
and and21271(N35558,R3,R4);
and and21272(N35559,N35564,N35565);
and and21280(N35573,N35578,N35579);
and and21281(N35574,N35580,R7);
and and21289(N35588,N35593,N35594);
and and21290(N35589,R6,N35595);
and and21298(N35603,N35608,N35609);
and and21299(N35604,R6,R7);
and and21307(N35617,N35622,R5);
and and21308(N35618,R6,N35623);
and and21316(N35631,N35635,N35636);
and and21317(N35632,R6,N35637);
and and21325(N35645,R4,N35650);
and and21326(N35646,R6,N35651);
and and21334(N35659,N35664,R5);
and and21335(N35660,N35665,R7);
and and21343(N35673,N35679,R4);
and and21344(N35674,R6,R7);
and and21352(N35687,R3,N35692);
and and21353(N35688,R5,N35693);
and and21361(N35701,N35706,R4);
and and21362(N35702,N35707,R7);
and and21370(N35715,R4,R5);
and and21371(N35716,N35720,N35721);
and and21379(N35729,N35734,R4);
and and21380(N35730,N35735,R6);
and and21388(N35743,R3,N35748);
and and21389(N35744,R6,N35749);
and and21397(N35757,N35761,N35762);
and and21398(N35758,R6,N35763);
and and21406(N35771,R3,R4);
and and21407(N35772,N35777,R7);
and and21415(N35785,N35789,N35790);
and and21416(N35786,R6,N35791);
and and21424(N35799,R3,R5);
and and21425(N35800,R6,N35805);
and and21433(N35813,N35818,R5);
and and21434(N35814,N35819,R7);
and and21442(N35827,R4,R5);
and and21443(N35828,N35833,R7);
and and21451(N35841,R3,N35846);
and and21452(N35842,R5,N35847);
and and21460(N35855,N35859,R4);
and and21461(N35856,N35860,N35861);
and and21469(N35869,N35873,R5);
and and21470(N35870,N35874,N35875);
and and21478(N35883,N35888,R5);
and and21479(N35884,N35889,R7);
and and21487(N35897,N35902,N35903);
and and21488(N35898,R6,R7);
and and21496(N35911,N35916,N35917);
and and21497(N35912,R6,R7);
and and21505(N35925,N35930,N35931);
and and21506(N35926,R6,R7);
and and21514(N35939,N35944,N35945);
and and21515(N35940,R6,R7);
and and21523(N35953,N35958,R5);
and and21524(N35954,N35959,R7);
and and21532(N35967,N35972,R5);
and and21533(N35968,N35973,R7);
and and21541(N35981,N35986,R5);
and and21542(N35982,N35987,R7);
and and21550(N35995,R3,N36000);
and and21551(N35996,R5,N36001);
and and21559(N36009,N36014,R5);
and and21560(N36010,R6,N36015);
and and21568(N36023,R4,N36029);
and and21569(N36024,R6,R7);
and and21577(N36037,R4,N36041);
and and21578(N36038,N36042,N36043);
and and21586(N36051,R4,N36056);
and and21587(N36052,R6,N36057);
and and21595(N36065,N36070,N36071);
and and21596(N36066,R6,R7);
and and21604(N36079,R4,N36085);
and and21605(N36080,R6,R7);
and and21613(N36093,N36097,N36098);
and and21614(N36094,N36099,R6);
and and21622(N36107,R4,R5);
and and21623(N36108,N36112,N36113);
and and21631(N36121,N36126,N36127);
and and21632(N36122,R6,R7);
and and21640(N36135,R3,N36139);
and and21641(N36136,N36140,N36141);
and and21649(N36149,N36154,N36155);
and and21650(N36150,R5,R6);
and and21658(N36163,R4,N36169);
and and21659(N36164,R6,R7);
and and21667(N36177,N36181,R4);
and and21668(N36178,N36182,N36183);
and and21676(N36191,R4,N36196);
and and21677(N36192,R6,R7);
and and21685(N36204,N36208,N36209);
and and21686(N36205,R6,R7);
and and21694(N36217,R4,N36222);
and and21695(N36218,R6,R7);
and and21703(N36230,R4,N36235);
and and21704(N36231,R6,R7);
and and21712(N36243,R3,N36248);
and and21713(N36244,R5,R7);
and and21721(N36256,R3,R4);
and and21722(N36257,N36261,R7);
and and21730(N36269,R4,R5);
and and21731(N36270,N36274,R7);
and and21739(N36282,R4,N36287);
and and21740(N36283,R6,R7);
and and21748(N36295,R4,N36300);
and and21749(N36296,R6,R7);
and and21757(N36308,N36312,R5);
and and21758(N36309,N36313,R7);
and and21766(N36321,N36324,N36325);
and and21767(N36322,R6,N36326);
and and21775(N36334,R4,R5);
and and21776(N36335,R6,R7);
and and21784(N36347,N36351,N36352);
and and21785(N36348,R6,R7);
and and21793(N36360,N36364,N36365);
and and21794(N36361,R6,R7);
and and21802(N36373,N36377,R4);
and and21803(N36374,N36378,R6);
and and21811(N36386,R3,N36390);
and and21812(N36387,N36391,R7);
and and21820(N36399,R3,R4);
and and21821(N36400,R6,N36404);
and and21829(N36412,R3,R4);
and and21830(N36413,N36417,R6);
and and21838(N36425,R4,R5);
and and21839(N36426,R6,N36430);
and and21847(N36438,R4,R5);
and and21848(N36439,R6,N36443);
and and21856(N36451,R4,R5);
and and21857(N36452,N36456,R7);
and and21865(N36464,R4,N36469);
and and21866(N36465,R6,R7);
and and21874(N36477,R3,R4);
and and21875(N36478,R5,R7);
and and21883(N36490,N36493,N36494);
and and21884(N36491,N36495,R7);
and and21892(N36503,R4,R5);
and and21893(N36504,N36508,R7);
and and21901(N36516,R3,R4);
and and21902(N36517,R6,N36521);
and and21910(N36529,R3,N36534);
and and21911(N36530,R6,R7);
and and21919(N36542,R3,N36547);
and and21920(N36543,R5,R6);
and and21928(N36555,R3,R4);
and and21929(N36556,R5,N36560);
and and21937(N36568,R3,R4);
and and21938(N36569,N36573,R7);
and and21946(N36581,R3,R4);
and and21947(N36582,N36585,N36586);
and and21955(N36594,R3,R4);
and and21956(N36595,R6,N36599);
and and21964(N36607,N36611,N36612);
and and21965(N36608,R6,R7);
and and21973(N36620,N36624,R5);
and and21974(N36621,N36625,R7);
and and21982(N36633,N36637,N36638);
and and21983(N36634,R6,R7);
and and21991(N36646,R4,R5);
and and21992(N36647,R6,R7);
and and22000(N36658,N36661,R5);
and and22001(N36659,N36662,R7);
and and22009(N36670,R3,R5);
and and22010(N36671,R6,R7);
and and22018(N36682,R4,N36686);
and and22019(N36683,R6,R7);
and and22027(N36694,N36697,R4);
and and22028(N36695,N36698,R7);
and and22036(N36706,R4,R5);
and and22037(N36707,R6,R7);
and and22045(N36718,R4,R5);
and and22046(N36719,N36722,R7);
and and22054(N36730,R4,N36734);
and and22055(N36731,R6,R7);
and and22063(N36742,R4,R5);
and and22064(N36743,R6,N36746);
and and22072(N36754,R4,R5);
and and22073(N36755,R6,R7);
and and22081(N36765,R4,R5);
and and22082(N36766,R6,R7);
and and22090(N36776,R4,R5);
and and22091(N36777,R6,R7);
and and22099(N36787,N36790,R5);
and and22100(N36788,R6,R7);
and and22108(N36798,R3,R4);
and and22109(N36799,R6,R7);
and and22117(N36809,R4,R5);
and and22118(N36810,N36812,R7);
and and22126(N36820,N36826,N36827);
and and22134(N36835,N36841,N36842);
and and22142(N36850,N36857,R7);
and and22150(N36865,N36871,N36872);
and and22158(N36880,N36887,R7);
and and22166(N36895,N36900,N36901);
and and22174(N36909,N36914,N36915);
and and22182(N36923,N36928,N36929);
and and22190(N36937,N36942,N36943);
and and22198(N36951,R6,N36957);
and and22206(N36965,N36970,N36971);
and and22214(N36979,N36984,N36985);
and and22222(N36993,N36998,N36999);
and and22230(N37007,N37013,R7);
and and22238(N37021,N37026,N37027);
and and22246(N37035,N37040,N37041);
and and22254(N37049,R6,N37054);
and and22262(N37062,R6,N37067);
and and22270(N37075,N37080,R7);
and and22278(N37088,R6,N37093);
and and22286(N37101,N37105,N37106);
and and22294(N37114,N37117,N37118);
and and22302(N37126,R5,R7);
and and22310(N37138,N37142,R7);
and and22318(N37150,N37154,R7);
and and22326(N37162,R5,N37166);
and and22334(N37174,R5,N37178);
and and22342(N37186,N37189,R7);
and and22350(N37197,R5,R7);
and and22358(N37208,R6,N37211);
and and22366(N37219,R5,R7);
and and22374(N37229,R6,R7);
and and22382(N37239,R5,R6);
and and22397(N37322,N37323,N37324);
and and22404(N37332,N37333,N37334);
and and22410(N37344,N37345,N37346);
and and22416(N37356,N37357,N37358);
and and22422(N37368,N37369,N37370);
and and22428(N37380,N37381,N37382);
and and22434(N37392,N37393,N37394);
and and22440(N37404,N37405,N37406);
and and22446(N37415,N37416,N37417);
and and22452(N37426,N37427,N37428);
and and22458(N37437,N37438,N37439);
and and22464(N37448,N37449,N37450);
and and22470(N37459,N37460,N37461);
and and22476(N37470,N37471,N37472);
and and22482(N37481,N37482,N37483);
and and22488(N37492,N37493,N37494);
and and22494(N37503,N37504,N37505);
and and22500(N37514,N37515,N37516);
and and22506(N37525,N37526,N37527);
and and22512(N37536,N37537,N37538);
and and22518(N37546,N37547,N37548);
and and22524(N37556,N37557,N37558);
and and22530(N37566,N37567,N37568);
and and22536(N37576,N37577,N37578);
and and22542(N37586,N37587,N37588);
and and22548(N37596,N37597,N37598);
and and22554(N37606,N37607,N37608);
and and22560(N37616,N37617,N37618);
and and22566(N37626,N37627,N37628);
and and22572(N37636,N37637,N37638);
and and22578(N37645,N37646,N37647);
and and22584(N37654,N37655,N37656);
and and22590(N37663,N37664,N37665);
and and22596(N37672,N37673,N37674);
and and22602(N37681,N37682,N37683);
and and22608(N37690,N37691,N37692);
and and22614(N37699,N37700,N37701);
and and22620(N37708,N37709,N37710);
and and22626(N37717,N37718,N37719);
and and22632(N37726,N37727,N37728);
and and22638(N37735,N37736,N37737);
and and22644(N37744,N37745,N37746);
and and22650(N37753,N37754,N37755);
and and22656(N37762,N37763,N37764);
and and22662(N37770,N37771,N37772);
and and22668(N37778,N37779,N37780);
and and22674(N37786,N37787,N37788);
and and22680(N37794,N37795,N37796);
and and22686(N37802,N37803,N37804);
and and22692(N37810,N37811,N37812);
and and22698(N37818,N37819,N37820);
and and22704(N37825,N37826,N37827);
and and22710(N37832,N37833,N37834);
and and22716(N37839,N37840,N37841);
and and22722(N37846,N37847,N37848);
and and22728(N37853,N37854,N37855);
and and22734(N37860,N37861,N37862);
and and22740(N37867,N37868,N37869);
and and22745(N37876,N37877,N37878);
and and22398(N37323,N37325,N37326);
and and22399(N37324,N37327,N37328);
and and22405(N37333,N37335,N37336);
and and22406(N37334,N37337,N37338);
and and22411(N37345,N37347,N37348);
and and22412(N37346,N37349,N37350);
and and22417(N37357,N37359,N37360);
and and22418(N37358,N37361,N37362);
and and22423(N37369,N37371,N37372);
and and22424(N37370,N37373,N37374);
and and22429(N37381,N37383,N37384);
and and22430(N37382,N37385,N37386);
and and22435(N37393,N37395,N37396);
and and22436(N37394,N37397,N37398);
and and22441(N37405,N37407,N37408);
and and22442(N37406,N37409,R0);
and and22447(N37416,N37418,N37419);
and and22448(N37417,N37420,N37421);
and and22453(N37427,N37429,N37430);
and and22454(N37428,N37431,N37432);
and and22459(N37438,N37440,N37441);
and and22460(N37439,N37442,R0);
and and22465(N37449,N37451,N37452);
and and22466(N37450,N37453,N37454);
and and22471(N37460,N37462,N37463);
and and22472(N37461,N37464,N37465);
and and22477(N37471,N37473,N37474);
and and22478(N37472,N37475,N37476);
and and22483(N37482,N37484,N37485);
and and22484(N37483,N37486,N37487);
and and22489(N37493,N37495,N37496);
and and22490(N37494,N37497,R0);
and and22495(N37504,N37506,N37507);
and and22496(N37505,N37508,N37509);
and and22501(N37515,N37517,N37518);
and and22502(N37516,N37519,N37520);
and and22507(N37526,N37528,N37529);
and and22508(N37527,N37530,N37531);
and and22513(N37537,N37539,N37540);
and and22514(N37538,N37541,N37542);
and and22519(N37547,N37549,N37550);
and and22520(N37548,N37551,N37552);
and and22525(N37557,N37559,N37560);
and and22526(N37558,N37561,R0);
and and22531(N37567,N37569,N37570);
and and22532(N37568,N37571,N37572);
and and22537(N37577,N37579,N37580);
and and22538(N37578,N37581,N37582);
and and22543(N37587,N37589,N37590);
and and22544(N37588,N37591,N37592);
and and22549(N37597,N37599,N37600);
and and22550(N37598,N37601,N37602);
and and22555(N37607,N37609,N37610);
and and22556(N37608,N37611,N37612);
and and22561(N37617,N37619,N37620);
and and22562(N37618,N37621,N37622);
and and22567(N37627,N37629,N37630);
and and22568(N37628,N37631,N37632);
and and22573(N37637,N37639,N37640);
and and22574(N37638,N37641,R0);
and and22579(N37646,N37648,N37649);
and and22580(N37647,N37650,R0);
and and22585(N37655,N37657,N37658);
and and22586(N37656,N37659,R0);
and and22591(N37664,N37666,N37667);
and and22592(N37665,N37668,R0);
and and22597(N37673,N37675,N37676);
and and22598(N37674,N37677,R0);
and and22603(N37682,N37684,N37685);
and and22604(N37683,N37686,N37687);
and and22609(N37691,N37693,N37694);
and and22610(N37692,N37695,R0);
and and22615(N37700,N37702,N37703);
and and22616(N37701,N37704,R0);
and and22621(N37709,N37711,N37712);
and and22622(N37710,N37713,R0);
and and22627(N37718,N37720,N37721);
and and22628(N37719,N37722,R0);
and and22633(N37727,N37729,N37730);
and and22634(N37728,N37731,R0);
and and22639(N37736,N37738,N37739);
and and22640(N37737,N37740,N37741);
and and22645(N37745,N37747,N37748);
and and22646(N37746,N37749,N37750);
and and22651(N37754,N37756,N37757);
and and22652(N37755,N37758,R0);
and and22657(N37763,N37765,N37766);
and and22658(N37764,N37767,R0);
and and22663(N37771,N37773,N37774);
and and22664(N37772,N37775,N37776);
and and22669(N37779,N37781,N37782);
and and22670(N37780,N37783,R0);
and and22675(N37787,N37789,N37790);
and and22676(N37788,N37791,R0);
and and22681(N37795,N37797,N37798);
and and22682(N37796,N37799,N37800);
and and22687(N37803,N37805,N37806);
and and22688(N37804,N37807,R0);
and and22693(N37811,N37813,N37814);
and and22694(N37812,N37815,N37816);
and and22699(N37819,N37821,N37822);
and and22700(N37820,N37823,R0);
and and22705(N37826,N37828,N37829);
and and22706(N37827,N37830,R1);
and and22711(N37833,N37835,N37836);
and and22712(N37834,N37837,R0);
and and22717(N37840,N37842,N37843);
and and22718(N37841,N37844,R0);
and and22723(N37847,N37849,N37850);
and and22724(N37848,N37851,R0);
and and22729(N37854,N37856,N37857);
and and22730(N37855,N37858,R1);
and and22735(N37861,N37863,N37864);
and and22736(N37862,N37865,R0);
and and22741(N37868,N37870,N37871);
and and22742(N37869,R0,N37872);
and and22746(N37877,N37879,N37880);
and and22747(N37878,R1,N37881);
and and22400(N37325,R0,N37329);
and and22401(N37326,R2,N37330);
and and22402(N37327,R4,R5);
and and22403(N37328,R6,N37331);
and and22407(N37335,R1,N37339);
and and22408(N37336,N37340,N37341);
and and22409(N37337,N37342,N37343);
and and22413(N37347,N37351,N37352);
and and22414(N37348,N37353,N37354);
and and22415(N37349,N37355,R7);
and and22419(N37359,N37363,N37364);
and and22420(N37360,N37365,N37366);
and and22421(N37361,R6,N37367);
and and22425(N37371,N37375,N37376);
and and22426(N37372,N37377,R4);
and and22427(N37373,N37378,N37379);
and and22431(N37383,N37387,R2);
and and22432(N37384,N37388,N37389);
and and22433(N37385,N37390,N37391);
and and22437(N37395,N37399,N37400);
and and22438(N37396,N37401,N37402);
and and22439(N37397,N37403,R7);
and and22443(N37407,N37410,N37411);
and and22444(N37408,N37412,R5);
and and22445(N37409,N37413,N37414);
and and22449(N37418,N37422,N37423);
and and22450(N37419,R3,N37424);
and and22451(N37420,N37425,R7);
and and22455(N37429,R2,R3);
and and22456(N37430,N37433,N37434);
and and22457(N37431,N37435,N37436);
and and22461(N37440,N37443,N37444);
and and22462(N37441,N37445,N37446);
and and22463(N37442,R6,N37447);
and and22467(N37451,N37455,R2);
and and22468(N37452,N37456,N37457);
and and22469(N37453,R6,N37458);
and and22473(N37462,R1,N37466);
and and22474(N37463,N37467,N37468);
and and22475(N37464,R5,N37469);
and and22479(N37473,N37477,N37478);
and and22480(N37474,R3,N37479);
and and22481(N37475,R5,N37480);
and and22485(N37484,R1,N37488);
and and22486(N37485,R4,N37489);
and and22487(N37486,N37490,N37491);
and and22491(N37495,N37498,N37499);
and and22492(N37496,N37500,N37501);
and and22493(N37497,N37502,R7);
and and22497(N37506,N37510,R2);
and and22498(N37507,R3,N37511);
and and22499(N37508,N37512,N37513);
and and22503(N37517,N37521,R2);
and and22504(N37518,N37522,R5);
and and22505(N37519,N37523,N37524);
and and22509(N37528,N37532,N37533);
and and22510(N37529,R4,R5);
and and22511(N37530,N37534,N37535);
and and22515(N37539,R1,R2);
and and22516(N37540,R3,N37543);
and and22517(N37541,N37544,N37545);
and and22521(N37549,N37553,R2);
and and22522(N37550,R3,N37554);
and and22523(N37551,N37555,R6);
and and22527(N37559,R1,N37562);
and and22528(N37560,R4,N37563);
and and22529(N37561,N37564,N37565);
and and22533(N37569,R1,N37573);
and and22534(N37570,N37574,N37575);
and and22535(N37571,R6,R7);
and and22539(N37579,N37583,N37584);
and and22540(N37580,R3,N37585);
and and22541(N37581,R6,R7);
and and22545(N37589,N37593,R3);
and and22546(N37590,R4,N37594);
and and22547(N37591,N37595,R7);
and and22551(N37599,R1,N37603);
and and22552(N37600,N37604,R4);
and and22553(N37601,N37605,R7);
and and22557(N37609,R1,R2);
and and22558(N37610,N37613,N37614);
and and22559(N37611,N37615,R6);
and and22563(N37619,R1,N37623);
and and22564(N37620,N37624,R4);
and and22565(N37621,R6,N37625);
and and22569(N37629,R1,N37633);
and and22570(N37630,N37634,R5);
and and22571(N37631,R6,N37635);
and and22575(N37639,R1,N37642);
and and22576(N37640,N37643,R5);
and and22577(N37641,R6,N37644);
and and22581(N37648,N37651,R3);
and and22582(N37649,N37652,R5);
and and22583(N37650,N37653,R7);
and and22587(N37657,N37660,R3);
and and22588(N37658,N37661,R5);
and and22589(N37659,R6,N37662);
and and22593(N37666,R1,N37669);
and and22594(N37667,N37670,R5);
and and22595(N37668,N37671,R7);
and and22599(N37675,R1,R2);
and and22600(N37676,N37678,N37679);
and and22601(N37677,R6,N37680);
and and22605(N37684,N37688,R2);
and and22606(N37685,R3,R5);
and and22607(N37686,N37689,R7);
and and22611(N37693,R2,N37696);
and and22612(N37694,N37697,R5);
and and22613(N37695,N37698,R7);
and and22617(N37702,N37705,R2);
and and22618(N37703,N37706,N37707);
and and22619(N37704,R6,R7);
and and22623(N37711,N37714,R2);
and and22624(N37712,R3,N37715);
and and22625(N37713,R5,N37716);
and and22629(N37720,R1,N37723);
and and22630(N37721,N37724,R4);
and and22631(N37722,N37725,R6);
and and22635(N37729,R1,N37732);
and and22636(N37730,N37733,N37734);
and and22637(N37731,R6,R7);
and and22641(N37738,R1,N37742);
and and22642(N37739,R4,R5);
and and22643(N37740,N37743,R7);
and and22647(N37747,R2,N37751);
and and22648(N37748,R4,N37752);
and and22649(N37749,R6,R7);
and and22653(N37756,R1,R2);
and and22654(N37757,R4,N37759);
and and22655(N37758,N37760,N37761);
and and22659(N37765,N37768,R2);
and and22660(N37766,R3,R4);
and and22661(N37767,N37769,R7);
and and22665(N37773,N37777,R2);
and and22666(N37774,R3,R4);
and and22667(N37775,R5,R6);
and and22671(N37781,R1,N37784);
and and22672(N37782,R3,R4);
and and22673(N37783,R5,N37785);
and and22677(N37789,R1,R2);
and and22678(N37790,R3,N37792);
and and22679(N37791,N37793,R7);
and and22683(N37797,R1,R2);
and and22684(N37798,R3,R4);
and and22685(N37799,R5,N37801);
and and22689(N37805,N37808,R2);
and and22690(N37806,R3,R4);
and and22691(N37807,N37809,R6);
and and22695(N37813,R1,R3);
and and22696(N37814,N37817,R5);
and and22697(N37815,R6,R7);
and and22701(N37821,R1,R2);
and and22702(N37822,N37824,R4);
and and22703(N37823,R5,R7);
and and22707(N37828,R2,N37831);
and and22708(N37829,R4,R5);
and and22709(N37830,R6,R7);
and and22713(N37835,N37838,R2);
and and22714(N37836,R3,R5);
and and22715(N37837,R6,R7);
and and22719(N37842,R1,R2);
and and22720(N37843,N37845,R5);
and and22721(N37844,R6,R7);
and and22725(N37849,R1,R2);
and and22726(N37850,R3,N37852);
and and22727(N37851,R6,R7);
and and22731(N37856,R2,R3);
and and22732(N37857,R4,R5);
and and22733(N37858,R6,N37859);
and and22737(N37863,R1,R3);
and and22738(N37864,R4,R5);
and and22739(N37865,N37866,R7);
and and22743(N37870,R3,N37873);
and and22744(N37871,N37874,N37875);
and and22748(N37879,R3,R5);
and and22749(N37880,R6,R7);
and and22750(N37913,N37914,N37915);
and and22757(N37928,N37929,N37930);
and and22763(N37939,N37940,N37941);
and and22769(N37950,N37951,N37952);
and and22775(N37961,N37962,N37963);
and and22781(N37972,N37973,N37974);
and and22787(N37983,N37984,N37985);
and and22793(N37993,N37994,N37995);
and and22799(N38003,N38004,N38005);
and and22805(N38013,N38014,N38015);
and and22811(N38023,N38024,N38025);
and and22817(N38033,N38034,N38035);
and and22823(N38043,N38044,N38045);
and and22829(N38052,N38053,N38054);
and and22835(N38061,N38062,N38063);
and and22841(N38070,N38071,N38072);
and and22847(N38079,N38080,N38081);
and and22853(N38088,N38089,N38090);
and and22859(N38097,N38098,N38099);
and and22865(N38106,N38107,N38108);
and and22871(N38115,N38116,N38117);
and and22877(N38124,N38125,N38126);
and and22883(N38133,N38134,N38135);
and and22889(N38141,N38142,N38143);
and and22895(N38149,N38150,N38151);
and and22901(N38157,N38158,N38159);
and and22907(N38165,N38166,N38167);
and and22913(N38173,N38174,N38175);
and and22919(N38181,N38182,N38183);
and and22925(N38189,N38190,N38191);
and and22931(N38197,N38198,N38199);
and and22937(N38205,N38206,N38207);
and and22751(N37914,N37916,N37917);
and and22752(N37915,N37918,N37919);
and and22758(N37929,N37931,N37932);
and and22759(N37930,N37933,N37934);
and and22764(N37940,N37942,N37943);
and and22765(N37941,N37944,N37945);
and and22770(N37951,N37953,N37954);
and and22771(N37952,N37955,N37956);
and and22776(N37962,N37964,N37965);
and and22777(N37963,N37966,N37967);
and and22782(N37973,N37975,N37976);
and and22783(N37974,N37977,R0);
and and22788(N37984,N37986,N37987);
and and22789(N37985,N37988,R1);
and and22794(N37994,N37996,N37997);
and and22795(N37995,N37998,R0);
and and22800(N38004,N38006,N38007);
and and22801(N38005,N38008,R0);
and and22806(N38014,N38016,N38017);
and and22807(N38015,N38018,N38019);
and and22812(N38024,N38026,N38027);
and and22813(N38025,N38028,N38029);
and and22818(N38034,N38036,N38037);
and and22819(N38035,N38038,N38039);
and and22824(N38044,N38046,N38047);
and and22825(N38045,N38048,R0);
and and22830(N38053,N38055,N38056);
and and22831(N38054,N38057,N38058);
and and22836(N38062,N38064,N38065);
and and22837(N38063,N38066,R0);
and and22842(N38071,N38073,N38074);
and and22843(N38072,N38075,R0);
and and22848(N38080,N38082,N38083);
and and22849(N38081,N38084,R0);
and and22854(N38089,N38091,N38092);
and and22855(N38090,N38093,N38094);
and and22860(N38098,N38100,N38101);
and and22861(N38099,N38102,R0);
and and22866(N38107,N38109,N38110);
and and22867(N38108,N38111,R1);
and and22872(N38116,N38118,N38119);
and and22873(N38117,N38120,R0);
and and22878(N38125,N38127,N38128);
and and22879(N38126,N38129,N38130);
and and22884(N38134,N38136,N38137);
and and22885(N38135,N38138,N38139);
and and22890(N38142,N38144,N38145);
and and22891(N38143,N38146,R1);
and and22896(N38150,N38152,N38153);
and and22897(N38151,N38154,R0);
and and22902(N38158,N38160,N38161);
and and22903(N38159,N38162,R0);
and and22908(N38166,N38168,N38169);
and and22909(N38167,N38170,R0);
and and22914(N38174,N38176,N38177);
and and22915(N38175,N38178,R0);
and and22920(N38182,N38184,N38185);
and and22921(N38183,N38186,N38187);
and and22926(N38190,N38192,N38193);
and and22927(N38191,N38194,R0);
and and22932(N38198,N38200,N38201);
and and22933(N38199,N38202,R0);
and and22938(N38206,N38208,N38209);
and and22939(N38207,N38210,R1);
and and22753(N37916,N37920,N37921);
and and22754(N37917,N37922,N37923);
and and22755(N37918,N37924,N37925);
and and22756(N37919,N37926,N37927);
and and22760(N37931,R1,N37935);
and and22761(N37932,R3,N37936);
and and22762(N37933,N37937,N37938);
and and22766(N37942,N37946,N37947);
and and22767(N37943,R3,R4);
and and22768(N37944,N37948,N37949);
and and22772(N37953,R2,N37957);
and and22773(N37954,R4,N37958);
and and22774(N37955,N37959,N37960);
and and22778(N37964,N37968,R3);
and and22779(N37965,N37969,N37970);
and and22780(N37966,R6,N37971);
and and22784(N37975,N37978,N37979);
and and22785(N37976,R4,N37980);
and and22786(N37977,N37981,N37982);
and and22790(N37986,N37989,R3);
and and22791(N37987,N37990,N37991);
and and22792(N37988,N37992,R7);
and and22796(N37996,R1,N37999);
and and22797(N37997,N38000,R5);
and and22798(N37998,N38001,N38002);
and and22802(N38006,N38009,N38010);
and and22803(N38007,R3,N38011);
and and22804(N38008,N38012,R7);
and and22808(N38016,N38020,R2);
and and22809(N38017,R3,N38021);
and and22810(N38018,R5,N38022);
and and22814(N38026,R2,N38030);
and and22815(N38027,R4,N38031);
and and22816(N38028,N38032,R7);
and and22820(N38036,N38040,R2);
and and22821(N38037,R4,N38041);
and and22822(N38038,N38042,R7);
and and22826(N38046,R1,R2);
and and22827(N38047,R3,N38049);
and and22828(N38048,N38050,N38051);
and and22832(N38055,R1,N38059);
and and22833(N38056,R3,R4);
and and22834(N38057,R5,N38060);
and and22838(N38064,R1,N38067);
and and22839(N38065,N38068,R4);
and and22840(N38066,N38069,R7);
and and22844(N38073,N38076,R2);
and and22845(N38074,R3,N38077);
and and22846(N38075,N38078,R6);
and and22850(N38082,R1,N38085);
and and22851(N38083,R3,N38086);
and and22852(N38084,R6,N38087);
and and22856(N38091,R1,N38095);
and and22857(N38092,R3,R5);
and and22858(N38093,R6,N38096);
and and22862(N38100,N38103,R2);
and and22863(N38101,N38104,R4);
and and22864(N38102,N38105,R7);
and and22868(N38109,R2,N38112);
and and22869(N38110,R4,N38113);
and and22870(N38111,R6,N38114);
and and22874(N38118,N38121,R2);
and and22875(N38119,R4,R5);
and and22876(N38120,N38122,N38123);
and and22880(N38127,R2,R3);
and and22881(N38128,R4,N38131);
and and22882(N38129,R6,N38132);
and and22886(N38136,R1,R2);
and and22887(N38137,R3,N38140);
and and22888(N38138,R6,R7);
and and22892(N38144,N38147,R3);
and and22893(N38145,R4,N38148);
and and22894(N38146,R6,R7);
and and22898(N38152,N38155,R3);
and and22899(N38153,R4,R5);
and and22900(N38154,R6,N38156);
and and22904(N38160,N38163,R3);
and and22905(N38161,R4,R5);
and and22906(N38162,N38164,R7);
and and22910(N38168,N38171,R3);
and and22911(N38169,R4,N38172);
and and22912(N38170,R6,R7);
and and22916(N38176,R1,R2);
and and22917(N38177,N38179,R4);
and and22918(N38178,N38180,R7);
and and22922(N38184,R1,R2);
and and22923(N38185,R4,R5);
and and22924(N38186,N38188,R7);
and and22928(N38192,R1,R2);
and and22929(N38193,N38195,R4);
and and22930(N38194,R6,N38196);
and and22934(N38200,R1,R2);
and and22935(N38201,R3,R5);
and and22936(N38202,N38203,N38204);
and and22940(N38208,R2,N38211);
and and22941(N38209,R5,N38212);
and and22942(N38225,N38226,N38227);
and and22949(N38237,N38238,N38239);
and and22956(N38249,N38250,N38251);
and and22963(N38260,N38261,N38262);
and and22970(N38271,N38272,N38273);
and and22977(N38282,N38283,N38284);
and and22984(N38293,N38294,N38295);
and and22991(N38304,N38305,N38306);
and and22998(N38314,N38315,N38316);
and and23005(N38323,N38324,N38325);
and and23012(N38332,N38333,N38334);
and and23018(N38343,N38344,N38345);
and and23024(N38354,N38355,N38356);
and and22943(N38226,N38228,N38229);
and and22944(N38227,N38230,N38231);
and and22950(N38238,N38240,N38241);
and and22951(N38239,N38242,N38243);
and and22957(N38250,N38252,N38253);
and and22958(N38251,N38254,N38255);
and and22964(N38261,N38263,N38264);
and and22965(N38262,N38265,N38266);
and and22971(N38272,N38274,N38275);
and and22972(N38273,N38276,N38277);
and and22978(N38283,N38285,N38286);
and and22979(N38284,N38287,N38288);
and and22985(N38294,N38296,N38297);
and and22986(N38295,N38298,N38299);
and and22992(N38305,N38307,N38308);
and and22993(N38306,N38309,N38310);
and and22999(N38315,N38317,N38318);
and and23000(N38316,N38319,N38320);
and and23006(N38324,N38326,N38327);
and and23007(N38325,N38328,N38329);
and and23013(N38333,N38335,N38336);
and and23014(N38334,N38337,R0);
and and23019(N38344,N38346,N38347);
and and23020(N38345,N38348,N38349);
and and23025(N38355,N38357,N38358);
and and23026(N38356,N38359,N38360);
and and22945(N38228,N38232,R1);
and and22946(N38229,R2,N38233);
and and22947(N38230,R4,N38234);
and and22948(N38231,N38235,N38236);
and and22952(N38240,R0,N38244);
and and22953(N38241,N38245,N38246);
and and22954(N38242,R4,N38247);
and and22955(N38243,N38248,R7);
and and22959(N38252,N38256,R1);
and and22960(N38253,R2,R3);
and and22961(N38254,N38257,N38258);
and and22962(N38255,R6,N38259);
and and22966(N38263,N38267,R1);
and and22967(N38264,R2,R3);
and and22968(N38265,N38268,R5);
and and22969(N38266,N38269,N38270);
and and22973(N38274,R0,N38278);
and and22974(N38275,N38279,R3);
and and22975(N38276,N38280,N38281);
and and22976(N38277,R6,R7);
and and22980(N38285,N38289,N38290);
and and22981(N38286,R2,R3);
and and22982(N38287,R4,R5);
and and22983(N38288,N38291,N38292);
and and22987(N38296,N38300,R1);
and and22988(N38297,N38301,R3);
and and22989(N38298,N38302,R5);
and and22990(N38299,N38303,R7);
and and22994(N38307,R0,R1);
and and22995(N38308,N38311,N38312);
and and22996(N38309,R4,R5);
and and22997(N38310,R6,N38313);
and and23001(N38317,R0,R1);
and and23002(N38318,R2,R3);
and and23003(N38319,R4,N38321);
and and23004(N38320,N38322,R7);
and and23008(N38326,R0,R1);
and and23009(N38327,R2,R3);
and and23010(N38328,N38330,R5);
and and23011(N38329,R6,N38331);
and and23015(N38335,R1,N38338);
and and23016(N38336,N38339,N38340);
and and23017(N38337,N38341,N38342);
and and23021(N38346,N38350,N38351);
and and23022(N38347,R4,N38352);
and and23023(N38348,R6,N38353);
and and23027(N38357,N38361,R2);
and and23028(N38358,N38362,R5);
and and23029(N38359,N38363,R7);
and and23030(N38403,N38404,N38405);
and and23037(N38418,N38419,N38420);
and and23043(N38429,N38430,N38431);
and and23049(N38440,N38441,N38442);
and and23055(N38451,N38452,N38453);
and and23061(N38462,N38463,N38464);
and and23067(N38472,N38473,N38474);
and and23073(N38482,N38483,N38484);
and and23079(N38492,N38493,N38494);
and and23085(N38502,N38503,N38504);
and and23091(N38512,N38513,N38514);
and and23097(N38522,N38523,N38524);
and and23103(N38532,N38533,N38534);
and and23109(N38541,N38542,N38543);
and and23115(N38550,N38551,N38552);
and and23121(N38559,N38560,N38561);
and and23127(N38568,N38569,N38570);
and and23133(N38577,N38578,N38579);
and and23139(N38586,N38587,N38588);
and and23145(N38595,N38596,N38597);
and and23151(N38604,N38605,N38606);
and and23157(N38613,N38614,N38615);
and and23163(N38622,N38623,N38624);
and and23169(N38631,N38632,N38633);
and and23175(N38640,N38641,N38642);
and and23181(N38649,N38650,N38651);
and and23187(N38657,N38658,N38659);
and and23193(N38665,N38666,N38667);
and and23199(N38673,N38674,N38675);
and and23205(N38681,N38682,N38683);
and and23211(N38689,N38690,N38691);
and and23217(N38697,N38698,N38699);
and and23223(N38705,N38706,N38707);
and and23229(N38713,N38714,N38715);
and and23235(N38721,N38722,N38723);
and and23241(N38729,N38730,N38731);
and and23247(N38737,N38738,N38739);
and and23252(N38746,N38747,N38748);
and and23257(N38755,N38756,N38757);
and and23262(N38764,N38765,N38766);
and and23031(N38404,N38406,N38407);
and and23032(N38405,N38408,N38409);
and and23038(N38419,N38421,N38422);
and and23039(N38420,N38423,N38424);
and and23044(N38430,N38432,N38433);
and and23045(N38431,N38434,N38435);
and and23050(N38441,N38443,N38444);
and and23051(N38442,N38445,N38446);
and and23056(N38452,N38454,N38455);
and and23057(N38453,N38456,N38457);
and and23062(N38463,N38465,N38466);
and and23063(N38464,N38467,R1);
and and23068(N38473,N38475,N38476);
and and23069(N38474,N38477,R0);
and and23074(N38483,N38485,N38486);
and and23075(N38484,N38487,N38488);
and and23080(N38493,N38495,N38496);
and and23081(N38494,N38497,N38498);
and and23086(N38503,N38505,N38506);
and and23087(N38504,N38507,N38508);
and and23092(N38513,N38515,N38516);
and and23093(N38514,N38517,N38518);
and and23098(N38523,N38525,N38526);
and and23099(N38524,N38527,N38528);
and and23104(N38533,N38535,N38536);
and and23105(N38534,N38537,R0);
and and23110(N38542,N38544,N38545);
and and23111(N38543,N38546,N38547);
and and23116(N38551,N38553,N38554);
and and23117(N38552,N38555,R0);
and and23122(N38560,N38562,N38563);
and and23123(N38561,N38564,R0);
and and23128(N38569,N38571,N38572);
and and23129(N38570,N38573,R0);
and and23134(N38578,N38580,N38581);
and and23135(N38579,N38582,N38583);
and and23140(N38587,N38589,N38590);
and and23141(N38588,N38591,N38592);
and and23146(N38596,N38598,N38599);
and and23147(N38597,N38600,R1);
and and23152(N38605,N38607,N38608);
and and23153(N38606,N38609,N38610);
and and23158(N38614,N38616,N38617);
and and23159(N38615,N38618,N38619);
and and23164(N38623,N38625,N38626);
and and23165(N38624,N38627,R1);
and and23170(N38632,N38634,N38635);
and and23171(N38633,N38636,N38637);
and and23176(N38641,N38643,N38644);
and and23177(N38642,N38645,R0);
and and23182(N38650,N38652,N38653);
and and23183(N38651,N38654,R1);
and and23188(N38658,N38660,N38661);
and and23189(N38659,N38662,R0);
and and23194(N38666,N38668,N38669);
and and23195(N38667,N38670,R0);
and and23200(N38674,N38676,N38677);
and and23201(N38675,N38678,R0);
and and23206(N38682,N38684,N38685);
and and23207(N38683,N38686,R0);
and and23212(N38690,N38692,N38693);
and and23213(N38691,N38694,N38695);
and and23218(N38698,N38700,N38701);
and and23219(N38699,N38702,R0);
and and23224(N38706,N38708,N38709);
and and23225(N38707,N38710,R0);
and and23230(N38714,N38716,N38717);
and and23231(N38715,N38718,R0);
and and23236(N38722,N38724,N38725);
and and23237(N38723,N38726,N38727);
and and23242(N38730,N38732,N38733);
and and23243(N38731,N38734,R0);
and and23248(N38738,N38740,N38741);
and and23249(N38739,N38742,R2);
and and23253(N38747,N38749,N38750);
and and23254(N38748,R0,R1);
and and23258(N38756,N38758,N38759);
and and23259(N38757,R0,N38760);
and and23263(N38765,N38767,N38768);
and and23264(N38766,R0,N38769);
and and23033(N38406,N38410,N38411);
and and23034(N38407,N38412,N38413);
and and23035(N38408,N38414,N38415);
and and23036(N38409,N38416,N38417);
and and23040(N38421,R1,N38425);
and and23041(N38422,R3,N38426);
and and23042(N38423,N38427,N38428);
and and23046(N38432,N38436,N38437);
and and23047(N38433,R3,R4);
and and23048(N38434,N38438,N38439);
and and23052(N38443,N38447,R3);
and and23053(N38444,N38448,N38449);
and and23054(N38445,R6,N38450);
and and23058(N38454,N38458,N38459);
and and23059(N38455,R4,N38460);
and and23060(N38456,R6,N38461);
and and23064(N38465,N38468,R3);
and and23065(N38466,N38469,N38470);
and and23066(N38467,N38471,R7);
and and23070(N38475,N38478,N38479);
and and23071(N38476,R3,N38480);
and and23072(N38477,N38481,R7);
and and23076(N38485,N38489,R2);
and and23077(N38486,R3,N38490);
and and23078(N38487,R5,N38491);
and and23082(N38495,R2,N38499);
and and23083(N38496,N38500,R5);
and and23084(N38497,N38501,R7);
and and23088(N38505,R1,R2);
and and23089(N38506,N38509,R5);
and and23090(N38507,N38510,N38511);
and and23094(N38515,R1,N38519);
and and23095(N38516,R3,N38520);
and and23096(N38517,N38521,R7);
and and23100(N38525,N38529,R2);
and and23101(N38526,R4,N38530);
and and23102(N38527,N38531,R7);
and and23106(N38535,R1,R2);
and and23107(N38536,R3,N38538);
and and23108(N38537,N38539,N38540);
and and23112(N38544,R1,N38548);
and and23113(N38545,R3,R4);
and and23114(N38546,R5,N38549);
and and23118(N38553,R1,N38556);
and and23119(N38554,N38557,R4);
and and23120(N38555,N38558,R7);
and and23124(N38562,N38565,R2);
and and23125(N38563,R3,N38566);
and and23126(N38564,N38567,R6);
and and23130(N38571,R1,N38574);
and and23131(N38572,R3,N38575);
and and23132(N38573,R6,N38576);
and and23136(N38580,R1,N38584);
and and23137(N38581,R3,R5);
and and23138(N38582,R6,N38585);
and and23142(N38589,R1,R2);
and and23143(N38590,R3,N38593);
and and23144(N38591,N38594,R6);
and and23148(N38598,R2,R3);
and and23149(N38599,N38601,R5);
and and23150(N38600,N38602,N38603);
and and23154(N38607,R2,R3);
and and23155(N38608,R4,R5);
and and23156(N38609,N38611,N38612);
and and23160(N38616,R2,N38620);
and and23161(N38617,R4,R5);
and and23162(N38618,N38621,R7);
and and23166(N38625,R2,N38628);
and and23167(N38626,R4,N38629);
and and23168(N38627,R6,N38630);
and and23172(N38634,R2,R3);
and and23173(N38635,R4,N38638);
and and23174(N38636,R6,N38639);
and and23178(N38643,N38646,N38647);
and and23179(N38644,R3,R4);
and and23180(N38645,N38648,R7);
and and23184(N38652,N38655,R3);
and and23185(N38653,R4,N38656);
and and23186(N38654,R6,R7);
and and23190(N38660,N38663,R3);
and and23191(N38661,R4,R5);
and and23192(N38662,R6,N38664);
and and23196(N38668,N38671,R3);
and and23197(N38669,R4,N38672);
and and23198(N38670,R6,R7);
and and23202(N38676,R1,N38679);
and and23203(N38677,R4,R5);
and and23204(N38678,R6,N38680);
and and23208(N38684,R1,R2);
and and23209(N38685,R4,N38687);
and and23210(N38686,N38688,R7);
and and23214(N38692,R1,R2);
and and23215(N38693,R4,R5);
and and23216(N38694,N38696,R7);
and and23220(N38700,R1,R2);
and and23221(N38701,R3,N38703);
and and23222(N38702,R5,N38704);
and and23226(N38708,R1,R2);
and and23227(N38709,R3,R5);
and and23228(N38710,N38711,N38712);
and and23232(N38716,N38719,R3);
and and23233(N38717,R4,R5);
and and23234(N38718,N38720,R7);
and and23238(N38724,R1,R2);
and and23239(N38725,R3,N38728);
and and23240(N38726,R6,R7);
and and23244(N38732,R1,R2);
and and23245(N38733,N38735,R4);
and and23246(N38734,N38736,R6);
and and23250(N38740,N38743,R4);
and and23251(N38741,N38744,N38745);
and and23255(N38749,N38751,N38752);
and and23256(N38750,N38753,N38754);
and and23260(N38758,N38761,R4);
and and23261(N38759,N38762,N38763);
and and23265(N38767,R2,N38770);
and and23266(N38768,R4,N38771);
and and23267(N38794,N38795,N38796);
and and23274(N38807,N38808,N38809);
and and23281(N38820,N38821,N38822);
and and23288(N38833,N38834,N38835);
and and23295(N38845,N38846,N38847);
and and23302(N38856,N38857,N38858);
and and23309(N38867,N38868,N38869);
and and23316(N38878,N38879,N38880);
and and23323(N38889,N38890,N38891);
and and23330(N38900,N38901,N38902);
and and23337(N38911,N38912,N38913);
and and23344(N38922,N38923,N38924);
and and23351(N38932,N38933,N38934);
and and23358(N38942,N38943,N38944);
and and23365(N38951,N38952,N38953);
and and23372(N38960,N38961,N38962);
and and23379(N38968,N38969,N38970);
and and23386(N38976,N38977,N38978);
and and23392(N38988,N38989,N38990);
and and23398(N39000,N39001,N39002);
and and23404(N39011,N39012,N39013);
and and23410(N39021,N39022,N39023);
and and23416(N39028,N39029,N39030);
and and23268(N38795,N38797,N38798);
and and23269(N38796,N38799,N38800);
and and23275(N38808,N38810,N38811);
and and23276(N38809,N38812,N38813);
and and23282(N38821,N38823,N38824);
and and23283(N38822,N38825,N38826);
and and23289(N38834,N38836,N38837);
and and23290(N38835,N38838,N38839);
and and23296(N38846,N38848,N38849);
and and23297(N38847,N38850,N38851);
and and23303(N38857,N38859,N38860);
and and23304(N38858,N38861,N38862);
and and23310(N38868,N38870,N38871);
and and23311(N38869,N38872,N38873);
and and23317(N38879,N38881,N38882);
and and23318(N38880,N38883,N38884);
and and23324(N38890,N38892,N38893);
and and23325(N38891,N38894,N38895);
and and23331(N38901,N38903,N38904);
and and23332(N38902,N38905,N38906);
and and23338(N38912,N38914,N38915);
and and23339(N38913,N38916,N38917);
and and23345(N38923,N38925,N38926);
and and23346(N38924,N38927,N38928);
and and23352(N38933,N38935,N38936);
and and23353(N38934,N38937,N38938);
and and23359(N38943,N38945,N38946);
and and23360(N38944,N38947,N38948);
and and23366(N38952,N38954,N38955);
and and23367(N38953,N38956,N38957);
and and23373(N38961,N38963,N38964);
and and23374(N38962,N38965,N38966);
and and23380(N38969,N38971,N38972);
and and23381(N38970,N38973,N38974);
and and23387(N38977,N38979,N38980);
and and23388(N38978,N38981,N38982);
and and23393(N38989,N38991,N38992);
and and23394(N38990,N38993,N38994);
and and23399(N39001,N39003,N39004);
and and23400(N39002,N39005,R0);
and and23405(N39012,N39014,N39015);
and and23406(N39013,N39016,N39017);
and and23411(N39022,N39024,N39025);
and and23412(N39023,N39026,R0);
and and23417(N39029,N39031,N39032);
and and23418(N39030,N39033,R0);
and and23270(N38797,N38801,R1);
and and23271(N38798,N38802,N38803);
and and23272(N38799,N38804,R5);
and and23273(N38800,N38805,N38806);
and and23277(N38810,N38814,N38815);
and and23278(N38811,N38816,R3);
and and23279(N38812,N38817,R5);
and and23280(N38813,N38818,N38819);
and and23284(N38823,R0,N38827);
and and23285(N38824,N38828,N38829);
and and23286(N38825,N38830,N38831);
and and23287(N38826,N38832,R7);
and and23291(N38836,R0,N38840);
and and23292(N38837,N38841,R3);
and and23293(N38838,R4,N38842);
and and23294(N38839,N38843,N38844);
and and23298(N38848,N38852,N38853);
and and23299(N38849,N38854,R3);
and and23300(N38850,R4,N38855);
and and23301(N38851,R6,R7);
and and23305(N38859,R0,N38863);
and and23306(N38860,R2,R3);
and and23307(N38861,N38864,R5);
and and23308(N38862,N38865,N38866);
and and23312(N38870,R0,R1);
and and23313(N38871,N38874,N38875);
and and23314(N38872,R4,N38876);
and and23315(N38873,R6,N38877);
and and23319(N38881,N38885,R1);
and and23320(N38882,N38886,R3);
and and23321(N38883,R4,N38887);
and and23322(N38884,N38888,R7);
and and23326(N38892,R0,R1);
and and23327(N38893,N38896,N38897);
and and23328(N38894,N38898,N38899);
and and23329(N38895,R6,R7);
and and23333(N38903,N38907,R1);
and and23334(N38904,N38908,N38909);
and and23335(N38905,R4,R5);
and and23336(N38906,N38910,R7);
and and23340(N38914,N38918,N38919);
and and23341(N38915,R2,N38920);
and and23342(N38916,R4,N38921);
and and23343(N38917,R6,R7);
and and23347(N38925,R0,N38929);
and and23348(N38926,R2,R3);
and and23349(N38927,R4,N38930);
and and23350(N38928,R6,N38931);
and and23354(N38935,R0,N38939);
and and23355(N38936,R2,N38940);
and and23356(N38937,R4,R5);
and and23357(N38938,R6,N38941);
and and23361(N38945,R0,R1);
and and23362(N38946,N38949,R3);
and and23363(N38947,N38950,R5);
and and23364(N38948,R6,R7);
and and23368(N38954,N38958,R1);
and and23369(N38955,N38959,R3);
and and23370(N38956,R4,R5);
and and23371(N38957,R6,R7);
and and23375(N38963,R0,R1);
and and23376(N38964,R2,R3);
and and23377(N38965,R4,R5);
and and23378(N38966,R6,N38967);
and and23382(N38971,R0,R1);
and and23383(N38972,R2,R3);
and and23384(N38973,R4,R5);
and and23385(N38974,N38975,R7);
and and23389(N38979,N38983,N38984);
and and23390(N38980,N38985,R4);
and and23391(N38981,N38986,N38987);
and and23395(N38991,N38995,N38996);
and and23396(N38992,R4,N38997);
and and23397(N38993,N38998,N38999);
and and23401(N39003,N39006,N39007);
and and23402(N39004,N39008,R5);
and and23403(N39005,N39009,N39010);
and and23407(N39014,R1,R2);
and and23408(N39015,R3,N39018);
and and23409(N39016,N39019,N39020);
and and23413(N39024,R1,R2);
and and23414(N39025,R3,N39027);
and and23415(N39026,R6,R7);
and and23419(N39031,R1,R2);
and and23420(N39032,N39034,R5);
and and23421(N39033,R6,R7);
and and23422(N39080,N39081,N39082);
and and23429(N39090,N39091,N39092);
and and23436(N39099,N39100,N39101);
and and23442(N39111,N39112,N39113);
and and23448(N39123,N39124,N39125);
and and23454(N39135,N39136,N39137);
and and23460(N39147,N39148,N39149);
and and23466(N39159,N39160,N39161);
and and23472(N39170,N39171,N39172);
and and23478(N39181,N39182,N39183);
and and23484(N39192,N39193,N39194);
and and23490(N39203,N39204,N39205);
and and23496(N39214,N39215,N39216);
and and23502(N39225,N39226,N39227);
and and23508(N39236,N39237,N39238);
and and23514(N39247,N39248,N39249);
and and23520(N39257,N39258,N39259);
and and23526(N39267,N39268,N39269);
and and23532(N39277,N39278,N39279);
and and23538(N39287,N39288,N39289);
and and23544(N39297,N39298,N39299);
and and23550(N39307,N39308,N39309);
and and23556(N39317,N39318,N39319);
and and23562(N39327,N39328,N39329);
and and23568(N39337,N39338,N39339);
and and23574(N39347,N39348,N39349);
and and23580(N39357,N39358,N39359);
and and23586(N39367,N39368,N39369);
and and23592(N39377,N39378,N39379);
and and23598(N39386,N39387,N39388);
and and23604(N39395,N39396,N39397);
and and23610(N39404,N39405,N39406);
and and23616(N39413,N39414,N39415);
and and23622(N39422,N39423,N39424);
and and23628(N39431,N39432,N39433);
and and23634(N39440,N39441,N39442);
and and23640(N39448,N39449,N39450);
and and23646(N39456,N39457,N39458);
and and23652(N39464,N39465,N39466);
and and23658(N39472,N39473,N39474);
and and23664(N39480,N39481,N39482);
and and23670(N39488,N39489,N39490);
and and23676(N39496,N39497,N39498);
and and23682(N39504,N39505,N39506);
and and23688(N39512,N39513,N39514);
and and23694(N39519,N39520,N39521);
and and23423(N39081,N39083,N39084);
and and23424(N39082,N39085,N39086);
and and23430(N39091,N39093,N39094);
and and23431(N39092,N39095,N39096);
and and23437(N39100,N39102,N39103);
and and23438(N39101,N39104,N39105);
and and23443(N39112,N39114,N39115);
and and23444(N39113,N39116,N39117);
and and23449(N39124,N39126,N39127);
and and23450(N39125,N39128,N39129);
and and23455(N39136,N39138,N39139);
and and23456(N39137,N39140,N39141);
and and23461(N39148,N39150,N39151);
and and23462(N39149,N39152,N39153);
and and23467(N39160,N39162,N39163);
and and23468(N39161,N39164,N39165);
and and23473(N39171,N39173,N39174);
and and23474(N39172,N39175,N39176);
and and23479(N39182,N39184,N39185);
and and23480(N39183,N39186,R0);
and and23485(N39193,N39195,N39196);
and and23486(N39194,N39197,R0);
and and23491(N39204,N39206,N39207);
and and23492(N39205,N39208,N39209);
and and23497(N39215,N39217,N39218);
and and23498(N39216,N39219,N39220);
and and23503(N39226,N39228,N39229);
and and23504(N39227,N39230,N39231);
and and23509(N39237,N39239,N39240);
and and23510(N39238,N39241,N39242);
and and23515(N39248,N39250,N39251);
and and23516(N39249,N39252,R1);
and and23521(N39258,N39260,N39261);
and and23522(N39259,N39262,R0);
and and23527(N39268,N39270,N39271);
and and23528(N39269,N39272,R0);
and and23533(N39278,N39280,N39281);
and and23534(N39279,N39282,N39283);
and and23539(N39288,N39290,N39291);
and and23540(N39289,N39292,R0);
and and23545(N39298,N39300,N39301);
and and23546(N39299,N39302,N39303);
and and23551(N39308,N39310,N39311);
and and23552(N39309,N39312,N39313);
and and23557(N39318,N39320,N39321);
and and23558(N39319,N39322,R1);
and and23563(N39328,N39330,N39331);
and and23564(N39329,N39332,N39333);
and and23569(N39338,N39340,N39341);
and and23570(N39339,N39342,N39343);
and and23575(N39348,N39350,N39351);
and and23576(N39349,N39352,N39353);
and and23581(N39358,N39360,N39361);
and and23582(N39359,N39362,N39363);
and and23587(N39368,N39370,N39371);
and and23588(N39369,N39372,N39373);
and and23593(N39378,N39380,N39381);
and and23594(N39379,N39382,R0);
and and23599(N39387,N39389,N39390);
and and23600(N39388,N39391,N39392);
and and23605(N39396,N39398,N39399);
and and23606(N39397,N39400,R0);
and and23611(N39405,N39407,N39408);
and and23612(N39406,N39409,R0);
and and23617(N39414,N39416,N39417);
and and23618(N39415,N39418,R0);
and and23623(N39423,N39425,N39426);
and and23624(N39424,N39427,R0);
and and23629(N39432,N39434,N39435);
and and23630(N39433,N39436,R1);
and and23635(N39441,N39443,N39444);
and and23636(N39442,N39445,R0);
and and23641(N39449,N39451,N39452);
and and23642(N39450,N39453,N39454);
and and23647(N39457,N39459,N39460);
and and23648(N39458,N39461,R0);
and and23653(N39465,N39467,N39468);
and and23654(N39466,N39469,R0);
and and23659(N39473,N39475,N39476);
and and23660(N39474,N39477,N39478);
and and23665(N39481,N39483,N39484);
and and23666(N39482,N39485,N39486);
and and23671(N39489,N39491,N39492);
and and23672(N39490,N39493,N39494);
and and23677(N39497,N39499,N39500);
and and23678(N39498,N39501,R1);
and and23683(N39505,N39507,N39508);
and and23684(N39506,N39509,R0);
and and23689(N39513,N39515,N39516);
and and23690(N39514,N39517,R0);
and and23695(N39520,N39522,N39523);
and and23696(N39521,N39524,N39525);
and and23425(N39083,R0,R1);
and and23426(N39084,R2,R3);
and and23427(N39085,N39087,N39088);
and and23428(N39086,N39089,R7);
and and23432(N39093,N39097,R1);
and and23433(N39094,R2,N39098);
and and23434(N39095,R4,R5);
and and23435(N39096,R6,R7);
and and23439(N39102,R1,N39106);
and and23440(N39103,N39107,N39108);
and and23441(N39104,N39109,N39110);
and and23445(N39114,N39118,N39119);
and and23446(N39115,N39120,N39121);
and and23447(N39116,N39122,R7);
and and23451(N39126,N39130,N39131);
and and23452(N39127,N39132,N39133);
and and23453(N39128,R6,N39134);
and and23457(N39138,N39142,R2);
and and23458(N39139,N39143,N39144);
and and23459(N39140,N39145,N39146);
and and23463(N39150,N39154,N39155);
and and23464(N39151,N39156,N39157);
and and23465(N39152,N39158,R7);
and and23469(N39162,N39166,N39167);
and and23470(N39163,R3,N39168);
and and23471(N39164,N39169,R7);
and and23475(N39173,R2,R3);
and and23476(N39174,N39177,N39178);
and and23477(N39175,N39179,N39180);
and and23481(N39184,N39187,R3);
and and23482(N39185,N39188,N39189);
and and23483(N39186,N39190,N39191);
and and23487(N39195,N39198,N39199);
and and23488(N39196,N39200,N39201);
and and23489(N39197,R6,N39202);
and and23493(N39206,N39210,R2);
and and23494(N39207,N39211,N39212);
and and23495(N39208,R6,N39213);
and and23499(N39217,N39221,R2);
and and23500(N39218,R3,N39222);
and and23501(N39219,N39223,N39224);
and and23505(N39228,N39232,R2);
and and23506(N39229,N39233,R5);
and and23507(N39230,N39234,N39235);
and and23511(N39239,N39243,N39244);
and and23512(N39240,R4,N39245);
and and23513(N39241,N39246,R7);
and and23517(N39250,N39253,R3);
and and23518(N39251,R4,N39254);
and and23519(N39252,N39255,N39256);
and and23523(N39260,R1,N39263);
and and23524(N39261,N39264,N39265);
and and23525(N39262,N39266,R7);
and and23529(N39270,N39273,N39274);
and and23530(N39271,R3,N39275);
and and23531(N39272,R5,N39276);
and and23535(N39280,N39284,R2);
and and23536(N39281,R3,N39285);
and and23537(N39282,N39286,R6);
and and23541(N39290,R1,N39293);
and and23542(N39291,R4,N39294);
and and23543(N39292,N39295,N39296);
and and23547(N39300,R1,N39304);
and and23548(N39301,N39305,N39306);
and and23549(N39302,R6,R7);
and and23553(N39310,N39314,R3);
and and23554(N39311,N39315,N39316);
and and23555(N39312,R6,R7);
and and23559(N39320,N39323,N39324);
and and23560(N39321,N39325,R5);
and and23561(N39322,R6,N39326);
and and23565(N39330,N39334,R3);
and and23566(N39331,N39335,R5);
and and23567(N39332,R6,N39336);
and and23571(N39340,R1,N39344);
and and23572(N39341,N39345,R4);
and and23573(N39342,N39346,R7);
and and23577(N39350,R1,R2);
and and23578(N39351,N39354,N39355);
and and23579(N39352,N39356,R6);
and and23583(N39360,R1,N39364);
and and23584(N39361,N39365,R4);
and and23585(N39362,R6,N39366);
and and23589(N39370,R1,N39374);
and and23590(N39371,N39375,R5);
and and23591(N39372,R6,N39376);
and and23595(N39380,R1,R2);
and and23596(N39381,N39383,N39384);
and and23597(N39382,R6,N39385);
and and23601(N39389,R2,R3);
and and23602(N39390,N39393,R5);
and and23603(N39391,N39394,R7);
and and23607(N39398,R2,N39401);
and and23608(N39399,N39402,R5);
and and23609(N39400,N39403,R7);
and and23613(N39407,N39410,R2);
and and23614(N39408,N39411,N39412);
and and23615(N39409,R6,R7);
and and23619(N39416,R1,R2);
and and23620(N39417,R4,N39419);
and and23621(N39418,N39420,N39421);
and and23625(N39425,R1,N39428);
and and23626(N39426,N39429,R5);
and and23627(N39427,R6,N39430);
and and23631(N39434,N39437,N39438);
and and23632(N39435,R4,N39439);
and and23633(N39436,R6,R7);
and and23637(N39443,N39446,R2);
and and23638(N39444,R3,R4);
and and23639(N39445,N39447,R7);
and and23643(N39451,N39455,R2);
and and23644(N39452,R3,R4);
and and23645(N39453,R5,R6);
and and23649(N39459,N39462,R2);
and and23650(N39460,R3,N39463);
and and23651(N39461,R5,R6);
and and23655(N39467,R1,N39470);
and and23656(N39468,R3,R4);
and and23657(N39469,R5,N39471);
and and23661(N39475,N39479,R2);
and and23662(N39476,R3,R4);
and and23663(N39477,R5,R7);
and and23667(N39483,R1,R2);
and and23668(N39484,R3,R4);
and and23669(N39485,R5,N39487);
and and23673(N39491,R1,R3);
and and23674(N39492,N39495,R5);
and and23675(N39493,R6,R7);
and and23679(N39499,N39502,R3);
and and23680(N39500,R4,R5);
and and23681(N39501,N39503,R7);
and and23685(N39507,R1,R2);
and and23686(N39508,N39510,R5);
and and23687(N39509,N39511,R7);
and and23691(N39515,R1,N39518);
and and23692(N39516,R3,R4);
and and23693(N39517,R5,R7);
and and23697(N39522,R2,R3);
and and23698(N39523,R4,R5);
and and23699(N39524,R6,R7);

or or0(N0,N1,N2);
or or1(N1,N3,N4);
or or2(N2,N5,N6);
or or3(N3,N7,N8);
or or4(N4,N9,N10);
or or5(N5,N11,N12);
or or6(N6,N13,N14);
or or7(N7,N15,N16);
or or8(N8,N17,N18);
or or9(N9,N19,N20);
or or10(N10,N21,N22);
or or11(N11,N23,N24);
or or12(N12,N25,N26);
or or13(N13,N27,N28);
or or14(N14,N29,N30);
or or15(N15,N31,N32);
or or16(N16,N33,N34);
or or17(N17,N35,N36);
or or18(N18,N37,N38);
or or19(N19,N39,N40);
or or20(N20,N41,N42);
or or21(N21,N43,N44);
or or22(N22,N45,N46);
or or23(N23,N47,N48);
or or24(N24,N49,N50);
or or25(N25,N51,N52);
or or26(N26,N53,N54);
or or27(N27,N55,N56);
or or28(N28,N57,N58);
or or29(N29,N59,N60);
or or30(N30,N61,N62);
or or31(N31,N63,N64);
or or32(N32,N65,N66);
or or33(N33,N67,N68);
or or34(N34,N69,N70);
or or35(N35,N71,N72);
or or36(N36,N73,N74);
or or37(N37,N75,N76);
or or38(N38,N77,N78);
or or39(N39,N79,N80);
or or40(N40,N81,N82);
or or41(N41,N83,N84);
or or42(N42,N85,N86);
or or43(N43,N87,N88);
or or44(N44,N89,N90);
or or45(N45,N91,N92);
or or46(N46,N93,N94);
or or47(N47,N95,N96);
or or48(N48,N97,N98);
or or49(N49,N99,N100);
or or50(N50,N101,N102);
or or51(N51,N103,N104);
or or52(N52,N105,N106);
or or53(N53,N107,N108);
or or54(N54,N109,N110);
or or55(N55,N111,N112);
or or56(N56,N113,N114);
or or57(N57,N115,N116);
or or58(N58,N117,N118);
or or59(N59,N119,N120);
or or60(N60,N121,N122);
or or61(N61,N123,N124);
or or62(N62,N125,N126);
or or63(N63,N127,N128);
or or64(N64,N129,N130);
or or65(N65,N131,N132);
or or66(N66,N133,N134);
or or67(N67,N135,N136);
or or68(N68,N137,N138);
or or69(N69,N139,N140);
or or70(N70,N141,N142);
or or71(N71,N143,N144);
or or72(N72,N145,N146);
or or73(N73,N147,N148);
or or74(N74,N149,N150);
or or75(N75,N151,N152);
or or76(N76,N153,N154);
or or77(N77,N155,N156);
or or78(N78,N157,N158);
or or79(N79,N159,N160);
or or80(N80,N161,N162);
or or81(N81,N163,N164);
or or82(N82,N165,N166);
or or83(N83,N167,N168);
or or84(N84,N169,N170);
or or85(N85,N171,N172);
or or86(N86,N173,N174);
or or87(N87,N175,N176);
or or88(N88,N177,N178);
or or89(N89,N179,N180);
or or90(N90,N181,N182);
or or91(N91,N183,N184);
or or92(N92,N185,N186);
or or93(N93,N187,N188);
or or94(N94,N189,N190);
or or95(N95,N191,N192);
or or96(N96,N193,N194);
or or97(N97,N195,N196);
or or98(N98,N197,N198);
or or99(N99,N199,N200);
or or100(N100,N201,N202);
or or101(N101,N203,N204);
or or102(N102,N205,N206);
or or103(N103,N207,N208);
or or104(N104,N209,N210);
or or105(N105,N211,N212);
or or106(N106,N213,N214);
or or107(N107,N215,N216);
or or108(N108,N217,N218);
or or109(N109,N219,N220);
or or110(N110,N221,N222);
or or111(N111,N223,N224);
or or112(N112,N225,N226);
or or113(N113,N227,N228);
or or114(N114,N229,N230);
or or115(N115,N231,N232);
or or116(N116,N233,N234);
or or117(N117,N235,N236);
or or118(N118,N237,N238);
or or119(N119,N239,N240);
or or120(N120,N241,N242);
or or121(N121,N243,N244);
or or122(N122,N245,N246);
or or123(N123,N247,N248);
or or124(N124,N249,N250);
or or125(N125,N251,N252);
or or126(N126,N253,N254);
or or127(N127,N255,N256);
or or128(N128,N257,N258);
or or129(N129,N259,N260);
or or130(N130,N261,N262);
or or131(N131,N263,N264);
or or132(N132,N265,N266);
or or133(N133,N267,N268);
or or134(N134,N269,N270);
or or135(N135,N271,N272);
or or136(N136,N273,N274);
or or137(N137,N275,N276);
or or138(N138,N277,N278);
or or139(N139,N279,N280);
or or140(N140,N281,N282);
or or141(N141,N283,N284);
or or142(N142,N285,N286);
or or143(N143,N287,N288);
or or144(N144,N289,N290);
or or145(N145,N291,N292);
or or146(N146,N293,N294);
or or147(N147,N295,N296);
or or148(N148,N297,N298);
or or149(N149,N299,N300);
or or150(N150,N301,N302);
or or151(N151,N303,N304);
or or152(N152,N305,N306);
or or153(N153,N307,N308);
or or154(N154,N309,N310);
or or155(N155,N311,N312);
or or156(N156,N313,N314);
or or157(N157,N315,N316);
or or158(N158,N317,N318);
or or159(N159,N319,N320);
or or160(N160,N321,N322);
or or161(N161,N323,N324);
or or162(N162,N325,N326);
or or163(N163,N327,N328);
or or164(N164,N329,N330);
or or165(N165,N331,N332);
or or166(N166,N333,N334);
or or167(N167,N335,N336);
or or168(N168,N337,N338);
or or169(N169,N339,N340);
or or170(N170,N341,N342);
or or171(N171,N343,N344);
or or172(N172,N345,N346);
or or173(N173,N347,N348);
or or174(N174,N349,N350);
or or175(N175,N351,N352);
or or176(N176,N353,N354);
or or177(N177,N355,N356);
or or178(N178,N357,N358);
or or179(N179,N359,N360);
or or180(N180,N361,N362);
or or181(N181,N363,N364);
or or182(N182,N365,N366);
or or183(N183,N367,N368);
or or184(N184,N369,N370);
or or185(N185,N371,N372);
or or186(N186,N373,N374);
or or187(N187,N375,N376);
or or188(N188,N377,N378);
or or189(N189,N379,N380);
or or190(N190,N381,N382);
or or191(N191,N383,N384);
or or192(N192,N385,N386);
or or193(N193,N387,N388);
or or194(N194,N405,N422);
or or195(N195,N439,N456);
or or196(N196,N473,N489);
or or197(N197,N505,N521);
or or198(N198,N537,N553);
or or199(N199,N569,N585);
or or200(N200,N601,N617);
or or201(N201,N633,N649);
or or202(N202,N665,N681);
or or203(N203,N697,N713);
or or204(N204,N729,N745);
or or205(N205,N761,N777);
or or206(N206,N793,N809);
or or207(N207,N824,N839);
or or208(N208,N854,N869);
or or209(N209,N884,N899);
or or210(N210,N914,N929);
or or211(N211,N944,N959);
or or212(N212,N974,N989);
or or213(N213,N1004,N1019);
or or214(N214,N1034,N1049);
or or215(N215,N1064,N1079);
or or216(N216,N1094,N1109);
or or217(N217,N1124,N1139);
or or218(N218,N1154,N1169);
or or219(N219,N1184,N1199);
or or220(N220,N1214,N1229);
or or221(N221,N1244,N1259);
or or222(N222,N1274,N1289);
or or223(N223,N1304,N1319);
or or224(N224,N1334,N1349);
or or225(N225,N1364,N1379);
or or226(N226,N1394,N1409);
or or227(N227,N1424,N1438);
or or228(N228,N1452,N1466);
or or229(N229,N1480,N1494);
or or230(N230,N1508,N1522);
or or231(N231,N1536,N1550);
or or232(N232,N1564,N1578);
or or233(N233,N1592,N1606);
or or234(N234,N1620,N1634);
or or235(N235,N1648,N1662);
or or236(N236,N1676,N1690);
or or237(N237,N1704,N1718);
or or238(N238,N1732,N1746);
or or239(N239,N1760,N1774);
or or240(N240,N1788,N1802);
or or241(N241,N1816,N1830);
or or242(N242,N1844,N1858);
or or243(N243,N1872,N1886);
or or244(N244,N1900,N1914);
or or245(N245,N1928,N1942);
or or246(N246,N1956,N1970);
or or247(N247,N1984,N1998);
or or248(N248,N2012,N2026);
or or249(N249,N2040,N2054);
or or250(N250,N2068,N2082);
or or251(N251,N2096,N2110);
or or252(N252,N2123,N2136);
or or253(N253,N2149,N2162);
or or254(N254,N2175,N2188);
or or255(N255,N2201,N2214);
or or256(N256,N2227,N2240);
or or257(N257,N2253,N2266);
or or258(N258,N2279,N2292);
or or259(N259,N2305,N2318);
or or260(N260,N2331,N2344);
or or261(N261,N2357,N2370);
or or262(N262,N2383,N2396);
or or263(N263,N2409,N2422);
or or264(N264,N2435,N2448);
or or265(N265,N2461,N2474);
or or266(N266,N2487,N2500);
or or267(N267,N2513,N2526);
or or268(N268,N2539,N2552);
or or269(N269,N2565,N2578);
or or270(N270,N2591,N2604);
or or271(N271,N2616,N2628);
or or272(N272,N2640,N2652);
or or273(N273,N2664,N2676);
or or274(N274,N2688,N2700);
or or275(N275,N2712,N2724);
or or276(N276,N2736,N2748);
or or277(N277,N2760,N2772);
or or278(N278,N2784,N2796);
or or279(N279,N2808,N2820);
or or280(N280,N2832,N2844);
or or281(N281,N2856,N2868);
or or282(N282,N2880,N2892);
or or283(N283,N2904,N2916);
or or284(N284,N2928,N2940);
or or285(N285,N2952,N2964);
or or286(N286,N2976,N2988);
or or287(N287,N3000,N3012);
or or288(N288,N3024,N3036);
or or289(N289,N3048,N3060);
or or290(N290,N3072,N3084);
or or291(N291,N3095,N3106);
or or292(N292,N3117,N3128);
or or293(N293,N3139,N3150);
or or294(N294,N3161,N3172);
or or295(N295,N3183,N3194);
or or296(N296,N3205,N3216);
or or297(N297,N3227,N3237);
or or298(N298,N3247,N3256);
or or299(N299,N3272,N3288);
or or300(N300,N3304,N3320);
or or301(N301,N3336,N3352);
or or302(N302,N3368,N3383);
or or303(N303,N3398,N3413);
or or304(N304,N3428,N3443);
or or305(N305,N3458,N3473);
or or306(N306,N3488,N3503);
or or307(N307,N3518,N3532);
or or308(N308,N3546,N3560);
or or309(N309,N3574,N3588);
or or310(N310,N3602,N3616);
or or311(N311,N3630,N3644);
or or312(N312,N3658,N3672);
or or313(N313,N3686,N3700);
or or314(N314,N3714,N3728);
or or315(N315,N3742,N3756);
or or316(N316,N3770,N3784);
or or317(N317,N3798,N3812);
or or318(N318,N3826,N3840);
or or319(N319,N3854,N3868);
or or320(N320,N3882,N3895);
or or321(N321,N3908,N3921);
or or322(N322,N3934,N3947);
or or323(N323,N3960,N3973);
or or324(N324,N3986,N3999);
or or325(N325,N4012,N4025);
or or326(N326,N4038,N4051);
or or327(N327,N4064,N4077);
or or328(N328,N4090,N4103);
or or329(N329,N4116,N4129);
or or330(N330,N4142,N4155);
or or331(N331,N4168,N4181);
or or332(N332,N4194,N4207);
or or333(N333,N4220,N4233);
or or334(N334,N4246,N4259);
or or335(N335,N4272,N4285);
or or336(N336,N4298,N4311);
or or337(N337,N4324,N4337);
or or338(N338,N4350,N4363);
or or339(N339,N4376,N4389);
or or340(N340,N4402,N4415);
or or341(N341,N4428,N4441);
or or342(N342,N4454,N4467);
or or343(N343,N4480,N4493);
or or344(N344,N4505,N4517);
or or345(N345,N4529,N4541);
or or346(N346,N4553,N4565);
or or347(N347,N4577,N4589);
or or348(N348,N4601,N4613);
or or349(N349,N4625,N4637);
or or350(N350,N4649,N4661);
or or351(N351,N4673,N4685);
or or352(N352,N4697,N4709);
or or353(N353,N4721,N4733);
or or354(N354,N4745,N4757);
or or355(N355,N4769,N4781);
or or356(N356,N4793,N4805);
or or357(N357,N4817,N4829);
or or358(N358,N4841,N4853);
or or359(N359,N4865,N4877);
or or360(N360,N4889,N4901);
or or361(N361,N4913,N4925);
or or362(N362,N4937,N4949);
or or363(N363,N4961,N4973);
or or364(N364,N4984,N4995);
or or365(N365,N5006,N5017);
or or366(N366,N5028,N5039);
or or367(N367,N5050,N5061);
or or368(N368,N5072,N5083);
or or369(N369,N5094,N5105);
or or370(N370,N5116,N5127);
or or371(N371,N5138,N5149);
or or372(N372,N5160,N5171);
or or373(N373,N5182,N5192);
or or374(N374,N5202,N5212);
or or375(N375,N5222,N5232);
or or376(N376,N5242,N5252);
or or377(N377,N5261,N5270);
or or378(N378,N5279,N5293);
or or379(N379,N5306,N5319);
or or380(N380,N5331,N5343);
or or381(N381,N5355,N5367);
or or382(N382,N5378,N5389);
or or383(N383,N5400,N5411);
or or384(N384,N5422,N5432);
or or385(N385,N5442,N5452);
or or386(N386,N5462,N5471);
or or387(N387,N5480,N5489);
or or388(N5497,N5498,N5499);
or or389(N5498,N5500,N5501);
or or390(N5499,N5502,N5503);
or or391(N5500,N5504,N5505);
or or392(N5501,N5506,N5507);
or or393(N5502,N5508,N5509);
or or394(N5503,N5510,N5511);
or or395(N5504,N5512,N5513);
or or396(N5505,N5514,N5515);
or or397(N5506,N5516,N5517);
or or398(N5507,N5518,N5519);
or or399(N5508,N5520,N5521);
or or400(N5509,N5522,N5523);
or or401(N5510,N5524,N5525);
or or402(N5511,N5526,N5527);
or or403(N5512,N5528,N5529);
or or404(N5513,N5530,N5531);
or or405(N5514,N5532,N5533);
or or406(N5515,N5534,N5535);
or or407(N5516,N5536,N5537);
or or408(N5517,N5538,N5539);
or or409(N5518,N5540,N5541);
or or410(N5519,N5542,N5543);
or or411(N5520,N5544,N5545);
or or412(N5521,N5546,N5547);
or or413(N5522,N5548,N5549);
or or414(N5523,N5550,N5551);
or or415(N5524,N5552,N5553);
or or416(N5525,N5554,N5555);
or or417(N5526,N5556,N5557);
or or418(N5527,N5558,N5559);
or or419(N5528,N5560,N5561);
or or420(N5529,N5562,N5563);
or or421(N5530,N5564,N5565);
or or422(N5531,N5566,N5567);
or or423(N5532,N5568,N5569);
or or424(N5533,N5570,N5571);
or or425(N5534,N5572,N5573);
or or426(N5535,N5574,N5575);
or or427(N5536,N5576,N5577);
or or428(N5537,N5578,N5579);
or or429(N5538,N5580,N5581);
or or430(N5539,N5582,N5583);
or or431(N5540,N5584,N5585);
or or432(N5541,N5586,N5587);
or or433(N5542,N5588,N5589);
or or434(N5543,N5590,N5591);
or or435(N5544,N5592,N5593);
or or436(N5545,N5594,N5595);
or or437(N5546,N5596,N5597);
or or438(N5547,N5598,N5599);
or or439(N5548,N5600,N5601);
or or440(N5549,N5602,N5603);
or or441(N5550,N5604,N5605);
or or442(N5551,N5606,N5607);
or or443(N5552,N5608,N5609);
or or444(N5553,N5610,N5611);
or or445(N5554,N5612,N5613);
or or446(N5555,N5614,N5615);
or or447(N5556,N5616,N5617);
or or448(N5557,N5618,N5619);
or or449(N5558,N5620,N5621);
or or450(N5559,N5622,N5623);
or or451(N5560,N5624,N5625);
or or452(N5561,N5626,N5627);
or or453(N5562,N5628,N5629);
or or454(N5563,N5630,N5631);
or or455(N5564,N5632,N5633);
or or456(N5565,N5634,N5635);
or or457(N5566,N5636,N5637);
or or458(N5567,N5638,N5639);
or or459(N5568,N5640,N5641);
or or460(N5569,N5642,N5643);
or or461(N5570,N5644,N5645);
or or462(N5571,N5646,N5647);
or or463(N5572,N5648,N5649);
or or464(N5573,N5650,N5651);
or or465(N5574,N5652,N5653);
or or466(N5575,N5654,N5655);
or or467(N5576,N5656,N5657);
or or468(N5577,N5658,N5659);
or or469(N5578,N5660,N5661);
or or470(N5579,N5662,N5663);
or or471(N5580,N5664,N5665);
or or472(N5581,N5666,N5667);
or or473(N5582,N5668,N5669);
or or474(N5583,N5670,N5671);
or or475(N5584,N5672,N5673);
or or476(N5585,N5674,N5675);
or or477(N5586,N5676,N5677);
or or478(N5587,N5678,N5679);
or or479(N5588,N5680,N5681);
or or480(N5589,N5682,N5683);
or or481(N5590,N5684,N5685);
or or482(N5591,N5686,N5687);
or or483(N5592,N5688,N5689);
or or484(N5593,N5690,N5691);
or or485(N5594,N5692,N5693);
or or486(N5595,N5694,N5695);
or or487(N5596,N5696,N5697);
or or488(N5597,N5698,N5699);
or or489(N5598,N5700,N5701);
or or490(N5599,N5702,N5703);
or or491(N5600,N5704,N5705);
or or492(N5601,N5706,N5707);
or or493(N5602,N5708,N5709);
or or494(N5603,N5710,N5711);
or or495(N5604,N5712,N5713);
or or496(N5605,N5714,N5715);
or or497(N5606,N5716,N5717);
or or498(N5607,N5718,N5719);
or or499(N5608,N5720,N5721);
or or500(N5609,N5722,N5723);
or or501(N5610,N5724,N5725);
or or502(N5611,N5726,N5727);
or or503(N5612,N5728,N5729);
or or504(N5613,N5730,N5731);
or or505(N5614,N5732,N5733);
or or506(N5615,N5734,N5735);
or or507(N5616,N5736,N5737);
or or508(N5617,N5738,N5739);
or or509(N5618,N5740,N5741);
or or510(N5619,N5742,N5743);
or or511(N5620,N5744,N5745);
or or512(N5621,N5746,N5747);
or or513(N5622,N5748,N5749);
or or514(N5623,N5750,N5751);
or or515(N5624,N5752,N5753);
or or516(N5625,N5754,N5755);
or or517(N5626,N5756,N5757);
or or518(N5627,N5758,N5759);
or or519(N5628,N5760,N5761);
or or520(N5629,N5762,N5763);
or or521(N5630,N5764,N5765);
or or522(N5631,N5766,N5767);
or or523(N5632,N5768,N5769);
or or524(N5633,N5770,N5771);
or or525(N5634,N5772,N5773);
or or526(N5635,N5774,N5775);
or or527(N5636,N5776,N5777);
or or528(N5637,N5778,N5779);
or or529(N5638,N5780,N5781);
or or530(N5639,N5782,N5783);
or or531(N5640,N5784,N5785);
or or532(N5641,N5786,N5787);
or or533(N5642,N5788,N5789);
or or534(N5643,N5790,N5791);
or or535(N5644,N5792,N5793);
or or536(N5645,N5794,N5795);
or or537(N5646,N5796,N5797);
or or538(N5647,N5798,N5799);
or or539(N5648,N5800,N5801);
or or540(N5649,N5802,N5803);
or or541(N5650,N5804,N5805);
or or542(N5651,N5806,N5807);
or or543(N5652,N5808,N5809);
or or544(N5653,N5810,N5811);
or or545(N5654,N5812,N5813);
or or546(N5655,N5814,N5815);
or or547(N5656,N5816,N5817);
or or548(N5657,N5818,N5819);
or or549(N5658,N5820,N5821);
or or550(N5659,N5822,N5823);
or or551(N5660,N5824,N5825);
or or552(N5661,N5826,N5827);
or or553(N5662,N5828,N5829);
or or554(N5663,N5830,N5831);
or or555(N5664,N5832,N5833);
or or556(N5665,N5834,N5835);
or or557(N5666,N5836,N5837);
or or558(N5667,N5838,N5839);
or or559(N5668,N5840,N5841);
or or560(N5669,N5842,N5843);
or or561(N5670,N5844,N5845);
or or562(N5671,N5846,N5847);
or or563(N5672,N5848,N5849);
or or564(N5673,N5850,N5851);
or or565(N5674,N5852,N5853);
or or566(N5675,N5854,N5855);
or or567(N5676,N5856,N5857);
or or568(N5677,N5858,N5859);
or or569(N5678,N5860,N5861);
or or570(N5679,N5862,N5863);
or or571(N5680,N5864,N5865);
or or572(N5681,N5866,N5867);
or or573(N5682,N5868,N5869);
or or574(N5683,N5870,N5871);
or or575(N5684,N5872,N5873);
or or576(N5685,N5874,N5875);
or or577(N5686,N5876,N5877);
or or578(N5687,N5878,N5879);
or or579(N5688,N5880,N5881);
or or580(N5689,N5882,N5883);
or or581(N5690,N5884,N5885);
or or582(N5691,N5886,N5887);
or or583(N5692,N5888,N5889);
or or584(N5693,N5890,N5891);
or or585(N5694,N5892,N5893);
or or586(N5695,N5894,N5895);
or or587(N5696,N5896,N5897);
or or588(N5697,N5898,N5899);
or or589(N5698,N5900,N5901);
or or590(N5699,N5902,N5903);
or or591(N5700,N5904,N5905);
or or592(N5701,N5906,N5907);
or or593(N5702,N5908,N5909);
or or594(N5703,N5910,N5911);
or or595(N5704,N5912,N5913);
or or596(N5705,N5914,N5915);
or or597(N5706,N5916,N5917);
or or598(N5707,N5918,N5919);
or or599(N5708,N5920,N5921);
or or600(N5709,N5922,N5923);
or or601(N5710,N5924,N5925);
or or602(N5711,N5926,N5927);
or or603(N5712,N5928,N5929);
or or604(N5713,N5930,N5931);
or or605(N5714,N5949,N5967);
or or606(N5715,N5985,N6002);
or or607(N5716,N6019,N6036);
or or608(N5717,N6053,N6069);
or or609(N5718,N6085,N6101);
or or610(N5719,N6117,N6133);
or or611(N5720,N6149,N6165);
or or612(N5721,N6181,N6197);
or or613(N5722,N6213,N6229);
or or614(N5723,N6245,N6261);
or or615(N5724,N6277,N6293);
or or616(N5725,N6308,N6323);
or or617(N5726,N6338,N6353);
or or618(N5727,N6368,N6383);
or or619(N5728,N6398,N6413);
or or620(N5729,N6428,N6443);
or or621(N5730,N6458,N6473);
or or622(N5731,N6488,N6503);
or or623(N5732,N6518,N6533);
or or624(N5733,N6548,N6563);
or or625(N5734,N6578,N6593);
or or626(N5735,N6608,N6623);
or or627(N5736,N6638,N6653);
or or628(N5737,N6668,N6683);
or or629(N5738,N6698,N6712);
or or630(N5739,N6726,N6740);
or or631(N5740,N6754,N6768);
or or632(N5741,N6782,N6796);
or or633(N5742,N6810,N6824);
or or634(N5743,N6838,N6852);
or or635(N5744,N6866,N6880);
or or636(N5745,N6894,N6908);
or or637(N5746,N6922,N6936);
or or638(N5747,N6950,N6964);
or or639(N5748,N6978,N6992);
or or640(N5749,N7006,N7020);
or or641(N5750,N7034,N7048);
or or642(N5751,N7062,N7076);
or or643(N5752,N7090,N7104);
or or644(N5753,N7118,N7131);
or or645(N5754,N7144,N7157);
or or646(N5755,N7170,N7183);
or or647(N5756,N7196,N7209);
or or648(N5757,N7222,N7235);
or or649(N5758,N7248,N7261);
or or650(N5759,N7274,N7287);
or or651(N5760,N7300,N7313);
or or652(N5761,N7326,N7339);
or or653(N5762,N7352,N7365);
or or654(N5763,N7378,N7391);
or or655(N5764,N7404,N7417);
or or656(N5765,N7430,N7443);
or or657(N5766,N7456,N7469);
or or658(N5767,N7482,N7495);
or or659(N5768,N7508,N7521);
or or660(N5769,N7534,N7547);
or or661(N5770,N7560,N7573);
or or662(N5771,N7586,N7599);
or or663(N5772,N7612,N7624);
or or664(N5773,N7636,N7648);
or or665(N5774,N7660,N7672);
or or666(N5775,N7684,N7696);
or or667(N5776,N7708,N7720);
or or668(N5777,N7732,N7744);
or or669(N5778,N7756,N7768);
or or670(N5779,N7780,N7792);
or or671(N5780,N7804,N7816);
or or672(N5781,N7828,N7840);
or or673(N5782,N7852,N7864);
or or674(N5783,N7876,N7888);
or or675(N5784,N7900,N7911);
or or676(N5785,N7922,N7933);
or or677(N5786,N7944,N7955);
or or678(N5787,N7966,N7977);
or or679(N5788,N7988,N7999);
or or680(N5789,N8010,N8021);
or or681(N5790,N8032,N8042);
or or682(N5791,N8052,N8062);
or or683(N5792,N8072,N8082);
or or684(N5793,N8092,N8102);
or or685(N5794,N8112,N8121);
or or686(N5795,N8137,N8153);
or or687(N5796,N8168,N8183);
or or688(N5797,N8198,N8213);
or or689(N5798,N8228,N8243);
or or690(N5799,N8258,N8273);
or or691(N5800,N8288,N8303);
or or692(N5801,N8318,N8333);
or or693(N5802,N8348,N8363);
or or694(N5803,N8377,N8391);
or or695(N5804,N8405,N8419);
or or696(N5805,N8433,N8447);
or or697(N5806,N8461,N8475);
or or698(N5807,N8489,N8503);
or or699(N5808,N8517,N8531);
or or700(N5809,N8545,N8559);
or or701(N5810,N8573,N8587);
or or702(N5811,N8601,N8615);
or or703(N5812,N8629,N8643);
or or704(N5813,N8657,N8671);
or or705(N5814,N8685,N8699);
or or706(N5815,N8713,N8727);
or or707(N5816,N8741,N8755);
or or708(N5817,N8769,N8783);
or or709(N5818,N8797,N8811);
or or710(N5819,N8825,N8839);
or or711(N5820,N8853,N8867);
or or712(N5821,N8881,N8895);
or or713(N5822,N8908,N8921);
or or714(N5823,N8934,N8947);
or or715(N5824,N8960,N8973);
or or716(N5825,N8986,N8999);
or or717(N5826,N9012,N9025);
or or718(N5827,N9038,N9051);
or or719(N5828,N9064,N9077);
or or720(N5829,N9090,N9103);
or or721(N5830,N9116,N9129);
or or722(N5831,N9142,N9155);
or or723(N5832,N9168,N9181);
or or724(N5833,N9194,N9207);
or or725(N5834,N9220,N9233);
or or726(N5835,N9246,N9259);
or or727(N5836,N9272,N9285);
or or728(N5837,N9298,N9311);
or or729(N5838,N9324,N9337);
or or730(N5839,N9350,N9363);
or or731(N5840,N9376,N9389);
or or732(N5841,N9402,N9415);
or or733(N5842,N9428,N9441);
or or734(N5843,N9454,N9467);
or or735(N5844,N9480,N9493);
or or736(N5845,N9506,N9519);
or or737(N5846,N9532,N9545);
or or738(N5847,N9558,N9571);
or or739(N5848,N9584,N9597);
or or740(N5849,N9610,N9623);
or or741(N5850,N9636,N9648);
or or742(N5851,N9660,N9672);
or or743(N5852,N9684,N9696);
or or744(N5853,N9708,N9720);
or or745(N5854,N9732,N9744);
or or746(N5855,N9756,N9768);
or or747(N5856,N9780,N9792);
or or748(N5857,N9804,N9816);
or or749(N5858,N9828,N9840);
or or750(N5859,N9852,N9864);
or or751(N5860,N9876,N9888);
or or752(N5861,N9900,N9912);
or or753(N5862,N9924,N9936);
or or754(N5863,N9948,N9960);
or or755(N5864,N9972,N9984);
or or756(N5865,N9996,N10008);
or or757(N5866,N10020,N10032);
or or758(N5867,N10044,N10056);
or or759(N5868,N10068,N10080);
or or760(N5869,N10092,N10104);
or or761(N5870,N10116,N10128);
or or762(N5871,N10140,N10152);
or or763(N5872,N10164,N10176);
or or764(N5873,N10188,N10200);
or or765(N5874,N10211,N10222);
or or766(N5875,N10233,N10244);
or or767(N5876,N10255,N10266);
or or768(N5877,N10277,N10288);
or or769(N5878,N10299,N10310);
or or770(N5879,N10321,N10332);
or or771(N5880,N10343,N10354);
or or772(N5881,N10365,N10376);
or or773(N5882,N10387,N10398);
or or774(N5883,N10409,N10420);
or or775(N5884,N10431,N10442);
or or776(N5885,N10453,N10464);
or or777(N5886,N10475,N10486);
or or778(N5887,N10497,N10508);
or or779(N5888,N10519,N10530);
or or780(N5889,N10541,N10552);
or or781(N5890,N10563,N10574);
or or782(N5891,N10585,N10596);
or or783(N5892,N10607,N10618);
or or784(N5893,N10629,N10640);
or or785(N5894,N10651,N10662);
or or786(N5895,N10673,N10683);
or or787(N5896,N10693,N10703);
or or788(N5897,N10713,N10723);
or or789(N5898,N10733,N10743);
or or790(N5899,N10753,N10763);
or or791(N5900,N10773,N10783);
or or792(N5901,N10793,N10803);
or or793(N5902,N10813,N10823);
or or794(N5903,N10833,N10843);
or or795(N5904,N10853,N10863);
or or796(N5905,N10873,N10883);
or or797(N5906,N10893,N10903);
or or798(N5907,N10913,N10923);
or or799(N5908,N10932,N10941);
or or800(N5909,N10950,N10959);
or or801(N5910,N10968,N10981);
or or802(N5911,N10994,N11007);
or or803(N5912,N11019,N11031);
or or804(N5913,N11043,N11055);
or or805(N5914,N11067,N11079);
or or806(N5915,N11091,N11103);
or or807(N5916,N11115,N11126);
or or808(N5917,N11137,N11148);
or or809(N5918,N11159,N11170);
or or810(N5919,N11181,N11192);
or or811(N5920,N11203,N11214);
or or812(N5921,N11225,N11236);
or or813(N5922,N11247,N11258);
or or814(N5923,N11269,N11279);
or or815(N5924,N11289,N11299);
or or816(N5925,N11309,N11319);
or or817(N5926,N11329,N11339);
or or818(N5927,N11349,N11359);
or or819(N5928,N11369,N11379);
or or820(N5929,N11389,N11399);
or or821(N5930,N11408,N11420);
or or822(N11430,N11431,N11432);
or or823(N11431,N11433,N11434);
or or824(N11432,N11435,N11436);
or or825(N11433,N11437,N11438);
or or826(N11434,N11439,N11440);
or or827(N11435,N11441,N11442);
or or828(N11436,N11443,N11444);
or or829(N11437,N11445,N11446);
or or830(N11438,N11447,N11448);
or or831(N11439,N11449,N11450);
or or832(N11440,N11451,N11452);
or or833(N11441,N11453,N11454);
or or834(N11442,N11455,N11456);
or or835(N11443,N11457,N11458);
or or836(N11444,N11459,N11460);
or or837(N11445,N11461,N11462);
or or838(N11446,N11463,N11464);
or or839(N11447,N11465,N11466);
or or840(N11448,N11467,N11468);
or or841(N11449,N11469,N11470);
or or842(N11450,N11471,N11472);
or or843(N11451,N11473,N11474);
or or844(N11452,N11475,N11476);
or or845(N11453,N11477,N11478);
or or846(N11454,N11479,N11480);
or or847(N11455,N11481,N11482);
or or848(N11456,N11483,N11484);
or or849(N11457,N11485,N11486);
or or850(N11458,N11487,N11488);
or or851(N11459,N11489,N11490);
or or852(N11460,N11491,N11492);
or or853(N11461,N11493,N11494);
or or854(N11462,N11495,N11496);
or or855(N11463,N11497,N11498);
or or856(N11464,N11499,N11500);
or or857(N11465,N11501,N11502);
or or858(N11466,N11503,N11504);
or or859(N11467,N11505,N11506);
or or860(N11468,N11507,N11508);
or or861(N11469,N11509,N11510);
or or862(N11470,N11511,N11512);
or or863(N11471,N11513,N11514);
or or864(N11472,N11515,N11516);
or or865(N11473,N11517,N11518);
or or866(N11474,N11519,N11520);
or or867(N11475,N11521,N11522);
or or868(N11476,N11523,N11524);
or or869(N11477,N11525,N11526);
or or870(N11478,N11527,N11528);
or or871(N11479,N11529,N11530);
or or872(N11480,N11531,N11532);
or or873(N11481,N11533,N11534);
or or874(N11482,N11535,N11536);
or or875(N11483,N11537,N11538);
or or876(N11484,N11539,N11540);
or or877(N11485,N11541,N11542);
or or878(N11486,N11543,N11544);
or or879(N11487,N11545,N11546);
or or880(N11488,N11547,N11548);
or or881(N11489,N11549,N11550);
or or882(N11490,N11551,N11552);
or or883(N11491,N11553,N11554);
or or884(N11492,N11555,N11556);
or or885(N11493,N11557,N11558);
or or886(N11494,N11559,N11560);
or or887(N11495,N11561,N11562);
or or888(N11496,N11563,N11564);
or or889(N11497,N11565,N11566);
or or890(N11498,N11567,N11568);
or or891(N11499,N11569,N11570);
or or892(N11500,N11571,N11572);
or or893(N11501,N11573,N11574);
or or894(N11502,N11575,N11576);
or or895(N11503,N11577,N11578);
or or896(N11504,N11579,N11580);
or or897(N11505,N11581,N11582);
or or898(N11506,N11583,N11584);
or or899(N11507,N11585,N11586);
or or900(N11508,N11587,N11588);
or or901(N11509,N11589,N11590);
or or902(N11510,N11591,N11592);
or or903(N11511,N11593,N11594);
or or904(N11512,N11595,N11596);
or or905(N11513,N11597,N11598);
or or906(N11514,N11599,N11600);
or or907(N11515,N11601,N11602);
or or908(N11516,N11603,N11604);
or or909(N11517,N11605,N11606);
or or910(N11518,N11607,N11608);
or or911(N11519,N11609,N11610);
or or912(N11520,N11611,N11612);
or or913(N11521,N11613,N11614);
or or914(N11522,N11615,N11616);
or or915(N11523,N11617,N11618);
or or916(N11524,N11619,N11620);
or or917(N11525,N11621,N11622);
or or918(N11526,N11623,N11624);
or or919(N11527,N11625,N11626);
or or920(N11528,N11627,N11628);
or or921(N11529,N11629,N11630);
or or922(N11530,N11631,N11632);
or or923(N11531,N11633,N11634);
or or924(N11532,N11635,N11636);
or or925(N11533,N11637,N11638);
or or926(N11534,N11639,N11640);
or or927(N11535,N11641,N11642);
or or928(N11536,N11643,N11644);
or or929(N11537,N11645,N11646);
or or930(N11538,N11647,N11648);
or or931(N11539,N11649,N11650);
or or932(N11540,N11651,N11652);
or or933(N11541,N11653,N11654);
or or934(N11542,N11655,N11656);
or or935(N11543,N11657,N11658);
or or936(N11544,N11659,N11660);
or or937(N11545,N11661,N11662);
or or938(N11546,N11663,N11664);
or or939(N11547,N11665,N11666);
or or940(N11548,N11667,N11668);
or or941(N11549,N11669,N11670);
or or942(N11550,N11671,N11672);
or or943(N11551,N11673,N11674);
or or944(N11552,N11675,N11676);
or or945(N11553,N11677,N11678);
or or946(N11554,N11679,N11680);
or or947(N11555,N11681,N11682);
or or948(N11556,N11683,N11684);
or or949(N11557,N11685,N11686);
or or950(N11558,N11687,N11688);
or or951(N11559,N11689,N11690);
or or952(N11560,N11691,N11692);
or or953(N11561,N11693,N11694);
or or954(N11562,N11695,N11696);
or or955(N11563,N11697,N11698);
or or956(N11564,N11699,N11700);
or or957(N11565,N11701,N11702);
or or958(N11566,N11703,N11704);
or or959(N11567,N11705,N11706);
or or960(N11568,N11707,N11708);
or or961(N11569,N11709,N11710);
or or962(N11570,N11711,N11712);
or or963(N11571,N11713,N11714);
or or964(N11572,N11715,N11716);
or or965(N11573,N11717,N11718);
or or966(N11574,N11719,N11720);
or or967(N11575,N11721,N11722);
or or968(N11576,N11723,N11724);
or or969(N11577,N11725,N11726);
or or970(N11578,N11727,N11728);
or or971(N11579,N11729,N11730);
or or972(N11580,N11731,N11732);
or or973(N11581,N11733,N11734);
or or974(N11582,N11735,N11736);
or or975(N11583,N11737,N11738);
or or976(N11584,N11739,N11740);
or or977(N11585,N11741,N11742);
or or978(N11586,N11743,N11744);
or or979(N11587,N11745,N11746);
or or980(N11588,N11747,N11748);
or or981(N11589,N11749,N11750);
or or982(N11590,N11751,N11752);
or or983(N11591,N11753,N11754);
or or984(N11592,N11755,N11756);
or or985(N11593,N11757,N11758);
or or986(N11594,N11759,N11760);
or or987(N11595,N11761,N11762);
or or988(N11596,N11763,N11764);
or or989(N11597,N11765,N11766);
or or990(N11598,N11767,N11768);
or or991(N11599,N11769,N11770);
or or992(N11600,N11771,N11772);
or or993(N11601,N11773,N11774);
or or994(N11602,N11775,N11776);
or or995(N11603,N11777,N11778);
or or996(N11604,N11779,N11780);
or or997(N11605,N11781,N11782);
or or998(N11606,N11783,N11784);
or or999(N11607,N11785,N11786);
or or1000(N11608,N11787,N11788);
or or1001(N11609,N11789,N11790);
or or1002(N11610,N11791,N11792);
or or1003(N11611,N11793,N11794);
or or1004(N11612,N11795,N11796);
or or1005(N11613,N11797,N11798);
or or1006(N11614,N11799,N11800);
or or1007(N11615,N11801,N11802);
or or1008(N11616,N11803,N11804);
or or1009(N11617,N11805,N11806);
or or1010(N11618,N11807,N11808);
or or1011(N11619,N11809,N11810);
or or1012(N11620,N11811,N11812);
or or1013(N11621,N11813,N11814);
or or1014(N11622,N11815,N11816);
or or1015(N11623,N11817,N11818);
or or1016(N11624,N11819,N11820);
or or1017(N11625,N11821,N11822);
or or1018(N11626,N11823,N11824);
or or1019(N11627,N11825,N11826);
or or1020(N11628,N11827,N11828);
or or1021(N11629,N11829,N11830);
or or1022(N11630,N11831,N11832);
or or1023(N11631,N11833,N11834);
or or1024(N11632,N11835,N11836);
or or1025(N11633,N11837,N11838);
or or1026(N11634,N11839,N11840);
or or1027(N11635,N11841,N11842);
or or1028(N11636,N11843,N11844);
or or1029(N11637,N11845,N11846);
or or1030(N11638,N11847,N11848);
or or1031(N11639,N11849,N11850);
or or1032(N11640,N11851,N11852);
or or1033(N11641,N11853,N11854);
or or1034(N11642,N11855,N11856);
or or1035(N11643,N11857,N11858);
or or1036(N11644,N11859,N11860);
or or1037(N11645,N11861,N11862);
or or1038(N11646,N11863,N11864);
or or1039(N11647,N11865,N11866);
or or1040(N11648,N11867,N11868);
or or1041(N11649,N11869,N11870);
or or1042(N11650,N11871,N11872);
or or1043(N11651,N11873,N11874);
or or1044(N11652,N11875,N11876);
or or1045(N11653,N11877,N11878);
or or1046(N11654,N11879,N11880);
or or1047(N11655,N11881,N11882);
or or1048(N11656,N11900,N11918);
or or1049(N11657,N11935,N11952);
or or1050(N11658,N11969,N11986);
or or1051(N11659,N12002,N12018);
or or1052(N11660,N12034,N12050);
or or1053(N11661,N12066,N12082);
or or1054(N11662,N12098,N12114);
or or1055(N11663,N12130,N12146);
or or1056(N11664,N12162,N12178);
or or1057(N11665,N12194,N12209);
or or1058(N11666,N12224,N12239);
or or1059(N11667,N12254,N12269);
or or1060(N11668,N12284,N12299);
or or1061(N11669,N12314,N12329);
or or1062(N11670,N12344,N12359);
or or1063(N11671,N12374,N12389);
or or1064(N11672,N12404,N12419);
or or1065(N11673,N12434,N12449);
or or1066(N11674,N12464,N12479);
or or1067(N11675,N12494,N12509);
or or1068(N11676,N12524,N12539);
or or1069(N11677,N12554,N12569);
or or1070(N11678,N12584,N12599);
or or1071(N11679,N12614,N12629);
or or1072(N11680,N12644,N12659);
or or1073(N11681,N12674,N12689);
or or1074(N11682,N12704,N12719);
or or1075(N11683,N12734,N12749);
or or1076(N11684,N12763,N12777);
or or1077(N11685,N12791,N12805);
or or1078(N11686,N12819,N12833);
or or1079(N11687,N12847,N12861);
or or1080(N11688,N12875,N12889);
or or1081(N11689,N12903,N12917);
or or1082(N11690,N12931,N12945);
or or1083(N11691,N12959,N12973);
or or1084(N11692,N12987,N13001);
or or1085(N11693,N13015,N13029);
or or1086(N11694,N13043,N13057);
or or1087(N11695,N13071,N13085);
or or1088(N11696,N13099,N13113);
or or1089(N11697,N13127,N13141);
or or1090(N11698,N13155,N13169);
or or1091(N11699,N13183,N13197);
or or1092(N11700,N13211,N13225);
or or1093(N11701,N13239,N13253);
or or1094(N11702,N13267,N13281);
or or1095(N11703,N13295,N13309);
or or1096(N11704,N13323,N13336);
or or1097(N11705,N13349,N13362);
or or1098(N11706,N13375,N13388);
or or1099(N11707,N13401,N13414);
or or1100(N11708,N13427,N13440);
or or1101(N11709,N13453,N13466);
or or1102(N11710,N13479,N13492);
or or1103(N11711,N13505,N13518);
or or1104(N11712,N13531,N13544);
or or1105(N11713,N13557,N13570);
or or1106(N11714,N13583,N13596);
or or1107(N11715,N13609,N13622);
or or1108(N11716,N13635,N13648);
or or1109(N11717,N13661,N13674);
or or1110(N11718,N13687,N13700);
or or1111(N11719,N13713,N13726);
or or1112(N11720,N13739,N13752);
or or1113(N11721,N13765,N13778);
or or1114(N11722,N13791,N13804);
or or1115(N11723,N13817,N13830);
or or1116(N11724,N13843,N13856);
or or1117(N11725,N13869,N13882);
or or1118(N11726,N13895,N13908);
or or1119(N11727,N13921,N13933);
or or1120(N11728,N13945,N13957);
or or1121(N11729,N13969,N13981);
or or1122(N11730,N13993,N14005);
or or1123(N11731,N14017,N14029);
or or1124(N11732,N14041,N14053);
or or1125(N11733,N14065,N14077);
or or1126(N11734,N14089,N14101);
or or1127(N11735,N14113,N14125);
or or1128(N11736,N14137,N14149);
or or1129(N11737,N14161,N14173);
or or1130(N11738,N14185,N14197);
or or1131(N11739,N14209,N14221);
or or1132(N11740,N14233,N14245);
or or1133(N11741,N14257,N14268);
or or1134(N11742,N14279,N14290);
or or1135(N11743,N14301,N14312);
or or1136(N11744,N14323,N14334);
or or1137(N11745,N14345,N14356);
or or1138(N11746,N14367,N14378);
or or1139(N11747,N14389,N14400);
or or1140(N11748,N14411,N14422);
or or1141(N11749,N14433,N14443);
or or1142(N11750,N14453,N14463);
or or1143(N11751,N14473,N14483);
or or1144(N11752,N14493,N14502);
or or1145(N11753,N14518,N14534);
or or1146(N11754,N14550,N14565);
or or1147(N11755,N14580,N14595);
or or1148(N11756,N14610,N14625);
or or1149(N11757,N14640,N14655);
or or1150(N11758,N14670,N14685);
or or1151(N11759,N14700,N14714);
or or1152(N11760,N14728,N14742);
or or1153(N11761,N14756,N14770);
or or1154(N11762,N14784,N14798);
or or1155(N11763,N14812,N14826);
or or1156(N11764,N14840,N14854);
or or1157(N11765,N14868,N14882);
or or1158(N11766,N14896,N14910);
or or1159(N11767,N14924,N14938);
or or1160(N11768,N14952,N14966);
or or1161(N11769,N14980,N14994);
or or1162(N11770,N15008,N15022);
or or1163(N11771,N15036,N15050);
or or1164(N11772,N15064,N15078);
or or1165(N11773,N15092,N15106);
or or1166(N11774,N15120,N15134);
or or1167(N11775,N15148,N15162);
or or1168(N11776,N15176,N15190);
or or1169(N11777,N15203,N15216);
or or1170(N11778,N15229,N15242);
or or1171(N11779,N15255,N15268);
or or1172(N11780,N15281,N15294);
or or1173(N11781,N15307,N15320);
or or1174(N11782,N15333,N15346);
or or1175(N11783,N15359,N15372);
or or1176(N11784,N15385,N15398);
or or1177(N11785,N15411,N15424);
or or1178(N11786,N15437,N15450);
or or1179(N11787,N15463,N15476);
or or1180(N11788,N15489,N15502);
or or1181(N11789,N15515,N15528);
or or1182(N11790,N15541,N15554);
or or1183(N11791,N15567,N15580);
or or1184(N11792,N15593,N15606);
or or1185(N11793,N15619,N15632);
or or1186(N11794,N15645,N15658);
or or1187(N11795,N15671,N15684);
or or1188(N11796,N15697,N15710);
or or1189(N11797,N15723,N15736);
or or1190(N11798,N15749,N15762);
or or1191(N11799,N15775,N15788);
or or1192(N11800,N15801,N15814);
or or1193(N11801,N15826,N15838);
or or1194(N11802,N15850,N15862);
or or1195(N11803,N15874,N15886);
or or1196(N11804,N15898,N15910);
or or1197(N11805,N15922,N15934);
or or1198(N11806,N15946,N15958);
or or1199(N11807,N15970,N15982);
or or1200(N11808,N15994,N16006);
or or1201(N11809,N16018,N16030);
or or1202(N11810,N16042,N16054);
or or1203(N11811,N16066,N16078);
or or1204(N11812,N16090,N16102);
or or1205(N11813,N16114,N16126);
or or1206(N11814,N16138,N16150);
or or1207(N11815,N16162,N16174);
or or1208(N11816,N16186,N16198);
or or1209(N11817,N16210,N16222);
or or1210(N11818,N16234,N16246);
or or1211(N11819,N16258,N16270);
or or1212(N11820,N16282,N16294);
or or1213(N11821,N16306,N16318);
or or1214(N11822,N16330,N16342);
or or1215(N11823,N16354,N16366);
or or1216(N11824,N16378,N16390);
or or1217(N11825,N16402,N16414);
or or1218(N11826,N16426,N16438);
or or1219(N11827,N16450,N16461);
or or1220(N11828,N16472,N16483);
or or1221(N11829,N16494,N16505);
or or1222(N11830,N16516,N16527);
or or1223(N11831,N16538,N16549);
or or1224(N11832,N16560,N16571);
or or1225(N11833,N16582,N16593);
or or1226(N11834,N16604,N16615);
or or1227(N11835,N16626,N16637);
or or1228(N11836,N16648,N16659);
or or1229(N11837,N16670,N16681);
or or1230(N11838,N16692,N16703);
or or1231(N11839,N16714,N16725);
or or1232(N11840,N16736,N16747);
or or1233(N11841,N16758,N16769);
or or1234(N11842,N16780,N16791);
or or1235(N11843,N16802,N16813);
or or1236(N11844,N16824,N16835);
or or1237(N11845,N16846,N16857);
or or1238(N11846,N16868,N16879);
or or1239(N11847,N16890,N16900);
or or1240(N11848,N16910,N16920);
or or1241(N11849,N16930,N16940);
or or1242(N11850,N16950,N16960);
or or1243(N11851,N16970,N16980);
or or1244(N11852,N16990,N17000);
or or1245(N11853,N17010,N17020);
or or1246(N11854,N17030,N17040);
or or1247(N11855,N17050,N17060);
or or1248(N11856,N17069,N17078);
or or1249(N11857,N17087,N17096);
or or1250(N11858,N17105,N17114);
or or1251(N11859,N17123,N17132);
or or1252(N11860,N17141,N17150);
or or1253(N11861,N17158,N17172);
or or1254(N11862,N17186,N17200);
or or1255(N11863,N17214,N17227);
or or1256(N11864,N17240,N17253);
or or1257(N11865,N17266,N17279);
or or1258(N11866,N17291,N17303);
or or1259(N11867,N17315,N17327);
or or1260(N11868,N17339,N17351);
or or1261(N11869,N17363,N17375);
or or1262(N11870,N17387,N17398);
or or1263(N11871,N17409,N17420);
or or1264(N11872,N17431,N17442);
or or1265(N11873,N17453,N17464);
or or1266(N11874,N17475,N17486);
or or1267(N11875,N17497,N17508);
or or1268(N11876,N17519,N17530);
or or1269(N11877,N17541,N17552);
or or1270(N11878,N17563,N17574);
or or1271(N11879,N17584,N17594);
or or1272(N11880,N17604,N17614);
or or1273(N11881,N17624,N17634);
or or1274(N17644,N17645,N17646);
or or1275(N17645,N17647,N17648);
or or1276(N17646,N17649,N17650);
or or1277(N17647,N17651,N17652);
or or1278(N17648,N17653,N17654);
or or1279(N17649,N17655,N17656);
or or1280(N17650,N17657,N17658);
or or1281(N17651,N17659,N17660);
or or1282(N17652,N17661,N17662);
or or1283(N17653,N17663,N17664);
or or1284(N17654,N17665,N17666);
or or1285(N17655,N17667,N17668);
or or1286(N17656,N17669,N17670);
or or1287(N17657,N17671,N17672);
or or1288(N17658,N17673,N17674);
or or1289(N17659,N17675,N17676);
or or1290(N17660,N17677,N17678);
or or1291(N17661,N17679,N17680);
or or1292(N17662,N17681,N17682);
or or1293(N17663,N17683,N17684);
or or1294(N17664,N17685,N17686);
or or1295(N17665,N17687,N17688);
or or1296(N17666,N17689,N17690);
or or1297(N17667,N17691,N17692);
or or1298(N17668,N17693,N17694);
or or1299(N17669,N17695,N17696);
or or1300(N17670,N17697,N17698);
or or1301(N17671,N17699,N17700);
or or1302(N17672,N17701,N17702);
or or1303(N17673,N17703,N17704);
or or1304(N17674,N17705,N17706);
or or1305(N17675,N17707,N17708);
or or1306(N17676,N17709,N17710);
or or1307(N17677,N17711,N17712);
or or1308(N17678,N17713,N17714);
or or1309(N17679,N17715,N17716);
or or1310(N17680,N17717,N17718);
or or1311(N17681,N17719,N17720);
or or1312(N17682,N17721,N17722);
or or1313(N17683,N17723,N17724);
or or1314(N17684,N17725,N17726);
or or1315(N17685,N17727,N17728);
or or1316(N17686,N17729,N17730);
or or1317(N17687,N17731,N17732);
or or1318(N17688,N17733,N17734);
or or1319(N17689,N17735,N17736);
or or1320(N17690,N17737,N17738);
or or1321(N17691,N17739,N17740);
or or1322(N17692,N17741,N17742);
or or1323(N17693,N17743,N17744);
or or1324(N17694,N17745,N17746);
or or1325(N17695,N17747,N17748);
or or1326(N17696,N17749,N17750);
or or1327(N17697,N17751,N17752);
or or1328(N17698,N17753,N17754);
or or1329(N17699,N17755,N17756);
or or1330(N17700,N17757,N17758);
or or1331(N17701,N17759,N17760);
or or1332(N17702,N17761,N17762);
or or1333(N17703,N17763,N17764);
or or1334(N17704,N17765,N17766);
or or1335(N17705,N17767,N17768);
or or1336(N17706,N17769,N17770);
or or1337(N17707,N17771,N17772);
or or1338(N17708,N17773,N17774);
or or1339(N17709,N17775,N17776);
or or1340(N17710,N17777,N17778);
or or1341(N17711,N17779,N17780);
or or1342(N17712,N17781,N17782);
or or1343(N17713,N17783,N17784);
or or1344(N17714,N17785,N17786);
or or1345(N17715,N17787,N17788);
or or1346(N17716,N17789,N17790);
or or1347(N17717,N17791,N17792);
or or1348(N17718,N17793,N17794);
or or1349(N17719,N17795,N17796);
or or1350(N17720,N17797,N17798);
or or1351(N17721,N17799,N17800);
or or1352(N17722,N17801,N17802);
or or1353(N17723,N17803,N17804);
or or1354(N17724,N17805,N17806);
or or1355(N17725,N17807,N17808);
or or1356(N17726,N17809,N17810);
or or1357(N17727,N17811,N17812);
or or1358(N17728,N17813,N17814);
or or1359(N17729,N17815,N17816);
or or1360(N17730,N17817,N17818);
or or1361(N17731,N17819,N17820);
or or1362(N17732,N17821,N17822);
or or1363(N17733,N17823,N17824);
or or1364(N17734,N17825,N17826);
or or1365(N17735,N17827,N17828);
or or1366(N17736,N17829,N17830);
or or1367(N17737,N17831,N17832);
or or1368(N17738,N17833,N17834);
or or1369(N17739,N17835,N17836);
or or1370(N17740,N17837,N17838);
or or1371(N17741,N17839,N17840);
or or1372(N17742,N17841,N17842);
or or1373(N17743,N17843,N17844);
or or1374(N17744,N17845,N17846);
or or1375(N17745,N17847,N17848);
or or1376(N17746,N17849,N17850);
or or1377(N17747,N17851,N17852);
or or1378(N17748,N17853,N17854);
or or1379(N17749,N17855,N17856);
or or1380(N17750,N17857,N17858);
or or1381(N17751,N17859,N17860);
or or1382(N17752,N17861,N17862);
or or1383(N17753,N17863,N17864);
or or1384(N17754,N17865,N17866);
or or1385(N17755,N17867,N17868);
or or1386(N17756,N17869,N17870);
or or1387(N17757,N17871,N17872);
or or1388(N17758,N17873,N17874);
or or1389(N17759,N17875,N17876);
or or1390(N17760,N17877,N17878);
or or1391(N17761,N17879,N17880);
or or1392(N17762,N17881,N17882);
or or1393(N17763,N17883,N17884);
or or1394(N17764,N17885,N17886);
or or1395(N17765,N17887,N17888);
or or1396(N17766,N17889,N17890);
or or1397(N17767,N17891,N17892);
or or1398(N17768,N17893,N17894);
or or1399(N17769,N17895,N17896);
or or1400(N17770,N17897,N17898);
or or1401(N17771,N17899,N17900);
or or1402(N17772,N17901,N17902);
or or1403(N17773,N17903,N17904);
or or1404(N17774,N17905,N17906);
or or1405(N17775,N17907,N17908);
or or1406(N17776,N17909,N17910);
or or1407(N17777,N17911,N17912);
or or1408(N17778,N17913,N17914);
or or1409(N17779,N17915,N17916);
or or1410(N17780,N17917,N17918);
or or1411(N17781,N17919,N17920);
or or1412(N17782,N17921,N17922);
or or1413(N17783,N17923,N17924);
or or1414(N17784,N17925,N17926);
or or1415(N17785,N17927,N17928);
or or1416(N17786,N17929,N17930);
or or1417(N17787,N17931,N17932);
or or1418(N17788,N17933,N17934);
or or1419(N17789,N17935,N17936);
or or1420(N17790,N17937,N17938);
or or1421(N17791,N17939,N17940);
or or1422(N17792,N17941,N17942);
or or1423(N17793,N17943,N17944);
or or1424(N17794,N17945,N17946);
or or1425(N17795,N17947,N17948);
or or1426(N17796,N17949,N17950);
or or1427(N17797,N17951,N17952);
or or1428(N17798,N17953,N17954);
or or1429(N17799,N17955,N17956);
or or1430(N17800,N17957,N17958);
or or1431(N17801,N17959,N17960);
or or1432(N17802,N17961,N17962);
or or1433(N17803,N17963,N17964);
or or1434(N17804,N17965,N17966);
or or1435(N17805,N17967,N17968);
or or1436(N17806,N17969,N17970);
or or1437(N17807,N17971,N17972);
or or1438(N17808,N17973,N17974);
or or1439(N17809,N17975,N17976);
or or1440(N17810,N17977,N17978);
or or1441(N17811,N17979,N17980);
or or1442(N17812,N17981,N17982);
or or1443(N17813,N17983,N17984);
or or1444(N17814,N17985,N17986);
or or1445(N17815,N17987,N17988);
or or1446(N17816,N17989,N17990);
or or1447(N17817,N17991,N17992);
or or1448(N17818,N17993,N17994);
or or1449(N17819,N17995,N17996);
or or1450(N17820,N17997,N17998);
or or1451(N17821,N17999,N18000);
or or1452(N17822,N18001,N18002);
or or1453(N17823,N18003,N18004);
or or1454(N17824,N18005,N18006);
or or1455(N17825,N18007,N18008);
or or1456(N17826,N18009,N18010);
or or1457(N17827,N18011,N18012);
or or1458(N17828,N18013,N18014);
or or1459(N17829,N18015,N18016);
or or1460(N17830,N18017,N18018);
or or1461(N17831,N18019,N18020);
or or1462(N17832,N18021,N18022);
or or1463(N17833,N18023,N18024);
or or1464(N17834,N18025,N18026);
or or1465(N17835,N18027,N18028);
or or1466(N17836,N18029,N18030);
or or1467(N17837,N18031,N18032);
or or1468(N17838,N18033,N18034);
or or1469(N17839,N18035,N18036);
or or1470(N17840,N18037,N18038);
or or1471(N17841,N18039,N18040);
or or1472(N17842,N18041,N18042);
or or1473(N17843,N18043,N18044);
or or1474(N17844,N18045,N18046);
or or1475(N17845,N18047,N18048);
or or1476(N17846,N18049,N18050);
or or1477(N17847,N18051,N18052);
or or1478(N17848,N18053,N18054);
or or1479(N17849,N18055,N18056);
or or1480(N17850,N18057,N18058);
or or1481(N17851,N18059,N18060);
or or1482(N17852,N18061,N18062);
or or1483(N17853,N18063,N18064);
or or1484(N17854,N18065,N18066);
or or1485(N17855,N18067,N18068);
or or1486(N17856,N18069,N18070);
or or1487(N17857,N18071,N18072);
or or1488(N17858,N18073,N18074);
or or1489(N17859,N18075,N18076);
or or1490(N17860,N18077,N18078);
or or1491(N17861,N18079,N18080);
or or1492(N17862,N18081,N18082);
or or1493(N17863,N18083,N18084);
or or1494(N17864,N18085,N18086);
or or1495(N17865,N18087,N18088);
or or1496(N17866,N18089,N18090);
or or1497(N17867,N18091,N18092);
or or1498(N17868,N18093,N18094);
or or1499(N17869,N18095,N18096);
or or1500(N17870,N18097,N18098);
or or1501(N17871,N18099,N18100);
or or1502(N17872,N18101,N18102);
or or1503(N17873,N18103,N18104);
or or1504(N17874,N18105,N18106);
or or1505(N17875,N18107,N18108);
or or1506(N17876,N18109,N18110);
or or1507(N17877,N18128,N18145);
or or1508(N17878,N18162,N18179);
or or1509(N17879,N18196,N18213);
or or1510(N17880,N18230,N18246);
or or1511(N17881,N18262,N18278);
or or1512(N17882,N18294,N18310);
or or1513(N17883,N18326,N18342);
or or1514(N17884,N18358,N18374);
or or1515(N17885,N18390,N18406);
or or1516(N17886,N18422,N18438);
or or1517(N17887,N18454,N18470);
or or1518(N17888,N18486,N18502);
or or1519(N17889,N18518,N18534);
or or1520(N17890,N18550,N18565);
or or1521(N17891,N18580,N18595);
or or1522(N17892,N18610,N18625);
or or1523(N17893,N18640,N18655);
or or1524(N17894,N18670,N18685);
or or1525(N17895,N18700,N18715);
or or1526(N17896,N18730,N18745);
or or1527(N17897,N18760,N18775);
or or1528(N17898,N18790,N18805);
or or1529(N17899,N18820,N18835);
or or1530(N17900,N18850,N18865);
or or1531(N17901,N18880,N18895);
or or1532(N17902,N18910,N18924);
or or1533(N17903,N18938,N18952);
or or1534(N17904,N18966,N18980);
or or1535(N17905,N18994,N19008);
or or1536(N17906,N19022,N19036);
or or1537(N17907,N19050,N19064);
or or1538(N17908,N19078,N19092);
or or1539(N17909,N19106,N19120);
or or1540(N17910,N19134,N19148);
or or1541(N17911,N19162,N19176);
or or1542(N17912,N19190,N19204);
or or1543(N17913,N19218,N19232);
or or1544(N17914,N19246,N19260);
or or1545(N17915,N19274,N19288);
or or1546(N17916,N19302,N19316);
or or1547(N17917,N19330,N19344);
or or1548(N17918,N19358,N19372);
or or1549(N17919,N19386,N19400);
or or1550(N17920,N19414,N19428);
or or1551(N17921,N19442,N19456);
or or1552(N17922,N19470,N19484);
or or1553(N17923,N19498,N19512);
or or1554(N17924,N19526,N19540);
or or1555(N17925,N19554,N19568);
or or1556(N17926,N19582,N19596);
or or1557(N17927,N19610,N19624);
or or1558(N17928,N19638,N19652);
or or1559(N17929,N19666,N19680);
or or1560(N17930,N19694,N19708);
or or1561(N17931,N19722,N19735);
or or1562(N17932,N19748,N19761);
or or1563(N17933,N19774,N19787);
or or1564(N17934,N19800,N19813);
or or1565(N17935,N19826,N19839);
or or1566(N17936,N19852,N19865);
or or1567(N17937,N19878,N19891);
or or1568(N17938,N19904,N19917);
or or1569(N17939,N19930,N19943);
or or1570(N17940,N19956,N19969);
or or1571(N17941,N19982,N19995);
or or1572(N17942,N20008,N20021);
or or1573(N17943,N20034,N20047);
or or1574(N17944,N20060,N20073);
or or1575(N17945,N20086,N20099);
or or1576(N17946,N20112,N20125);
or or1577(N17947,N20138,N20151);
or or1578(N17948,N20164,N20177);
or or1579(N17949,N20190,N20203);
or or1580(N17950,N20216,N20229);
or or1581(N17951,N20242,N20254);
or or1582(N17952,N20266,N20278);
or or1583(N17953,N20290,N20302);
or or1584(N17954,N20314,N20326);
or or1585(N17955,N20338,N20350);
or or1586(N17956,N20362,N20374);
or or1587(N17957,N20386,N20398);
or or1588(N17958,N20410,N20422);
or or1589(N17959,N20434,N20446);
or or1590(N17960,N20458,N20470);
or or1591(N17961,N20482,N20494);
or or1592(N17962,N20506,N20518);
or or1593(N17963,N20530,N20542);
or or1594(N17964,N20554,N20566);
or or1595(N17965,N20578,N20590);
or or1596(N17966,N20602,N20614);
or or1597(N17967,N20626,N20638);
or or1598(N17968,N20650,N20662);
or or1599(N17969,N20673,N20684);
or or1600(N17970,N20695,N20706);
or or1601(N17971,N20717,N20728);
or or1602(N17972,N20738,N20748);
or or1603(N17973,N20758,N20768);
or or1604(N17974,N20778,N20788);
or or1605(N17975,N20798,N20808);
or or1606(N17976,N20818,N20828);
or or1607(N17977,N20838,N20848);
or or1608(N17978,N20864,N20880);
or or1609(N17979,N20895,N20910);
or or1610(N17980,N20925,N20940);
or or1611(N17981,N20955,N20970);
or or1612(N17982,N20985,N21000);
or or1613(N17983,N21015,N21030);
or or1614(N17984,N21045,N21060);
or or1615(N17985,N21075,N21089);
or or1616(N17986,N21103,N21117);
or or1617(N17987,N21131,N21145);
or or1618(N17988,N21159,N21173);
or or1619(N17989,N21187,N21201);
or or1620(N17990,N21215,N21229);
or or1621(N17991,N21243,N21257);
or or1622(N17992,N21271,N21285);
or or1623(N17993,N21299,N21313);
or or1624(N17994,N21327,N21341);
or or1625(N17995,N21355,N21369);
or or1626(N17996,N21383,N21397);
or or1627(N17997,N21411,N21425);
or or1628(N17998,N21439,N21453);
or or1629(N17999,N21467,N21481);
or or1630(N18000,N21495,N21509);
or or1631(N18001,N21523,N21536);
or or1632(N18002,N21549,N21562);
or or1633(N18003,N21575,N21588);
or or1634(N18004,N21601,N21614);
or or1635(N18005,N21627,N21640);
or or1636(N18006,N21653,N21666);
or or1637(N18007,N21679,N21692);
or or1638(N18008,N21705,N21718);
or or1639(N18009,N21731,N21744);
or or1640(N18010,N21757,N21770);
or or1641(N18011,N21783,N21796);
or or1642(N18012,N21809,N21822);
or or1643(N18013,N21835,N21848);
or or1644(N18014,N21861,N21874);
or or1645(N18015,N21887,N21900);
or or1646(N18016,N21913,N21926);
or or1647(N18017,N21939,N21952);
or or1648(N18018,N21965,N21978);
or or1649(N18019,N21991,N22004);
or or1650(N18020,N22017,N22030);
or or1651(N18021,N22043,N22056);
or or1652(N18022,N22069,N22082);
or or1653(N18023,N22095,N22108);
or or1654(N18024,N22121,N22134);
or or1655(N18025,N22147,N22160);
or or1656(N18026,N22173,N22186);
or or1657(N18027,N22199,N22212);
or or1658(N18028,N22225,N22237);
or or1659(N18029,N22249,N22261);
or or1660(N18030,N22273,N22285);
or or1661(N18031,N22297,N22309);
or or1662(N18032,N22321,N22333);
or or1663(N18033,N22345,N22357);
or or1664(N18034,N22369,N22381);
or or1665(N18035,N22393,N22405);
or or1666(N18036,N22417,N22429);
or or1667(N18037,N22441,N22453);
or or1668(N18038,N22465,N22477);
or or1669(N18039,N22489,N22501);
or or1670(N18040,N22513,N22525);
or or1671(N18041,N22537,N22549);
or or1672(N18042,N22561,N22573);
or or1673(N18043,N22585,N22597);
or or1674(N18044,N22609,N22621);
or or1675(N18045,N22633,N22645);
or or1676(N18046,N22657,N22669);
or or1677(N18047,N22681,N22693);
or or1678(N18048,N22705,N22717);
or or1679(N18049,N22729,N22741);
or or1680(N18050,N22753,N22765);
or or1681(N18051,N22777,N22789);
or or1682(N18052,N22801,N22813);
or or1683(N18053,N22825,N22836);
or or1684(N18054,N22847,N22858);
or or1685(N18055,N22869,N22880);
or or1686(N18056,N22891,N22902);
or or1687(N18057,N22913,N22924);
or or1688(N18058,N22935,N22946);
or or1689(N18059,N22957,N22968);
or or1690(N18060,N22979,N22990);
or or1691(N18061,N23001,N23012);
or or1692(N18062,N23023,N23034);
or or1693(N18063,N23045,N23056);
or or1694(N18064,N23067,N23078);
or or1695(N18065,N23089,N23100);
or or1696(N18066,N23111,N23122);
or or1697(N18067,N23133,N23144);
or or1698(N18068,N23155,N23166);
or or1699(N18069,N23177,N23188);
or or1700(N18070,N23199,N23210);
or or1701(N18071,N23221,N23232);
or or1702(N18072,N23243,N23254);
or or1703(N18073,N23265,N23276);
or or1704(N18074,N23287,N23298);
or or1705(N18075,N23309,N23320);
or or1706(N18076,N23331,N23342);
or or1707(N18077,N23353,N23364);
or or1708(N18078,N23375,N23386);
or or1709(N18079,N23397,N23407);
or or1710(N18080,N23417,N23427);
or or1711(N18081,N23437,N23447);
or or1712(N18082,N23457,N23467);
or or1713(N18083,N23477,N23487);
or or1714(N18084,N23497,N23507);
or or1715(N18085,N23517,N23527);
or or1716(N18086,N23537,N23547);
or or1717(N18087,N23556,N23565);
or or1718(N18088,N23574,N23583);
or or1719(N18089,N23592,N23601);
or or1720(N18090,N23610,N23619);
or or1721(N18091,N23628,N23636);
or or1722(N18092,N23650,N23664);
or or1723(N18093,N23677,N23690);
or or1724(N18094,N23703,N23716);
or or1725(N18095,N23729,N23742);
or or1726(N18096,N23754,N23766);
or or1727(N18097,N23778,N23790);
or or1728(N18098,N23802,N23814);
or or1729(N18099,N23826,N23838);
or or1730(N18100,N23850,N23861);
or or1731(N18101,N23872,N23883);
or or1732(N18102,N23894,N23905);
or or1733(N18103,N23916,N23927);
or or1734(N18104,N23938,N23948);
or or1735(N18105,N23958,N23968);
or or1736(N18106,N23978,N23988);
or or1737(N18107,N23998,N24008);
or or1738(N18108,N24018,N24028);
or or1739(N18109,N24038,N24047);
or or1740(N24056,N24057,N24058);
or or1741(N24057,N24059,N24060);
or or1742(N24058,N24061,N24062);
or or1743(N24059,N24063,N24064);
or or1744(N24060,N24065,N24066);
or or1745(N24061,N24067,N24068);
or or1746(N24062,N24069,N24070);
or or1747(N24063,N24071,N24072);
or or1748(N24064,N24073,N24074);
or or1749(N24065,N24075,N24076);
or or1750(N24066,N24077,N24078);
or or1751(N24067,N24079,N24080);
or or1752(N24068,N24081,N24082);
or or1753(N24069,N24083,N24084);
or or1754(N24070,N24085,N24086);
or or1755(N24071,N24087,N24088);
or or1756(N24072,N24089,N24090);
or or1757(N24073,N24091,N24092);
or or1758(N24074,N24093,N24094);
or or1759(N24075,N24095,N24096);
or or1760(N24076,N24097,N24098);
or or1761(N24077,N24099,N24100);
or or1762(N24078,N24101,N24102);
or or1763(N24079,N24103,N24104);
or or1764(N24080,N24105,N24106);
or or1765(N24081,N24107,N24108);
or or1766(N24082,N24109,N24110);
or or1767(N24083,N24111,N24112);
or or1768(N24084,N24113,N24114);
or or1769(N24085,N24115,N24116);
or or1770(N24086,N24117,N24118);
or or1771(N24087,N24119,N24120);
or or1772(N24088,N24121,N24122);
or or1773(N24089,N24123,N24124);
or or1774(N24090,N24125,N24126);
or or1775(N24091,N24127,N24128);
or or1776(N24092,N24129,N24130);
or or1777(N24093,N24131,N24132);
or or1778(N24094,N24133,N24134);
or or1779(N24095,N24135,N24136);
or or1780(N24096,N24137,N24138);
or or1781(N24097,N24139,N24140);
or or1782(N24098,N24141,N24142);
or or1783(N24099,N24143,N24144);
or or1784(N24100,N24145,N24146);
or or1785(N24101,N24147,N24148);
or or1786(N24102,N24149,N24150);
or or1787(N24103,N24151,N24152);
or or1788(N24104,N24153,N24154);
or or1789(N24105,N24155,N24156);
or or1790(N24106,N24157,N24158);
or or1791(N24107,N24159,N24160);
or or1792(N24108,N24161,N24162);
or or1793(N24109,N24163,N24164);
or or1794(N24110,N24165,N24166);
or or1795(N24111,N24167,N24168);
or or1796(N24112,N24169,N24170);
or or1797(N24113,N24171,N24172);
or or1798(N24114,N24173,N24174);
or or1799(N24115,N24175,N24176);
or or1800(N24116,N24177,N24178);
or or1801(N24117,N24179,N24180);
or or1802(N24118,N24181,N24182);
or or1803(N24119,N24183,N24184);
or or1804(N24120,N24185,N24186);
or or1805(N24121,N24187,N24188);
or or1806(N24122,N24189,N24190);
or or1807(N24123,N24191,N24192);
or or1808(N24124,N24193,N24194);
or or1809(N24125,N24195,N24196);
or or1810(N24126,N24197,N24198);
or or1811(N24127,N24199,N24200);
or or1812(N24128,N24201,N24202);
or or1813(N24129,N24203,N24204);
or or1814(N24130,N24205,N24206);
or or1815(N24131,N24207,N24208);
or or1816(N24132,N24209,N24210);
or or1817(N24133,N24211,N24212);
or or1818(N24134,N24213,N24214);
or or1819(N24135,N24215,N24216);
or or1820(N24136,N24217,N24218);
or or1821(N24137,N24219,N24220);
or or1822(N24138,N24221,N24222);
or or1823(N24139,N24223,N24224);
or or1824(N24140,N24225,N24226);
or or1825(N24141,N24227,N24228);
or or1826(N24142,N24229,N24230);
or or1827(N24143,N24231,N24232);
or or1828(N24144,N24233,N24234);
or or1829(N24145,N24235,N24236);
or or1830(N24146,N24237,N24238);
or or1831(N24147,N24239,N24240);
or or1832(N24148,N24241,N24242);
or or1833(N24149,N24243,N24244);
or or1834(N24150,N24245,N24246);
or or1835(N24151,N24247,N24248);
or or1836(N24152,N24249,N24250);
or or1837(N24153,N24251,N24252);
or or1838(N24154,N24253,N24254);
or or1839(N24155,N24255,N24256);
or or1840(N24156,N24257,N24258);
or or1841(N24157,N24259,N24260);
or or1842(N24158,N24261,N24262);
or or1843(N24159,N24263,N24264);
or or1844(N24160,N24265,N24266);
or or1845(N24161,N24267,N24268);
or or1846(N24162,N24269,N24270);
or or1847(N24163,N24271,N24272);
or or1848(N24164,N24273,N24274);
or or1849(N24165,N24275,N24276);
or or1850(N24166,N24277,N24278);
or or1851(N24167,N24279,N24280);
or or1852(N24168,N24281,N24282);
or or1853(N24169,N24283,N24284);
or or1854(N24170,N24285,N24286);
or or1855(N24171,N24287,N24288);
or or1856(N24172,N24289,N24290);
or or1857(N24173,N24291,N24292);
or or1858(N24174,N24293,N24294);
or or1859(N24175,N24295,N24296);
or or1860(N24176,N24297,N24298);
or or1861(N24177,N24299,N24300);
or or1862(N24178,N24301,N24302);
or or1863(N24179,N24303,N24304);
or or1864(N24180,N24305,N24306);
or or1865(N24181,N24307,N24308);
or or1866(N24182,N24309,N24310);
or or1867(N24183,N24311,N24312);
or or1868(N24184,N24313,N24314);
or or1869(N24185,N24315,N24316);
or or1870(N24186,N24317,N24318);
or or1871(N24187,N24319,N24320);
or or1872(N24188,N24321,N24322);
or or1873(N24189,N24323,N24324);
or or1874(N24190,N24325,N24326);
or or1875(N24191,N24327,N24328);
or or1876(N24192,N24329,N24330);
or or1877(N24193,N24331,N24332);
or or1878(N24194,N24333,N24334);
or or1879(N24195,N24335,N24336);
or or1880(N24196,N24337,N24338);
or or1881(N24197,N24339,N24340);
or or1882(N24198,N24341,N24342);
or or1883(N24199,N24343,N24344);
or or1884(N24200,N24345,N24346);
or or1885(N24201,N24347,N24348);
or or1886(N24202,N24349,N24350);
or or1887(N24203,N24351,N24352);
or or1888(N24204,N24353,N24354);
or or1889(N24205,N24355,N24356);
or or1890(N24206,N24357,N24358);
or or1891(N24207,N24359,N24360);
or or1892(N24208,N24361,N24362);
or or1893(N24209,N24363,N24364);
or or1894(N24210,N24365,N24366);
or or1895(N24211,N24367,N24368);
or or1896(N24212,N24369,N24370);
or or1897(N24213,N24371,N24372);
or or1898(N24214,N24373,N24374);
or or1899(N24215,N24375,N24376);
or or1900(N24216,N24377,N24378);
or or1901(N24217,N24379,N24380);
or or1902(N24218,N24381,N24382);
or or1903(N24219,N24383,N24384);
or or1904(N24220,N24385,N24386);
or or1905(N24221,N24387,N24388);
or or1906(N24222,N24389,N24390);
or or1907(N24223,N24391,N24392);
or or1908(N24224,N24393,N24394);
or or1909(N24225,N24395,N24396);
or or1910(N24226,N24397,N24398);
or or1911(N24227,N24399,N24400);
or or1912(N24228,N24401,N24402);
or or1913(N24229,N24403,N24404);
or or1914(N24230,N24405,N24406);
or or1915(N24231,N24407,N24408);
or or1916(N24232,N24409,N24410);
or or1917(N24233,N24411,N24412);
or or1918(N24234,N24413,N24414);
or or1919(N24235,N24415,N24416);
or or1920(N24236,N24417,N24418);
or or1921(N24237,N24419,N24420);
or or1922(N24238,N24421,N24422);
or or1923(N24239,N24423,N24424);
or or1924(N24240,N24425,N24426);
or or1925(N24241,N24427,N24444);
or or1926(N24242,N24461,N24478);
or or1927(N24243,N24495,N24512);
or or1928(N24244,N24529,N24546);
or or1929(N24245,N24563,N24579);
or or1930(N24246,N24595,N24611);
or or1931(N24247,N24627,N24643);
or or1932(N24248,N24659,N24675);
or or1933(N24249,N24691,N24707);
or or1934(N24250,N24723,N24739);
or or1935(N24251,N24755,N24771);
or or1936(N24252,N24787,N24803);
or or1937(N24253,N24819,N24835);
or or1938(N24254,N24851,N24867);
or or1939(N24255,N24882,N24897);
or or1940(N24256,N24912,N24927);
or or1941(N24257,N24942,N24957);
or or1942(N24258,N24972,N24987);
or or1943(N24259,N25002,N25017);
or or1944(N24260,N25032,N25047);
or or1945(N24261,N25062,N25077);
or or1946(N24262,N25092,N25107);
or or1947(N24263,N25122,N25137);
or or1948(N24264,N25152,N25167);
or or1949(N24265,N25182,N25197);
or or1950(N24266,N25212,N25227);
or or1951(N24267,N25242,N25257);
or or1952(N24268,N25271,N25285);
or or1953(N24269,N25299,N25313);
or or1954(N24270,N25327,N25341);
or or1955(N24271,N25355,N25369);
or or1956(N24272,N25383,N25397);
or or1957(N24273,N25411,N25425);
or or1958(N24274,N25439,N25453);
or or1959(N24275,N25467,N25481);
or or1960(N24276,N25495,N25509);
or or1961(N24277,N25523,N25537);
or or1962(N24278,N25551,N25565);
or or1963(N24279,N25579,N25593);
or or1964(N24280,N25607,N25621);
or or1965(N24281,N25635,N25649);
or or1966(N24282,N25663,N25677);
or or1967(N24283,N25691,N25705);
or or1968(N24284,N25719,N25733);
or or1969(N24285,N25747,N25761);
or or1970(N24286,N25775,N25789);
or or1971(N24287,N25803,N25817);
or or1972(N24288,N25831,N25845);
or or1973(N24289,N25859,N25873);
or or1974(N24290,N25887,N25901);
or or1975(N24291,N25915,N25929);
or or1976(N24292,N25943,N25957);
or or1977(N24293,N25971,N25985);
or or1978(N24294,N25999,N26013);
or or1979(N24295,N26027,N26041);
or or1980(N24296,N26055,N26069);
or or1981(N24297,N26083,N26097);
or or1982(N24298,N26111,N26125);
or or1983(N24299,N26139,N26152);
or or1984(N24300,N26165,N26178);
or or1985(N24301,N26191,N26204);
or or1986(N24302,N26217,N26230);
or or1987(N24303,N26243,N26256);
or or1988(N24304,N26269,N26282);
or or1989(N24305,N26295,N26308);
or or1990(N24306,N26321,N26334);
or or1991(N24307,N26347,N26360);
or or1992(N24308,N26373,N26386);
or or1993(N24309,N26399,N26412);
or or1994(N24310,N26425,N26438);
or or1995(N24311,N26451,N26464);
or or1996(N24312,N26477,N26490);
or or1997(N24313,N26503,N26515);
or or1998(N24314,N26527,N26539);
or or1999(N24315,N26551,N26563);
or or2000(N24316,N26575,N26587);
or or2001(N24317,N26599,N26611);
or or2002(N24318,N26623,N26635);
or or2003(N24319,N26647,N26659);
or or2004(N24320,N26671,N26683);
or or2005(N24321,N26695,N26707);
or or2006(N24322,N26719,N26731);
or or2007(N24323,N26743,N26755);
or or2008(N24324,N26767,N26779);
or or2009(N24325,N26791,N26803);
or or2010(N24326,N26815,N26827);
or or2011(N24327,N26839,N26851);
or or2012(N24328,N26863,N26875);
or or2013(N24329,N26887,N26899);
or or2014(N24330,N26911,N26923);
or or2015(N24331,N26935,N26947);
or or2016(N24332,N26959,N26971);
or or2017(N24333,N26982,N26993);
or or2018(N24334,N27004,N27015);
or or2019(N24335,N27026,N27037);
or or2020(N24336,N27048,N27059);
or or2021(N24337,N27070,N27081);
or or2022(N24338,N27092,N27103);
or or2023(N24339,N27114,N27125);
or or2024(N24340,N27136,N27147);
or or2025(N24341,N27157,N27167);
or or2026(N24342,N27177,N27187);
or or2027(N24343,N27197,N27213);
or or2028(N24344,N27229,N27245);
or or2029(N24345,N27260,N27275);
or or2030(N24346,N27290,N27305);
or or2031(N24347,N27320,N27335);
or or2032(N24348,N27350,N27365);
or or2033(N24349,N27380,N27395);
or or2034(N24350,N27410,N27424);
or or2035(N24351,N27438,N27452);
or or2036(N24352,N27466,N27480);
or or2037(N24353,N27494,N27508);
or or2038(N24354,N27522,N27536);
or or2039(N24355,N27550,N27564);
or or2040(N24356,N27578,N27592);
or or2041(N24357,N27606,N27620);
or or2042(N24358,N27634,N27648);
or or2043(N24359,N27662,N27676);
or or2044(N24360,N27690,N27704);
or or2045(N24361,N27718,N27732);
or or2046(N24362,N27746,N27759);
or or2047(N24363,N27772,N27785);
or or2048(N24364,N27798,N27811);
or or2049(N24365,N27824,N27837);
or or2050(N24366,N27850,N27863);
or or2051(N24367,N27876,N27889);
or or2052(N24368,N27902,N27915);
or or2053(N24369,N27928,N27941);
or or2054(N24370,N27954,N27967);
or or2055(N24371,N27980,N27993);
or or2056(N24372,N28006,N28019);
or or2057(N24373,N28032,N28045);
or or2058(N24374,N28058,N28071);
or or2059(N24375,N28084,N28097);
or or2060(N24376,N28110,N28123);
or or2061(N24377,N28136,N28149);
or or2062(N24378,N28162,N28174);
or or2063(N24379,N28186,N28198);
or or2064(N24380,N28210,N28222);
or or2065(N24381,N28234,N28246);
or or2066(N24382,N28258,N28270);
or or2067(N24383,N28282,N28294);
or or2068(N24384,N28306,N28318);
or or2069(N24385,N28330,N28342);
or or2070(N24386,N28354,N28366);
or or2071(N24387,N28378,N28390);
or or2072(N24388,N28402,N28414);
or or2073(N24389,N28426,N28438);
or or2074(N24390,N28450,N28462);
or or2075(N24391,N28474,N28486);
or or2076(N24392,N28498,N28510);
or or2077(N24393,N28522,N28534);
or or2078(N24394,N28546,N28558);
or or2079(N24395,N28570,N28582);
or or2080(N24396,N28594,N28606);
or or2081(N24397,N28618,N28630);
or or2082(N24398,N28642,N28654);
or or2083(N24399,N28665,N28676);
or or2084(N24400,N28687,N28698);
or or2085(N24401,N28709,N28720);
or or2086(N24402,N28731,N28742);
or or2087(N24403,N28753,N28764);
or or2088(N24404,N28775,N28786);
or or2089(N24405,N28797,N28808);
or or2090(N24406,N28819,N28830);
or or2091(N24407,N28841,N28852);
or or2092(N24408,N28863,N28874);
or or2093(N24409,N28885,N28896);
or or2094(N24410,N28907,N28918);
or or2095(N24411,N28929,N28939);
or or2096(N24412,N28949,N28959);
or or2097(N24413,N28969,N28979);
or or2098(N24414,N28989,N28999);
or or2099(N24415,N29009,N29019);
or or2100(N24416,N29029,N29039);
or or2101(N24417,N29049,N29058);
or or2102(N24418,N29071,N29084);
or or2103(N24419,N29097,N29109);
or or2104(N24420,N29121,N29133);
or or2105(N24421,N29145,N29157);
or or2106(N24422,N29168,N29179);
or or2107(N24423,N29190,N29201);
or or2108(N24424,N29212,N29223);
or or2109(N24425,N29234,N29244);
or or2110(N24426,N29254,N29263);
or or2111(N29273,N29274,N29275);
or or2112(N29274,N29276,N29277);
or or2113(N29275,N29278,N29279);
or or2114(N29276,N29280,N29281);
or or2115(N29277,N29282,N29283);
or or2116(N29278,N29284,N29285);
or or2117(N29279,N29286,N29287);
or or2118(N29280,N29288,N29289);
or or2119(N29281,N29290,N29291);
or or2120(N29282,N29292,N29293);
or or2121(N29283,N29294,N29295);
or or2122(N29284,N29296,N29297);
or or2123(N29285,N29298,N29299);
or or2124(N29286,N29300,N29301);
or or2125(N29287,N29302,N29303);
or or2126(N29288,N29304,N29305);
or or2127(N29289,N29306,N29307);
or or2128(N29290,N29308,N29309);
or or2129(N29291,N29310,N29311);
or or2130(N29292,N29312,N29313);
or or2131(N29293,N29314,N29315);
or or2132(N29294,N29316,N29317);
or or2133(N29295,N29318,N29319);
or or2134(N29296,N29320,N29321);
or or2135(N29297,N29322,N29323);
or or2136(N29298,N29324,N29325);
or or2137(N29299,N29326,N29327);
or or2138(N29300,N29328,N29329);
or or2139(N29301,N29330,N29331);
or or2140(N29302,N29332,N29333);
or or2141(N29303,N29334,N29335);
or or2142(N29304,N29336,N29337);
or or2143(N29305,N29338,N29339);
or or2144(N29306,N29340,N29341);
or or2145(N29307,N29342,N29343);
or or2146(N29308,N29344,N29345);
or or2147(N29309,N29346,N29347);
or or2148(N29310,N29348,N29349);
or or2149(N29311,N29350,N29351);
or or2150(N29312,N29352,N29353);
or or2151(N29313,N29354,N29355);
or or2152(N29314,N29356,N29357);
or or2153(N29315,N29358,N29359);
or or2154(N29316,N29360,N29361);
or or2155(N29317,N29362,N29363);
or or2156(N29318,N29364,N29365);
or or2157(N29319,N29366,N29367);
or or2158(N29320,N29368,N29369);
or or2159(N29321,N29370,N29371);
or or2160(N29322,N29372,N29373);
or or2161(N29323,N29374,N29375);
or or2162(N29324,N29376,N29377);
or or2163(N29325,N29378,N29379);
or or2164(N29326,N29380,N29381);
or or2165(N29327,N29382,N29383);
or or2166(N29328,N29384,N29385);
or or2167(N29329,N29386,N29387);
or or2168(N29330,N29388,N29389);
or or2169(N29331,N29390,N29391);
or or2170(N29332,N29392,N29393);
or or2171(N29333,N29394,N29395);
or or2172(N29334,N29396,N29397);
or or2173(N29335,N29398,N29399);
or or2174(N29336,N29400,N29401);
or or2175(N29337,N29402,N29403);
or or2176(N29338,N29404,N29405);
or or2177(N29339,N29406,N29407);
or or2178(N29340,N29408,N29409);
or or2179(N29341,N29410,N29411);
or or2180(N29342,N29412,N29413);
or or2181(N29343,N29414,N29415);
or or2182(N29344,N29416,N29417);
or or2183(N29345,N29418,N29419);
or or2184(N29346,N29420,N29421);
or or2185(N29347,N29422,N29423);
or or2186(N29348,N29424,N29425);
or or2187(N29349,N29426,N29427);
or or2188(N29350,N29428,N29429);
or or2189(N29351,N29430,N29431);
or or2190(N29352,N29432,N29433);
or or2191(N29353,N29434,N29452);
or or2192(N29354,N29470,N29487);
or or2193(N29355,N29504,N29520);
or or2194(N29356,N29536,N29550);
or or2195(N29357,N29568,N29586);
or or2196(N29358,N29604,N29621);
or or2197(N29359,N29638,N29655);
or or2198(N29360,N29672,N29689);
or or2199(N29361,N29706,N29722);
or or2200(N29362,N29738,N29754);
or or2201(N29363,N29770,N29786);
or or2202(N29364,N29802,N29818);
or or2203(N29365,N29834,N29850);
or or2204(N29366,N29866,N29882);
or or2205(N29367,N29898,N29914);
or or2206(N29368,N29930,N29946);
or or2207(N29369,N29962,N29978);
or or2208(N29370,N29994,N30009);
or or2209(N29371,N30024,N30039);
or or2210(N29372,N30054,N30069);
or or2211(N29373,N30084,N30099);
or or2212(N29374,N30114,N30129);
or or2213(N29375,N30144,N30159);
or or2214(N29376,N30174,N30189);
or or2215(N29377,N30204,N30219);
or or2216(N29378,N30234,N30249);
or or2217(N29379,N30264,N30279);
or or2218(N29380,N30294,N30309);
or or2219(N29381,N30324,N30339);
or or2220(N29382,N30354,N30369);
or or2221(N29383,N30384,N30399);
or or2222(N29384,N30414,N30429);
or or2223(N29385,N30444,N30459);
or or2224(N29386,N30474,N30488);
or or2225(N29387,N30502,N30516);
or or2226(N29388,N30530,N30544);
or or2227(N29389,N30558,N30572);
or or2228(N29390,N30586,N30600);
or or2229(N29391,N30614,N30628);
or or2230(N29392,N30642,N30656);
or or2231(N29393,N30670,N30684);
or or2232(N29394,N30698,N30712);
or or2233(N29395,N30726,N30740);
or or2234(N29396,N30754,N30768);
or or2235(N29397,N30782,N30796);
or or2236(N29398,N30810,N30824);
or or2237(N29399,N30838,N30852);
or or2238(N29400,N30866,N30880);
or or2239(N29401,N30894,N30908);
or or2240(N29402,N30922,N30936);
or or2241(N29403,N30950,N30964);
or or2242(N29404,N30977,N30990);
or or2243(N29405,N31003,N31016);
or or2244(N29406,N31029,N31042);
or or2245(N29407,N31055,N31068);
or or2246(N29408,N31081,N31094);
or or2247(N29409,N31107,N31120);
or or2248(N29410,N31133,N31146);
or or2249(N29411,N31159,N31172);
or or2250(N29412,N31185,N31198);
or or2251(N29413,N31211,N31224);
or or2252(N29414,N31237,N31249);
or or2253(N29415,N31261,N31273);
or or2254(N29416,N31285,N31297);
or or2255(N29417,N31309,N31321);
or or2256(N29418,N31333,N31345);
or or2257(N29419,N31357,N31367);
or or2258(N29420,N31377,N31387);
or or2259(N29421,N31397,N31407);
or or2260(N29422,N31423,N31439);
or or2261(N29423,N31455,N31470);
or or2262(N29424,N31485,N31500);
or or2263(N29425,N31514,N31528);
or or2264(N29426,N31542,N31556);
or or2265(N29427,N31570,N31584);
or or2266(N29428,N31597,N31610);
or or2267(N29429,N31623,N31635);
or or2268(N29430,N31647,N31659);
or or2269(N29431,N31671,N31683);
or or2270(N29432,N31694,N31705);
or or2271(N29433,N31716,N31726);
or or2272(N31740,N31741,N31742);
or or2273(N31741,N31743,N31744);
or or2274(N31742,N31745,N31746);
or or2275(N31743,N31747,N31748);
or or2276(N31744,N31749,N31750);
or or2277(N31745,N31751,N31752);
or or2278(N31746,N31753,N31754);
or or2279(N31747,N31755,N31756);
or or2280(N31748,N31757,N31758);
or or2281(N31749,N31759,N31760);
or or2282(N31750,N31761,N31762);
or or2283(N31751,N31763,N31764);
or or2284(N31752,N31765,N31766);
or or2285(N31753,N31767,N31768);
or or2286(N31754,N31769,N31770);
or or2287(N31755,N31771,N31772);
or or2288(N31756,N31773,N31774);
or or2289(N31757,N31775,N31776);
or or2290(N31758,N31777,N31778);
or or2291(N31759,N31779,N31780);
or or2292(N31760,N31781,N31782);
or or2293(N31761,N31783,N31784);
or or2294(N31762,N31785,N31786);
or or2295(N31763,N31787,N31788);
or or2296(N31764,N31789,N31790);
or or2297(N31765,N31791,N31792);
or or2298(N31766,N31793,N31794);
or or2299(N31767,N31795,N31796);
or or2300(N31768,N31797,N31798);
or or2301(N31769,N31799,N31800);
or or2302(N31770,N31801,N31802);
or or2303(N31771,N31803,N31804);
or or2304(N31772,N31805,N31806);
or or2305(N31773,N31807,N31808);
or or2306(N31774,N31809,N31810);
or or2307(N31775,N31811,N31812);
or or2308(N31776,N31813,N31814);
or or2309(N31777,N31815,N31816);
or or2310(N31778,N31817,N31818);
or or2311(N31779,N31819,N31820);
or or2312(N31780,N31821,N31822);
or or2313(N31781,N31823,N31824);
or or2314(N31782,N31825,N31826);
or or2315(N31783,N31827,N31828);
or or2316(N31784,N31829,N31830);
or or2317(N31785,N31831,N31832);
or or2318(N31786,N31833,N31834);
or or2319(N31787,N31835,N31836);
or or2320(N31788,N31837,N31838);
or or2321(N31789,N31839,N31840);
or or2322(N31790,N31841,N31842);
or or2323(N31791,N31843,N31844);
or or2324(N31792,N31845,N31846);
or or2325(N31793,N31847,N31848);
or or2326(N31794,N31849,N31850);
or or2327(N31795,N31851,N31852);
or or2328(N31796,N31853,N31854);
or or2329(N31797,N31855,N31856);
or or2330(N31798,N31857,N31858);
or or2331(N31799,N31859,N31860);
or or2332(N31800,N31861,N31862);
or or2333(N31801,N31863,N31864);
or or2334(N31802,N31865,N31866);
or or2335(N31803,N31867,N31868);
or or2336(N31804,N31869,N31870);
or or2337(N31805,N31871,N31872);
or or2338(N31806,N31873,N31874);
or or2339(N31807,N31875,N31876);
or or2340(N31808,N31877,N31878);
or or2341(N31809,N31879,N31880);
or or2342(N31810,N31881,N31882);
or or2343(N31811,N31883,N31884);
or or2344(N31812,N31885,N31886);
or or2345(N31813,N31887,N31888);
or or2346(N31814,N31889,N31890);
or or2347(N31815,N31891,N31892);
or or2348(N31816,N31893,N31894);
or or2349(N31817,N31895,N31896);
or or2350(N31818,N31897,N31898);
or or2351(N31819,N31899,N31900);
or or2352(N31820,N31901,N31902);
or or2353(N31821,N31903,N31904);
or or2354(N31822,N31905,N31906);
or or2355(N31823,N31907,N31908);
or or2356(N31824,N31909,N31910);
or or2357(N31825,N31911,N31912);
or or2358(N31826,N31929,N31945);
or or2359(N31827,N31960,N31975);
or or2360(N31828,N31993,N32011);
or or2361(N31829,N32029,N32046);
or or2362(N31830,N32063,N32080);
or or2363(N31831,N32097,N32114);
or or2364(N31832,N32131,N32148);
or or2365(N31833,N32165,N32182);
or or2366(N31834,N32199,N32216);
or or2367(N31835,N32233,N32250);
or or2368(N31836,N32266,N32282);
or or2369(N31837,N32298,N32314);
or or2370(N31838,N32330,N32346);
or or2371(N31839,N32362,N32378);
or or2372(N31840,N32394,N32410);
or or2373(N31841,N32426,N32442);
or or2374(N31842,N32458,N32474);
or or2375(N31843,N32490,N32506);
or or2376(N31844,N32522,N32538);
or or2377(N31845,N32554,N32570);
or or2378(N31846,N32586,N32602);
or or2379(N31847,N32617,N32632);
or or2380(N31848,N32647,N32662);
or or2381(N31849,N32677,N32692);
or or2382(N31850,N32707,N32722);
or or2383(N31851,N32737,N32752);
or or2384(N31852,N32767,N32782);
or or2385(N31853,N32797,N32812);
or or2386(N31854,N32827,N32842);
or or2387(N31855,N32857,N32872);
or or2388(N31856,N32887,N32902);
or or2389(N31857,N32917,N32932);
or or2390(N31858,N32947,N32962);
or or2391(N31859,N32977,N32992);
or or2392(N31860,N33007,N33022);
or or2393(N31861,N33037,N33052);
or or2394(N31862,N33067,N33082);
or or2395(N31863,N33097,N33112);
or or2396(N31864,N33127,N33141);
or or2397(N31865,N33155,N33169);
or or2398(N31866,N33183,N33197);
or or2399(N31867,N33211,N33225);
or or2400(N31868,N33239,N33253);
or or2401(N31869,N33267,N33281);
or or2402(N31870,N33295,N33309);
or or2403(N31871,N33323,N33337);
or or2404(N31872,N33351,N33365);
or or2405(N31873,N33379,N33393);
or or2406(N31874,N33407,N33421);
or or2407(N31875,N33435,N33449);
or or2408(N31876,N33463,N33477);
or or2409(N31877,N33491,N33505);
or or2410(N31878,N33519,N33533);
or or2411(N31879,N33547,N33561);
or or2412(N31880,N33575,N33589);
or or2413(N31881,N33602,N33615);
or or2414(N31882,N33628,N33641);
or or2415(N31883,N33654,N33667);
or or2416(N31884,N33680,N33693);
or or2417(N31885,N33706,N33719);
or or2418(N31886,N33732,N33745);
or or2419(N31887,N33758,N33771);
or or2420(N31888,N33784,N33797);
or or2421(N31889,N33810,N33823);
or or2422(N31890,N33836,N33849);
or or2423(N31891,N33862,N33874);
or or2424(N31892,N33886,N33898);
or or2425(N31893,N33910,N33922);
or or2426(N31894,N33934,N33946);
or or2427(N31895,N33958,N33970);
or or2428(N31896,N33982,N33994);
or or2429(N31897,N34006,N34018);
or or2430(N31898,N34030,N34042);
or or2431(N31899,N34053,N34064);
or or2432(N31900,N34080,N34095);
or or2433(N31901,N34110,N34125);
or or2434(N31902,N34140,N34154);
or or2435(N31903,N34168,N34182);
or or2436(N31904,N34196,N34210);
or or2437(N31905,N34224,N34238);
or or2438(N31906,N34251,N34264);
or or2439(N31907,N34277,N34290);
or or2440(N31908,N34302,N34314);
or or2441(N31909,N34326,N34337);
or or2442(N31910,N34348,N34359);
or or2443(N31911,N34370,N34381);
or or2444(N34392,N34393,N34394);
or or2445(N34393,N34395,N34396);
or or2446(N34394,N34397,N34398);
or or2447(N34395,N34399,N34400);
or or2448(N34396,N34401,N34402);
or or2449(N34397,N34403,N34404);
or or2450(N34398,N34405,N34406);
or or2451(N34399,N34407,N34408);
or or2452(N34400,N34409,N34410);
or or2453(N34401,N34411,N34412);
or or2454(N34402,N34413,N34414);
or or2455(N34403,N34415,N34416);
or or2456(N34404,N34417,N34418);
or or2457(N34405,N34419,N34420);
or or2458(N34406,N34421,N34422);
or or2459(N34407,N34423,N34424);
or or2460(N34408,N34425,N34426);
or or2461(N34409,N34427,N34428);
or or2462(N34410,N34429,N34430);
or or2463(N34411,N34431,N34432);
or or2464(N34412,N34433,N34434);
or or2465(N34413,N34435,N34436);
or or2466(N34414,N34437,N34438);
or or2467(N34415,N34439,N34440);
or or2468(N34416,N34441,N34442);
or or2469(N34417,N34443,N34444);
or or2470(N34418,N34445,N34446);
or or2471(N34419,N34447,N34448);
or or2472(N34420,N34449,N34450);
or or2473(N34421,N34451,N34452);
or or2474(N34422,N34453,N34454);
or or2475(N34423,N34455,N34456);
or or2476(N34424,N34457,N34458);
or or2477(N34425,N34459,N34460);
or or2478(N34426,N34461,N34462);
or or2479(N34427,N34463,N34464);
or or2480(N34428,N34465,N34466);
or or2481(N34429,N34467,N34468);
or or2482(N34430,N34469,N34470);
or or2483(N34431,N34471,N34472);
or or2484(N34432,N34473,N34474);
or or2485(N34433,N34475,N34476);
or or2486(N34434,N34477,N34478);
or or2487(N34435,N34479,N34480);
or or2488(N34436,N34481,N34482);
or or2489(N34437,N34483,N34484);
or or2490(N34438,N34485,N34486);
or or2491(N34439,N34487,N34488);
or or2492(N34440,N34489,N34490);
or or2493(N34441,N34491,N34492);
or or2494(N34442,N34493,N34494);
or or2495(N34443,N34495,N34496);
or or2496(N34444,N34497,N34498);
or or2497(N34445,N34499,N34500);
or or2498(N34446,N34501,N34502);
or or2499(N34447,N34503,N34504);
or or2500(N34448,N34505,N34506);
or or2501(N34449,N34507,N34508);
or or2502(N34450,N34509,N34510);
or or2503(N34451,N34511,N34512);
or or2504(N34452,N34513,N34514);
or or2505(N34453,N34515,N34516);
or or2506(N34454,N34517,N34518);
or or2507(N34455,N34519,N34520);
or or2508(N34456,N34521,N34522);
or or2509(N34457,N34523,N34524);
or or2510(N34458,N34525,N34526);
or or2511(N34459,N34527,N34528);
or or2512(N34460,N34529,N34530);
or or2513(N34461,N34531,N34532);
or or2514(N34462,N34533,N34534);
or or2515(N34463,N34535,N34536);
or or2516(N34464,N34537,N34538);
or or2517(N34465,N34539,N34540);
or or2518(N34466,N34541,N34542);
or or2519(N34467,N34543,N34544);
or or2520(N34468,N34545,N34546);
or or2521(N34469,N34547,N34548);
or or2522(N34470,N34549,N34550);
or or2523(N34471,N34551,N34552);
or or2524(N34472,N34553,N34554);
or or2525(N34473,N34555,N34556);
or or2526(N34474,N34557,N34558);
or or2527(N34475,N34559,N34560);
or or2528(N34476,N34561,N34562);
or or2529(N34477,N34563,N34564);
or or2530(N34478,N34565,N34566);
or or2531(N34479,N34567,N34568);
or or2532(N34480,N34569,N34570);
or or2533(N34481,N34571,N34572);
or or2534(N34482,N34573,N34574);
or or2535(N34483,N34575,N34576);
or or2536(N34484,N34577,N34578);
or or2537(N34485,N34579,N34580);
or or2538(N34486,N34581,N34582);
or or2539(N34487,N34602,N34620);
or or2540(N34488,N34637,N34655);
or or2541(N34489,N34673,N34691);
or or2542(N34490,N34709,N34727);
or or2543(N34491,N34744,N34761);
or or2544(N34492,N34778,N34794);
or or2545(N34493,N34810,N34826);
or or2546(N34494,N34842,N34858);
or or2547(N34495,N34874,N34890);
or or2548(N34496,N34906,N34922);
or or2549(N34497,N34938,N34954);
or or2550(N34498,N34970,N34986);
or or2551(N34499,N35002,N35018);
or or2552(N34500,N35034,N35050);
or or2553(N34501,N35066,N35082);
or or2554(N34502,N35098,N35114);
or or2555(N34503,N35130,N35146);
or or2556(N34504,N35161,N35176);
or or2557(N34505,N35191,N35206);
or or2558(N34506,N35221,N35236);
or or2559(N34507,N35251,N35266);
or or2560(N34508,N35281,N35296);
or or2561(N34509,N35311,N35326);
or or2562(N34510,N35341,N35356);
or or2563(N34511,N35371,N35386);
or or2564(N34512,N35401,N35416);
or or2565(N34513,N35431,N35446);
or or2566(N34514,N35461,N35476);
or or2567(N34515,N35491,N35506);
or or2568(N34516,N35521,N35536);
or or2569(N34517,N35551,N35566);
or or2570(N34518,N35581,N35596);
or or2571(N34519,N35610,N35624);
or or2572(N34520,N35638,N35652);
or or2573(N34521,N35666,N35680);
or or2574(N34522,N35694,N35708);
or or2575(N34523,N35722,N35736);
or or2576(N34524,N35750,N35764);
or or2577(N34525,N35778,N35792);
or or2578(N34526,N35806,N35820);
or or2579(N34527,N35834,N35848);
or or2580(N34528,N35862,N35876);
or or2581(N34529,N35890,N35904);
or or2582(N34530,N35918,N35932);
or or2583(N34531,N35946,N35960);
or or2584(N34532,N35974,N35988);
or or2585(N34533,N36002,N36016);
or or2586(N34534,N36030,N36044);
or or2587(N34535,N36058,N36072);
or or2588(N34536,N36086,N36100);
or or2589(N34537,N36114,N36128);
or or2590(N34538,N36142,N36156);
or or2591(N34539,N36170,N36184);
or or2592(N34540,N36197,N36210);
or or2593(N34541,N36223,N36236);
or or2594(N34542,N36249,N36262);
or or2595(N34543,N36275,N36288);
or or2596(N34544,N36301,N36314);
or or2597(N34545,N36327,N36340);
or or2598(N34546,N36353,N36366);
or or2599(N34547,N36379,N36392);
or or2600(N34548,N36405,N36418);
or or2601(N34549,N36431,N36444);
or or2602(N34550,N36457,N36470);
or or2603(N34551,N36483,N36496);
or or2604(N34552,N36509,N36522);
or or2605(N34553,N36535,N36548);
or or2606(N34554,N36561,N36574);
or or2607(N34555,N36587,N36600);
or or2608(N34556,N36613,N36626);
or or2609(N34557,N36639,N36651);
or or2610(N34558,N36663,N36675);
or or2611(N34559,N36687,N36699);
or or2612(N34560,N36711,N36723);
or or2613(N34561,N36735,N36747);
or or2614(N34562,N36758,N36769);
or or2615(N34563,N36780,N36791);
or or2616(N34564,N36802,N36813);
or or2617(N34565,N36828,N36843);
or or2618(N34566,N36858,N36873);
or or2619(N34567,N36888,N36902);
or or2620(N34568,N36916,N36930);
or or2621(N34569,N36944,N36958);
or or2622(N34570,N36972,N36986);
or or2623(N34571,N37000,N37014);
or or2624(N34572,N37028,N37042);
or or2625(N34573,N37055,N37068);
or or2626(N34574,N37081,N37094);
or or2627(N34575,N37107,N37119);
or or2628(N34576,N37131,N37143);
or or2629(N34577,N37155,N37167);
or or2630(N34578,N37179,N37190);
or or2631(N34579,N37201,N37212);
or or2632(N34580,N37222,N37232);
or or2633(N34581,N37242,N37253);
or or2634(N37264,N37265,N37266);
or or2635(N37265,N37267,N37268);
or or2636(N37266,N37269,N37270);
or or2637(N37267,N37271,N37272);
or or2638(N37268,N37273,N37274);
or or2639(N37269,N37275,N37276);
or or2640(N37270,N37277,N37278);
or or2641(N37271,N37279,N37280);
or or2642(N37272,N37281,N37282);
or or2643(N37273,N37283,N37284);
or or2644(N37274,N37285,N37286);
or or2645(N37275,N37287,N37288);
or or2646(N37276,N37289,N37290);
or or2647(N37277,N37291,N37292);
or or2648(N37278,N37293,N37294);
or or2649(N37279,N37295,N37296);
or or2650(N37280,N37297,N37298);
or or2651(N37281,N37299,N37300);
or or2652(N37282,N37301,N37302);
or or2653(N37283,N37303,N37304);
or or2654(N37284,N37305,N37306);
or or2655(N37285,N37307,N37308);
or or2656(N37286,N37309,N37310);
or or2657(N37287,N37311,N37312);
or or2658(N37288,N37313,N37314);
or or2659(N37289,N37315,N37316);
or or2660(N37290,N37317,N37318);
or or2661(N37291,N37319,N37320);
or or2662(N37292,N37321,N37322);
or or2663(N37293,N37332,N37344);
or or2664(N37294,N37356,N37368);
or or2665(N37295,N37380,N37392);
or or2666(N37296,N37404,N37415);
or or2667(N37297,N37426,N37437);
or or2668(N37298,N37448,N37459);
or or2669(N37299,N37470,N37481);
or or2670(N37300,N37492,N37503);
or or2671(N37301,N37514,N37525);
or or2672(N37302,N37536,N37546);
or or2673(N37303,N37556,N37566);
or or2674(N37304,N37576,N37586);
or or2675(N37305,N37596,N37606);
or or2676(N37306,N37616,N37626);
or or2677(N37307,N37636,N37645);
or or2678(N37308,N37654,N37663);
or or2679(N37309,N37672,N37681);
or or2680(N37310,N37690,N37699);
or or2681(N37311,N37708,N37717);
or or2682(N37312,N37726,N37735);
or or2683(N37313,N37744,N37753);
or or2684(N37314,N37762,N37770);
or or2685(N37315,N37778,N37786);
or or2686(N37316,N37794,N37802);
or or2687(N37317,N37810,N37818);
or or2688(N37318,N37825,N37832);
or or2689(N37319,N37839,N37846);
or or2690(N37320,N37853,N37860);
or or2691(N37321,N37867,N37876);
or or2692(N37882,N37883,N37884);
or or2693(N37883,N37885,N37886);
or or2694(N37884,N37887,N37888);
or or2695(N37885,N37889,N37890);
or or2696(N37886,N37891,N37892);
or or2697(N37887,N37893,N37894);
or or2698(N37888,N37895,N37896);
or or2699(N37889,N37897,N37898);
or or2700(N37890,N37899,N37900);
or or2701(N37891,N37901,N37902);
or or2702(N37892,N37903,N37904);
or or2703(N37893,N37905,N37906);
or or2704(N37894,N37907,N37908);
or or2705(N37895,N37909,N37910);
or or2706(N37896,N37911,N37912);
or or2707(N37897,N37913,N37928);
or or2708(N37898,N37939,N37950);
or or2709(N37899,N37961,N37972);
or or2710(N37900,N37983,N37993);
or or2711(N37901,N38003,N38013);
or or2712(N37902,N38023,N38033);
or or2713(N37903,N38043,N38052);
or or2714(N37904,N38061,N38070);
or or2715(N37905,N38079,N38088);
or or2716(N37906,N38097,N38106);
or or2717(N37907,N38115,N38124);
or or2718(N37908,N38133,N38141);
or or2719(N37909,N38149,N38157);
or or2720(N37910,N38165,N38173);
or or2721(N37911,N38181,N38189);
or or2722(N37912,N38197,N38205);
or or2723(N38213,N38214,N38215);
or or2724(N38214,N38216,N38217);
or or2725(N38215,N38218,N38219);
or or2726(N38216,N38220,N38221);
or or2727(N38217,N38222,N38223);
or or2728(N38218,N38224,N38225);
or or2729(N38219,N38237,N38249);
or or2730(N38220,N38260,N38271);
or or2731(N38221,N38282,N38293);
or or2732(N38222,N38304,N38314);
or or2733(N38223,N38323,N38332);
or or2734(N38224,N38343,N38354);
or or2735(N38364,N38365,N38366);
or or2736(N38365,N38367,N38368);
or or2737(N38366,N38369,N38370);
or or2738(N38367,N38371,N38372);
or or2739(N38368,N38373,N38374);
or or2740(N38369,N38375,N38376);
or or2741(N38370,N38377,N38378);
or or2742(N38371,N38379,N38380);
or or2743(N38372,N38381,N38382);
or or2744(N38373,N38383,N38384);
or or2745(N38374,N38385,N38386);
or or2746(N38375,N38387,N38388);
or or2747(N38376,N38389,N38390);
or or2748(N38377,N38391,N38392);
or or2749(N38378,N38393,N38394);
or or2750(N38379,N38395,N38396);
or or2751(N38380,N38397,N38398);
or or2752(N38381,N38399,N38400);
or or2753(N38382,N38401,N38402);
or or2754(N38383,N38403,N38418);
or or2755(N38384,N38429,N38440);
or or2756(N38385,N38451,N38462);
or or2757(N38386,N38472,N38482);
or or2758(N38387,N38492,N38502);
or or2759(N38388,N38512,N38522);
or or2760(N38389,N38532,N38541);
or or2761(N38390,N38550,N38559);
or or2762(N38391,N38568,N38577);
or or2763(N38392,N38586,N38595);
or or2764(N38393,N38604,N38613);
or or2765(N38394,N38622,N38631);
or or2766(N38395,N38640,N38649);
or or2767(N38396,N38657,N38665);
or or2768(N38397,N38673,N38681);
or or2769(N38398,N38689,N38697);
or or2770(N38399,N38705,N38713);
or or2771(N38400,N38721,N38729);
or or2772(N38401,N38737,N38746);
or or2773(N38402,N38755,N38764);
or or2774(N38772,N38773,N38774);
or or2775(N38773,N38775,N38776);
or or2776(N38774,N38777,N38778);
or or2777(N38775,N38779,N38780);
or or2778(N38776,N38781,N38782);
or or2779(N38777,N38783,N38784);
or or2780(N38778,N38785,N38786);
or or2781(N38779,N38787,N38788);
or or2782(N38780,N38789,N38790);
or or2783(N38781,N38791,N38792);
or or2784(N38782,N38793,N38794);
or or2785(N38783,N38807,N38820);
or or2786(N38784,N38833,N38845);
or or2787(N38785,N38856,N38867);
or or2788(N38786,N38878,N38889);
or or2789(N38787,N38900,N38911);
or or2790(N38788,N38922,N38932);
or or2791(N38789,N38942,N38951);
or or2792(N38790,N38960,N38968);
or or2793(N38791,N38976,N38988);
or or2794(N38792,N39000,N39011);
or or2795(N38793,N39021,N39028);
or or2796(N39035,N39036,N39037);
or or2797(N39036,N39038,N39039);
or or2798(N39037,N39040,N39041);
or or2799(N39038,N39042,N39043);
or or2800(N39039,N39044,N39045);
or or2801(N39040,N39046,N39047);
or or2802(N39041,N39048,N39049);
or or2803(N39042,N39050,N39051);
or or2804(N39043,N39052,N39053);
or or2805(N39044,N39054,N39055);
or or2806(N39045,N39056,N39057);
or or2807(N39046,N39058,N39059);
or or2808(N39047,N39060,N39061);
or or2809(N39048,N39062,N39063);
or or2810(N39049,N39064,N39065);
or or2811(N39050,N39066,N39067);
or or2812(N39051,N39068,N39069);
or or2813(N39052,N39070,N39071);
or or2814(N39053,N39072,N39073);
or or2815(N39054,N39074,N39075);
or or2816(N39055,N39076,N39077);
or or2817(N39056,N39078,N39079);
or or2818(N39057,N39080,N39090);
or or2819(N39058,N39099,N39111);
or or2820(N39059,N39123,N39135);
or or2821(N39060,N39147,N39159);
or or2822(N39061,N39170,N39181);
or or2823(N39062,N39192,N39203);
or or2824(N39063,N39214,N39225);
or or2825(N39064,N39236,N39247);
or or2826(N39065,N39257,N39267);
or or2827(N39066,N39277,N39287);
or or2828(N39067,N39297,N39307);
or or2829(N39068,N39317,N39327);
or or2830(N39069,N39337,N39347);
or or2831(N39070,N39357,N39367);
or or2832(N39071,N39377,N39386);
or or2833(N39072,N39395,N39404);
or or2834(N39073,N39413,N39422);
or or2835(N39074,N39431,N39440);
or or2836(N39075,N39448,N39456);
or or2837(N39076,N39464,N39472);
or or2838(N39077,N39480,N39488);
or or2839(N39078,N39496,N39504);
or or2840(N39079,N39512,N39519);

not not0(N397,in0);
not not1(N398,in2);
not not2(N399,R0);
not not3(N400,R1);
not not4(N414,in2);
not not5(N415,R0);
not not6(N416,R1);
not not7(N417,R2);
not not8(N418,R3);
not not9(N431,in0);
not not10(N432,in1);
not not11(N433,R0);
not not12(N434,R1);
not not13(N435,R2);
not not14(N436,R3);
not not15(N448,in0);
not not16(N449,in1);
not not17(N450,in2);
not not18(N451,R0);
not not19(N452,R2);
not not20(N465,in0);
not not21(N466,in1);
not not22(N467,R1);
not not23(N468,R2);
not not24(N469,R3);
not not25(N482,in2);
not not26(N483,R0);
not not27(N484,R1);
not not28(N485,R2);
not not29(N486,R3);
not not30(N498,in0);
not not31(N499,in2);
not not32(N500,R0);
not not33(N501,R1);
not not34(N502,R2);
not not35(N514,in0);
not not36(N515,R1);
not not37(N516,R2);
not not38(N517,R3);
not not39(N530,in2);
not not40(N531,R0);
not not41(N532,R1);
not not42(N533,R2);
not not43(N546,in0);
not not44(N547,R0);
not not45(N548,R1);
not not46(N549,R2);
not not47(N562,in1);
not not48(N563,R0);
not not49(N564,R3);
not not50(N578,in2);
not not51(N579,R0);
not not52(N580,R1);
not not53(N581,R3);
not not54(N594,in0);
not not55(N595,in2);
not not56(N596,R2);
not not57(N597,R3);
not not58(N610,in1);
not not59(N611,in2);
not not60(N612,R0);
not not61(N613,R1);
not not62(N626,in0);
not not63(N627,in1);
not not64(N628,R1);
not not65(N642,in1);
not not66(N643,in2);
not not67(N644,R0);
not not68(N645,R1);
not not69(N646,R2);
not not70(N658,in0);
not not71(N659,in2);
not not72(N660,R0);
not not73(N661,R1);
not not74(N662,R2);
not not75(N674,in0);
not not76(N675,in1);
not not77(N676,in2);
not not78(N677,R1);
not not79(N678,R2);
not not80(N690,in0);
not not81(N691,in2);
not not82(N692,R3);
not not83(N706,in0);
not not84(N707,in2);
not not85(N708,R1);
not not86(N709,R2);
not not87(N710,R3);
not not88(N722,in1);
not not89(N723,in2);
not not90(N724,R0);
not not91(N725,R2);
not not92(N738,in0);
not not93(N739,in1);
not not94(N740,in2);
not not95(N741,R0);
not not96(N742,R2);
not not97(N754,in0);
not not98(N755,R0);
not not99(N756,R1);
not not100(N770,in0);
not not101(N771,in1);
not not102(N772,in2);
not not103(N773,R2);
not not104(N774,R3);
not not105(N786,in2);
not not106(N787,R0);
not not107(N788,R1);
not not108(N802,in0);
not not109(N803,in1);
not not110(N804,in2);
not not111(N805,R1);
not not112(N818,in1);
not not113(N819,in2);
not not114(N820,R0);
not not115(N833,in1);
not not116(N834,R0);
not not117(N835,R2);
not not118(N848,in0);
not not119(N849,in2);
not not120(N850,R1);
not not121(N851,R2);
not not122(N863,in0);
not not123(N864,in1);
not not124(N865,in2);
not not125(N866,R0);
not not126(N878,in0);
not not127(N879,in1);
not not128(N880,in2);
not not129(N881,R0);
not not130(N893,in1);
not not131(N894,in2);
not not132(N895,R1);
not not133(N896,R3);
not not134(N908,in0);
not not135(N909,in2);
not not136(N910,R1);
not not137(N923,in1);
not not138(N924,in2);
not not139(N925,R1);
not not140(N926,R2);
not not141(N938,in0);
not not142(N939,in1);
not not143(N940,R0);
not not144(N941,R1);
not not145(N953,in0);
not not146(N954,in2);
not not147(N955,R0);
not not148(N956,R2);
not not149(N968,in0);
not not150(N969,in1);
not not151(N970,in2);
not not152(N971,R3);
not not153(N983,in2);
not not154(N984,R1);
not not155(N985,R2);
not not156(N998,in1);
not not157(N999,R0);
not not158(N1000,R1);
not not159(N1001,R3);
not not160(N1013,in0);
not not161(N1014,in1);
not not162(N1015,R1);
not not163(N1028,in1);
not not164(N1029,R1);
not not165(N1030,R2);
not not166(N1043,in2);
not not167(N1044,R1);
not not168(N1045,R2);
not not169(N1058,in0);
not not170(N1059,in1);
not not171(N1060,R1);
not not172(N1061,R2);
not not173(N1073,in0);
not not174(N1074,in2);
not not175(N1075,R0);
not not176(N1076,R1);
not not177(N1088,in2);
not not178(N1089,R0);
not not179(N1090,R2);
not not180(N1091,R3);
not not181(N1103,R0);
not not182(N1104,R2);
not not183(N1105,R3);
not not184(N1118,in0);
not not185(N1119,in1);
not not186(N1120,R0);
not not187(N1121,R3);
not not188(N1133,in0);
not not189(N1134,in1);
not not190(N1135,in2);
not not191(N1136,R3);
not not192(N1148,R0);
not not193(N1149,R1);
not not194(N1150,R3);
not not195(N1163,in0);
not not196(N1164,R1);
not not197(N1178,in0);
not not198(N1179,R0);
not not199(N1180,R2);
not not200(N1181,R3);
not not201(N1193,in0);
not not202(N1194,in2);
not not203(N1195,R0);
not not204(N1196,R2);
not not205(N1208,in1);
not not206(N1209,R1);
not not207(N1210,R2);
not not208(N1223,in2);
not not209(N1224,R1);
not not210(N1225,R2);
not not211(N1238,in0);
not not212(N1239,in2);
not not213(N1240,R1);
not not214(N1241,R2);
not not215(N1253,in0);
not not216(N1254,R1);
not not217(N1255,R3);
not not218(N1268,in0);
not not219(N1269,in1);
not not220(N1270,R0);
not not221(N1271,R2);
not not222(N1272,R3);
not not223(N1283,in0);
not not224(N1284,R1);
not not225(N1285,R2);
not not226(N1298,in0);
not not227(N1299,in2);
not not228(N1300,R0);
not not229(N1313,in0);
not not230(N1314,in1);
not not231(N1315,R1);
not not232(N1328,in2);
not not233(N1329,R1);
not not234(N1330,R3);
not not235(N1343,in0);
not not236(N1344,in1);
not not237(N1345,R0);
not not238(N1346,R3);
not not239(N1358,in0);
not not240(N1359,in2);
not not241(N1360,R0);
not not242(N1361,R1);
not not243(N1373,in0);
not not244(N1374,in1);
not not245(N1375,in2);
not not246(N1388,in0);
not not247(N1389,in1);
not not248(N1390,R0);
not not249(N1391,R1);
not not250(N1403,in0);
not not251(N1404,R0);
not not252(N1405,R3);
not not253(N1418,in0);
not not254(N1419,in1);
not not255(N1420,R0);
not not256(N1421,R1);
not not257(N1433,in1);
not not258(N1434,R0);
not not259(N1435,R2);
not not260(N1447,in0);
not not261(N1448,in1);
not not262(N1449,R0);
not not263(N1450,R2);
not not264(N1461,in0);
not not265(N1462,R0);
not not266(N1475,in1);
not not267(N1476,R0);
not not268(N1489,R0);
not not269(N1503,in0);
not not270(N1504,in2);
not not271(N1505,R0);
not not272(N1506,R2);
not not273(N1517,in2);
not not274(N1518,R0);
not not275(N1519,R2);
not not276(N1531,R1);
not not277(N1532,R3);
not not278(N1545,R1);
not not279(N1546,R2);
not not280(N1559,in2);
not not281(N1573,R3);
not not282(N1587,in2);
not not283(N1588,R2);
not not284(N1601,in0);
not not285(N1602,R0);
not not286(N1615,in1);
not not287(N1616,in2);
not not288(N1617,R1);
not not289(N1618,R2);
not not290(N1629,in1);
not not291(N1630,R0);
not not292(N1631,R1);
not not293(N1643,in2);
not not294(N1644,R0);
not not295(N1657,in1);
not not296(N1658,in2);
not not297(N1659,R0);
not not298(N1671,in0);
not not299(N1672,R3);
not not300(N1685,in0);
not not301(N1686,in2);
not not302(N1687,R1);
not not303(N1699,in2);
not not304(N1700,R0);
not not305(N1701,R3);
not not306(N1713,R0);
not not307(N1714,R1);
not not308(N1715,R2);
not not309(N1727,in2);
not not310(N1728,R0);
not not311(N1729,R2);
not not312(N1741,in2);
not not313(N1742,R1);
not not314(N1743,R3);
not not315(N1755,in0);
not not316(N1756,in2);
not not317(N1757,R1);
not not318(N1758,R2);
not not319(N1769,in2);
not not320(N1770,R0);
not not321(N1771,R1);
not not322(N1783,in0);
not not323(N1784,R0);
not not324(N1785,R2);
not not325(N1797,in0);
not not326(N1798,R0);
not not327(N1799,R1);
not not328(N1811,in0);
not not329(N1812,in1);
not not330(N1813,in2);
not not331(N1814,R2);
not not332(N1825,R0);
not not333(N1826,R1);
not not334(N1827,R2);
not not335(N1839,in0);
not not336(N1840,R0);
not not337(N1841,R1);
not not338(N1842,R2);
not not339(N1853,R1);
not not340(N1867,in0);
not not341(N1868,in2);
not not342(N1869,R0);
not not343(N1870,R1);
not not344(N1881,in2);
not not345(N1882,R0);
not not346(N1895,in0);
not not347(N1896,in2);
not not348(N1897,R2);
not not349(N1909,in0);
not not350(N1910,in2);
not not351(N1911,R2);
not not352(N1923,in0);
not not353(N1924,in1);
not not354(N1925,R1);
not not355(N1926,R3);
not not356(N1937,in0);
not not357(N1938,in2);
not not358(N1939,R1);
not not359(N1940,R3);
not not360(N1951,in0);
not not361(N1952,in2);
not not362(N1953,R2);
not not363(N1954,R3);
not not364(N1965,in0);
not not365(N1966,in1);
not not366(N1967,R0);
not not367(N1968,R3);
not not368(N1979,in0);
not not369(N1980,in1);
not not370(N1981,in2);
not not371(N1982,R0);
not not372(N1983,R2);
not not373(N1993,R0);
not not374(N1994,R3);
not not375(N2007,in0);
not not376(N2008,R0);
not not377(N2021,in2);
not not378(N2022,R1);
not not379(N2035,in0);
not not380(N2036,in1);
not not381(N2037,R2);
not not382(N2049,in0);
not not383(N2050,in1);
not not384(N2051,R1);
not not385(N2063,in2);
not not386(N2064,R3);
not not387(N2077,in0);
not not388(N2078,in1);
not not389(N2079,R0);
not not390(N2080,R1);
not not391(N2091,in0);
not not392(N2092,R3);
not not393(N2105,in0);
not not394(N2106,in1);
not not395(N2107,R2);
not not396(N2132,R2);
not not397(N2145,R1);
not not398(N2158,in1);
not not399(N2159,R0);
not not400(N2171,in0);
not not401(N2172,in2);
not not402(N2173,R0);
not not403(N2184,R1);
not not404(N2185,R3);
not not405(N2197,in0);
not not406(N2198,R1);
not not407(N2210,in0);
not not408(N2211,R2);
not not409(N2223,in1);
not not410(N2224,R1);
not not411(N2236,R1);
not not412(N2237,R3);
not not413(N2249,R0);
not not414(N2262,in0);
not not415(N2263,in1);
not not416(N2264,R1);
not not417(N2275,in0);
not not418(N2276,in1);
not not419(N2277,R3);
not not420(N2288,R1);
not not421(N2289,R2);
not not422(N2301,in1);
not not423(N2314,in0);
not not424(N2315,R0);
not not425(N2327,in0);
not not426(N2328,in2);
not not427(N2340,in0);
not not428(N2341,R2);
not not429(N2342,R3);
not not430(N2353,in1);
not not431(N2354,R0);
not not432(N2355,R1);
not not433(N2366,in1);
not not434(N2367,R2);
not not435(N2379,in2);
not not436(N2380,R0);
not not437(N2381,R1);
not not438(N2392,in1);
not not439(N2393,R1);
not not440(N2405,R1);
not not441(N2406,R2);
not not442(N2418,in1);
not not443(N2419,in2);
not not444(N2431,in0);
not not445(N2432,in2);
not not446(N2444,in0);
not not447(N2445,R0);
not not448(N2457,R0);
not not449(N2458,R2);
not not450(N2470,in1);
not not451(N2471,R0);
not not452(N2472,R2);
not not453(N2483,in2);
not not454(N2484,R0);
not not455(N2485,R2);
not not456(N2496,in0);
not not457(N2497,R1);
not not458(N2509,in0);
not not459(N2510,in2);
not not460(N2511,R0);
not not461(N2522,in1);
not not462(N2523,R2);
not not463(N2535,R3);
not not464(N2548,in0);
not not465(N2549,R1);
not not466(N2550,R2);
not not467(N2561,in0);
not not468(N2562,in1);
not not469(N2563,R1);
not not470(N2574,in0);
not not471(N2575,in1);
not not472(N2576,in2);
not not473(N2587,in0);
not not474(N2588,R1);
not not475(N2600,in0);
not not476(N2601,in2);
not not477(N2602,R0);
not not478(N2613,R3);
not not479(N2625,R0);
not not480(N2626,R2);
not not481(N2637,in0);
not not482(N2649,R3);
not not483(N2661,R3);
not not484(N2673,R1);
not not485(N2685,in0);
not not486(N2686,R0);
not not487(N2697,R2);
not not488(N2698,R3);
not not489(N2709,R0);
not not490(N2721,in0);
not not491(N2722,R3);
not not492(N2733,in2);
not not493(N2734,R3);
not not494(N2745,R1);
not not495(N2746,R2);
not not496(N2757,R1);
not not497(N2758,R2);
not not498(N2769,R0);
not not499(N2770,R1);
not not500(N2781,in0);
not not501(N2782,in2);
not not502(N2793,in2);
not not503(N2805,R2);
not not504(N2817,R1);
not not505(N2829,R0);
not not506(N2830,R1);
not not507(N2841,R0);
not not508(N2842,R2);
not not509(N2853,in0);
not not510(N2854,R0);
not not511(N2855,R2);
not not512(N2865,in2);
not not513(N2866,R0);
not not514(N2877,in0);
not not515(N2889,in0);
not not516(N2890,in1);
not not517(N2891,in2);
not not518(N2901,in0);
not not519(N2902,in1);
not not520(N2903,in2);
not not521(N2913,R0);
not not522(N2925,in0);
not not523(N2926,in1);
not not524(N2927,R2);
not not525(N2937,in0);
not not526(N2938,R1);
not not527(N2949,in0);
not not528(N2950,in2);
not not529(N2961,in0);
not not530(N2962,in2);
not not531(N2973,in0);
not not532(N2974,in1);
not not533(N2985,in0);
not not534(N2986,R3);
not not535(N2997,in0);
not not536(N2998,in1);
not not537(N2999,R0);
not not538(N3009,R0);
not not539(N3010,R1);
not not540(N3033,in0);
not not541(N3034,R0);
not not542(N3045,R3);
not not543(N3057,R2);
not not544(N3069,in0);
not not545(N3070,in2);
not not546(N3081,in0);
not not547(N3093,R2);
not not548(N3115,in0);
not not549(N3126,R1);
not not550(N3170,in0);
not not551(N3171,R1);
not not552(N3181,R1);
not not553(N3192,R0);
not not554(N3203,in1);
not not555(N3204,R0);
not not556(N3214,in0);
not not557(N3215,R0);
not not558(N3236,in2);
not not559(N3246,R0);
not not560(N3264,in0);
not not561(N3265,in1);
not not562(N3266,R0);
not not563(N3267,R2);
not not564(N3268,R4);
not not565(N3269,R5);
not not566(N3280,in1);
not not567(N3281,in2);
not not568(N3282,R0);
not not569(N3283,R1);
not not570(N3284,R2);
not not571(N3285,R4);
not not572(N3286,R5);
not not573(N3296,in0);
not not574(N3297,in1);
not not575(N3298,R0);
not not576(N3299,R1);
not not577(N3300,R2);
not not578(N3301,R3);
not not579(N3312,in0);
not not580(N3313,in1);
not not581(N3314,R0);
not not582(N3315,R1);
not not583(N3316,R3);
not not584(N3317,R4);
not not585(N3328,in0);
not not586(N3329,in1);
not not587(N3330,in2);
not not588(N3331,R0);
not not589(N3332,R2);
not not590(N3333,R5);
not not591(N3344,in1);
not not592(N3345,in2);
not not593(N3346,R1);
not not594(N3347,R2);
not not595(N3348,R4);
not not596(N3349,R5);
not not597(N3360,in0);
not not598(N3361,in1);
not not599(N3362,in2);
not not600(N3363,R0);
not not601(N3364,R1);
not not602(N3365,R4);
not not603(N3366,R5);
not not604(N3376,in1);
not not605(N3377,R0);
not not606(N3378,R1);
not not607(N3379,R2);
not not608(N3380,R3);
not not609(N3381,R5);
not not610(N3391,in0);
not not611(N3392,in2);
not not612(N3393,R0);
not not613(N3394,R1);
not not614(N3395,R5);
not not615(N3406,in0);
not not616(N3407,in1);
not not617(N3408,in2);
not not618(N3409,R4);
not not619(N3410,R5);
not not620(N3421,in0);
not not621(N3422,R0);
not not622(N3423,R1);
not not623(N3424,R2);
not not624(N3425,R4);
not not625(N3436,in0);
not not626(N3437,in1);
not not627(N3438,R0);
not not628(N3439,R2);
not not629(N3440,R4);
not not630(N3441,R5);
not not631(N3451,in0);
not not632(N3452,in2);
not not633(N3453,R2);
not not634(N3454,R3);
not not635(N3455,R5);
not not636(N3466,in0);
not not637(N3467,in2);
not not638(N3468,R0);
not not639(N3469,R2);
not not640(N3470,R4);
not not641(N3481,in1);
not not642(N3482,R0);
not not643(N3483,R1);
not not644(N3484,R2);
not not645(N3485,R4);
not not646(N3496,in0);
not not647(N3497,in2);
not not648(N3498,R0);
not not649(N3499,R2);
not not650(N3500,R4);
not not651(N3501,R5);
not not652(N3511,in0);
not not653(N3512,in1);
not not654(N3513,R0);
not not655(N3514,R2);
not not656(N3515,R3);
not not657(N3526,in0);
not not658(N3527,in2);
not not659(N3528,R0);
not not660(N3529,R3);
not not661(N3530,R4);
not not662(N3540,in1);
not not663(N3541,in2);
not not664(N3542,R2);
not not665(N3543,R4);
not not666(N3554,in0);
not not667(N3555,R0);
not not668(N3556,R3);
not not669(N3557,R5);
not not670(N3568,in2);
not not671(N3569,R0);
not not672(N3570,R4);
not not673(N3571,R5);
not not674(N3582,in1);
not not675(N3583,in2);
not not676(N3584,R0);
not not677(N3585,R4);
not not678(N3596,in1);
not not679(N3597,R1);
not not680(N3598,R3);
not not681(N3599,R4);
not not682(N3600,R5);
not not683(N3610,in1);
not not684(N3611,R1);
not not685(N3612,R4);
not not686(N3613,R5);
not not687(N3624,R0);
not not688(N3625,R1);
not not689(N3626,R2);
not not690(N3627,R4);
not not691(N3628,R5);
not not692(N3638,in0);
not not693(N3639,in2);
not not694(N3640,R4);
not not695(N3641,R5);
not not696(N3652,in0);
not not697(N3653,in2);
not not698(N3654,R2);
not not699(N3655,R4);
not not700(N3656,R5);
not not701(N3666,in0);
not not702(N3667,R2);
not not703(N3668,R3);
not not704(N3669,R4);
not not705(N3680,in1);
not not706(N3681,R2);
not not707(N3682,R3);
not not708(N3683,R4);
not not709(N3694,in2);
not not710(N3695,R0);
not not711(N3696,R1);
not not712(N3697,R3);
not not713(N3698,R5);
not not714(N3708,in2);
not not715(N3709,R0);
not not716(N3710,R1);
not not717(N3711,R3);
not not718(N3712,R5);
not not719(N3722,in1);
not not720(N3723,R3);
not not721(N3724,R4);
not not722(N3725,R5);
not not723(N3736,in0);
not not724(N3737,in1);
not not725(N3738,in2);
not not726(N3739,R2);
not not727(N3740,R4);
not not728(N3750,in0);
not not729(N3751,in1);
not not730(N3752,R0);
not not731(N3753,R4);
not not732(N3754,R5);
not not733(N3764,R1);
not not734(N3765,R2);
not not735(N3766,R4);
not not736(N3767,R5);
not not737(N3778,in2);
not not738(N3779,R1);
not not739(N3780,R4);
not not740(N3781,R5);
not not741(N3792,R0);
not not742(N3793,R1);
not not743(N3794,R2);
not not744(N3795,R3);
not not745(N3796,R5);
not not746(N3806,in0);
not not747(N3807,R0);
not not748(N3808,R2);
not not749(N3809,R4);
not not750(N3810,R5);
not not751(N3820,in0);
not not752(N3821,in2);
not not753(N3822,R2);
not not754(N3823,R3);
not not755(N3834,in0);
not not756(N3835,R1);
not not757(N3836,R3);
not not758(N3837,R5);
not not759(N3848,in2);
not not760(N3849,R0);
not not761(N3850,R2);
not not762(N3851,R3);
not not763(N3852,R5);
not not764(N3862,in0);
not not765(N3863,R0);
not not766(N3864,R2);
not not767(N3865,R4);
not not768(N3866,R5);
not not769(N3876,in0);
not not770(N3877,in1);
not not771(N3878,R2);
not not772(N3879,R4);
not not773(N3880,R5);
not not774(N3890,in2);
not not775(N3891,R0);
not not776(N3892,R5);
not not777(N3903,R0);
not not778(N3904,R1);
not not779(N3905,R5);
not not780(N3916,in2);
not not781(N3917,R4);
not not782(N3918,R5);
not not783(N3929,in1);
not not784(N3930,R2);
not not785(N3931,R5);
not not786(N3942,in0);
not not787(N3943,in1);
not not788(N3944,in2);
not not789(N3955,in1);
not not790(N3956,R2);
not not791(N3957,R5);
not not792(N3968,in0);
not not793(N3969,in1);
not not794(N3970,in2);
not not795(N3971,R2);
not not796(N3981,R0);
not not797(N3982,R1);
not not798(N3983,R3);
not not799(N3994,in2);
not not800(N3995,R0);
not not801(N3996,R1);
not not802(N3997,R4);
not not803(N4007,in1);
not not804(N4008,R0);
not not805(N4009,R4);
not not806(N4010,R5);
not not807(N4020,in1);
not not808(N4021,R3);
not not809(N4022,R5);
not not810(N4033,in1);
not not811(N4034,R2);
not not812(N4035,R3);
not not813(N4036,R4);
not not814(N4046,R0);
not not815(N4047,R3);
not not816(N4048,R5);
not not817(N4059,in2);
not not818(N4060,R3);
not not819(N4061,R4);
not not820(N4062,R5);
not not821(N4072,in1);
not not822(N4073,R0);
not not823(N4074,R1);
not not824(N4075,R4);
not not825(N4085,in0);
not not826(N4086,R0);
not not827(N4087,R1);
not not828(N4088,R4);
not not829(N4098,in1);
not not830(N4099,in2);
not not831(N4100,R0);
not not832(N4101,R1);
not not833(N4111,in1);
not not834(N4112,in2);
not not835(N4113,R0);
not not836(N4114,R2);
not not837(N4115,R4);
not not838(N4124,in1);
not not839(N4125,in2);
not not840(N4126,R1);
not not841(N4127,R3);
not not842(N4137,in1);
not not843(N4138,R0);
not not844(N4139,R3);
not not845(N4140,R4);
not not846(N4150,in1);
not not847(N4151,R0);
not not848(N4152,R3);
not not849(N4153,R4);
not not850(N4163,R1);
not not851(N4164,R2);
not not852(N4165,R3);
not not853(N4166,R5);
not not854(N4176,in1);
not not855(N4177,R2);
not not856(N4178,R3);
not not857(N4179,R5);
not not858(N4189,in1);
not not859(N4190,R0);
not not860(N4191,R2);
not not861(N4192,R5);
not not862(N4202,R0);
not not863(N4203,R1);
not not864(N4204,R2);
not not865(N4205,R5);
not not866(N4215,R0);
not not867(N4216,R1);
not not868(N4217,R2);
not not869(N4218,R5);
not not870(N4228,in0);
not not871(N4229,in1);
not not872(N4230,in2);
not not873(N4241,in0);
not not874(N4242,R0);
not not875(N4243,R2);
not not876(N4254,in1);
not not877(N4255,R1);
not not878(N4256,R5);
not not879(N4267,in0);
not not880(N4268,R1);
not not881(N4269,R2);
not not882(N4270,R4);
not not883(N4280,in0);
not not884(N4281,in2);
not not885(N4282,R2);
not not886(N4283,R3);
not not887(N4284,R5);
not not888(N4293,R0);
not not889(N4294,R1);
not not890(N4295,R2);
not not891(N4306,in1);
not not892(N4307,R0);
not not893(N4308,R1);
not not894(N4309,R4);
not not895(N4319,in1);
not not896(N4320,in2);
not not897(N4321,R1);
not not898(N4322,R4);
not not899(N4332,in0);
not not900(N4333,R0);
not not901(N4334,R1);
not not902(N4335,R3);
not not903(N4345,in0);
not not904(N4346,in1);
not not905(N4347,R2);
not not906(N4348,R5);
not not907(N4358,in0);
not not908(N4359,R4);
not not909(N4360,R5);
not not910(N4371,R1);
not not911(N4372,R4);
not not912(N4373,R5);
not not913(N4384,in2);
not not914(N4385,R0);
not not915(N4386,R3);
not not916(N4387,R4);
not not917(N4397,in2);
not not918(N4398,R1);
not not919(N4399,R5);
not not920(N4410,in0);
not not921(N4411,R0);
not not922(N4412,R2);
not not923(N4413,R5);
not not924(N4423,in2);
not not925(N4424,R0);
not not926(N4425,R2);
not not927(N4426,R3);
not not928(N4436,in1);
not not929(N4437,R0);
not not930(N4438,R4);
not not931(N4439,R5);
not not932(N4449,in0);
not not933(N4450,in2);
not not934(N4451,R4);
not not935(N4462,in1);
not not936(N4463,R1);
not not937(N4464,R3);
not not938(N4465,R4);
not not939(N4475,in0);
not not940(N4476,R2);
not not941(N4477,R3);
not not942(N4488,in1);
not not943(N4489,in2);
not not944(N4490,R4);
not not945(N4491,R5);
not not946(N4501,R1);
not not947(N4502,R4);
not not948(N4513,in1);
not not949(N4514,R1);
not not950(N4515,R5);
not not951(N4525,R0);
not not952(N4526,R4);
not not953(N4537,in2);
not not954(N4538,R2);
not not955(N4539,R4);
not not956(N4549,in0);
not not957(N4550,R3);
not not958(N4551,R5);
not not959(N4561,in1);
not not960(N4562,R2);
not not961(N4563,R4);
not not962(N4573,R0);
not not963(N4574,R1);
not not964(N4575,R4);
not not965(N4585,in0);
not not966(N4586,R0);
not not967(N4587,R5);
not not968(N4597,in1);
not not969(N4598,R1);
not not970(N4599,R2);
not not971(N4609,R0);
not not972(N4610,R4);
not not973(N4621,in2);
not not974(N4622,R1);
not not975(N4623,R4);
not not976(N4633,in1);
not not977(N4634,in2);
not not978(N4635,R1);
not not979(N4645,in1);
not not980(N4646,R3);
not not981(N4647,R4);
not not982(N4657,in2);
not not983(N4658,R3);
not not984(N4659,R4);
not not985(N4669,in1);
not not986(N4670,R4);
not not987(N4671,R5);
not not988(N4681,R0);
not not989(N4682,R2);
not not990(N4683,R3);
not not991(N4693,in2);
not not992(N4694,R0);
not not993(N4695,R4);
not not994(N4705,in1);
not not995(N4706,R3);
not not996(N4707,R4);
not not997(N4708,R5);
not not998(N4717,in2);
not not999(N4718,R1);
not not1000(N4719,R5);
not not1001(N4729,in0);
not not1002(N4730,in1);
not not1003(N4731,R3);
not not1004(N4741,R0);
not not1005(N4742,R3);
not not1006(N4743,R4);
not not1007(N4753,R0);
not not1008(N4754,R2);
not not1009(N4755,R3);
not not1010(N4765,in1);
not not1011(N4766,R1);
not not1012(N4767,R5);
not not1013(N4777,in0);
not not1014(N4778,R1);
not not1015(N4779,R3);
not not1016(N4789,in0);
not not1017(N4790,in2);
not not1018(N4801,in1);
not not1019(N4802,R2);
not not1020(N4813,R3);
not not1021(N4814,R5);
not not1022(N4825,in0);
not not1023(N4826,in1);
not not1024(N4827,R2);
not not1025(N4837,in1);
not not1026(N4838,in2);
not not1027(N4839,R4);
not not1028(N4849,R1);
not not1029(N4850,R2);
not not1030(N4851,R5);
not not1031(N4861,in1);
not not1032(N4862,R0);
not not1033(N4863,R2);
not not1034(N4864,R4);
not not1035(N4873,in2);
not not1036(N4874,R0);
not not1037(N4875,R2);
not not1038(N4876,R4);
not not1039(N4885,R2);
not not1040(N4886,R3);
not not1041(N4887,R5);
not not1042(N4897,in0);
not not1043(N4898,in1);
not not1044(N4899,in2);
not not1045(N4900,R4);
not not1046(N4909,R2);
not not1047(N4910,R4);
not not1048(N4921,in0);
not not1049(N4922,R0);
not not1050(N4923,R3);
not not1051(N4933,in2);
not not1052(N4934,R2);
not not1053(N4945,in2);
not not1054(N4946,R2);
not not1055(N4947,R3);
not not1056(N4957,in1);
not not1057(N4958,in2);
not not1058(N4959,R0);
not not1059(N4969,in0);
not not1060(N4970,R0);
not not1061(N4971,R1);
not not1062(N4981,R5);
not not1063(N4992,in1);
not not1064(N5003,R0);
not not1065(N5014,in0);
not not1066(N5015,R2);
not not1067(N5025,in2);
not not1068(N5026,R2);
not not1069(N5036,R0);
not not1070(N5037,R1);
not not1071(N5038,R5);
not not1072(N5047,in2);
not not1073(N5048,R4);
not not1074(N5058,R2);
not not1075(N5059,R5);
not not1076(N5069,in1);
not not1077(N5070,R0);
not not1078(N5071,R1);
not not1079(N5080,R1);
not not1080(N5081,R2);
not not1081(N5091,in2);
not not1082(N5092,R4);
not not1083(N5102,R0);
not not1084(N5113,R1);
not not1085(N5114,R4);
not not1086(N5124,in2);
not not1087(N5125,R4);
not not1088(N5126,R5);
not not1089(N5135,R1);
not not1090(N5136,R3);
not not1091(N5146,in1);
not not1092(N5147,R3);
not not1093(N5157,in2);
not not1094(N5158,R4);
not not1095(N5159,R5);
not not1096(N5168,R1);
not not1097(N5169,R2);
not not1098(N5179,in0);
not not1099(N5180,in1);
not not1100(N5181,R5);
not not1101(N5190,R3);
not not1102(N5200,in2);
not not1103(N5201,R1);
not not1104(N5210,R3);
not not1105(N5220,in1);
not not1106(N5221,in2);
not not1107(N5230,in2);
not not1108(N5231,R4);
not not1109(N5250,R4);
not not1110(N5251,R5);
not not1111(N5260,R4);
not not1112(N5269,in1);
not not1113(N5278,R1);
not not1114(N5286,R0);
not not1115(N5287,R2);
not not1116(N5288,R3);
not not1117(N5289,R4);
not not1118(N5290,R5);
not not1119(N5291,R6);
not not1120(N5292,R7);
not not1121(N5300,in1);
not not1122(N5301,R0);
not not1123(N5302,R2);
not not1124(N5303,R3);
not not1125(N5304,R5);
not not1126(N5305,R6);
not not1127(N5313,in1);
not not1128(N5314,in2);
not not1129(N5315,R3);
not not1130(N5316,R4);
not not1131(N5317,R5);
not not1132(N5318,R7);
not not1133(N5326,in1);
not not1134(N5327,R0);
not not1135(N5328,R3);
not not1136(N5329,R4);
not not1137(N5330,R5);
not not1138(N5338,R2);
not not1139(N5339,R3);
not not1140(N5340,R4);
not not1141(N5341,R5);
not not1142(N5342,R6);
not not1143(N5350,R0);
not not1144(N5351,R2);
not not1145(N5352,R3);
not not1146(N5353,R6);
not not1147(N5354,R7);
not not1148(N5362,in1);
not not1149(N5363,R0);
not not1150(N5364,R2);
not not1151(N5365,R3);
not not1152(N5366,R5);
not not1153(N5374,R2);
not not1154(N5375,R3);
not not1155(N5376,R4);
not not1156(N5377,R7);
not not1157(N5385,R3);
not not1158(N5386,R4);
not not1159(N5387,R5);
not not1160(N5388,R7);
not not1161(N5396,in1);
not not1162(N5397,R1);
not not1163(N5398,R4);
not not1164(N5399,R5);
not not1165(N5407,in1);
not not1166(N5408,R0);
not not1167(N5409,R5);
not not1168(N5410,R6);
not not1169(N5418,R0);
not not1170(N5419,R3);
not not1171(N5420,R4);
not not1172(N5421,R5);
not not1173(N5429,in1);
not not1174(N5430,R3);
not not1175(N5431,R7);
not not1176(N5439,in1);
not not1177(N5440,R3);
not not1178(N5441,R6);
not not1179(N5449,R0);
not not1180(N5450,R5);
not not1181(N5451,R6);
not not1182(N5459,in1);
not not1183(N5460,R4);
not not1184(N5461,R5);
not not1185(N5469,R0);
not not1186(N5470,R3);
not not1187(N5478,R4);
not not1188(N5479,R7);
not not1189(N5487,R4);
not not1190(N5488,R7);
not not1191(N5496,R2);
not not1192(N401,R4);
not not1193(N402,R5);
not not1194(N403,R6);
not not1195(N404,R7);
not not1196(N419,R4);
not not1197(N420,R5);
not not1198(N421,R7);
not not1199(N437,R5);
not not1200(N438,R7);
not not1201(N453,R4);
not not1202(N454,R6);
not not1203(N455,R7);
not not1204(N470,R4);
not not1205(N471,R5);
not not1206(N472,R6);
not not1207(N487,R5);
not not1208(N488,R6);
not not1209(N503,R6);
not not1210(N504,R7);
not not1211(N518,R4);
not not1212(N519,R6);
not not1213(N520,R7);
not not1214(N534,R4);
not not1215(N535,R5);
not not1216(N536,R6);
not not1217(N550,R5);
not not1218(N551,R6);
not not1219(N552,R7);
not not1220(N565,R4);
not not1221(N566,R5);
not not1222(N567,R6);
not not1223(N568,R7);
not not1224(N582,R4);
not not1225(N583,R5);
not not1226(N584,R6);
not not1227(N598,R4);
not not1228(N599,R6);
not not1229(N600,R7);
not not1230(N614,R4);
not not1231(N615,R6);
not not1232(N616,R7);
not not1233(N629,R4);
not not1234(N630,R5);
not not1235(N631,R6);
not not1236(N632,R7);
not not1237(N647,R4);
not not1238(N648,R5);
not not1239(N663,R5);
not not1240(N664,R7);
not not1241(N679,R5);
not not1242(N680,R7);
not not1243(N693,R4);
not not1244(N694,R5);
not not1245(N695,R6);
not not1246(N696,R7);
not not1247(N711,R6);
not not1248(N712,R7);
not not1249(N726,R4);
not not1250(N727,R6);
not not1251(N728,R7);
not not1252(N743,R3);
not not1253(N744,R5);
not not1254(N757,R3);
not not1255(N758,R4);
not not1256(N759,R5);
not not1257(N760,R7);
not not1258(N775,R5);
not not1259(N776,R7);
not not1260(N789,R4);
not not1261(N790,R5);
not not1262(N791,R6);
not not1263(N792,R7);
not not1264(N806,R4);
not not1265(N807,R5);
not not1266(N808,R6);
not not1267(N821,R5);
not not1268(N822,R6);
not not1269(N823,R7);
not not1270(N836,R5);
not not1271(N837,R6);
not not1272(N838,R7);
not not1273(N852,R4);
not not1274(N853,R6);
not not1275(N867,R6);
not not1276(N868,R7);
not not1277(N882,R3);
not not1278(N883,R6);
not not1279(N897,R5);
not not1280(N898,R7);
not not1281(N911,R4);
not not1282(N912,R5);
not not1283(N913,R7);
not not1284(N927,R5);
not not1285(N928,R7);
not not1286(N942,R6);
not not1287(N943,R7);
not not1288(N957,R4);
not not1289(N958,R5);
not not1290(N972,R4);
not not1291(N973,R5);
not not1292(N986,R4);
not not1293(N987,R5);
not not1294(N988,R7);
not not1295(N1002,R5);
not not1296(N1003,R7);
not not1297(N1016,R4);
not not1298(N1017,R5);
not not1299(N1018,R7);
not not1300(N1031,R4);
not not1301(N1032,R5);
not not1302(N1033,R6);
not not1303(N1046,R4);
not not1304(N1047,R5);
not not1305(N1048,R6);
not not1306(N1062,R4);
not not1307(N1063,R6);
not not1308(N1077,R4);
not not1309(N1078,R7);
not not1310(N1092,R4);
not not1311(N1093,R5);
not not1312(N1106,R4);
not not1313(N1107,R5);
not not1314(N1108,R7);
not not1315(N1122,R4);
not not1316(N1123,R7);
not not1317(N1137,R4);
not not1318(N1138,R6);
not not1319(N1151,R4);
not not1320(N1152,R5);
not not1321(N1153,R7);
not not1322(N1165,R4);
not not1323(N1166,R5);
not not1324(N1167,R6);
not not1325(N1168,R7);
not not1326(N1182,R4);
not not1327(N1183,R7);
not not1328(N1197,R4);
not not1329(N1198,R7);
not not1330(N1211,R4);
not not1331(N1212,R6);
not not1332(N1213,R7);
not not1333(N1226,R4);
not not1334(N1227,R6);
not not1335(N1228,R7);
not not1336(N1242,R5);
not not1337(N1243,R7);
not not1338(N1256,R4);
not not1339(N1257,R5);
not not1340(N1258,R6);
not not1341(N1273,R6);
not not1342(N1286,R3);
not not1343(N1287,R6);
not not1344(N1288,R7);
not not1345(N1301,R3);
not not1346(N1302,R5);
not not1347(N1303,R6);
not not1348(N1316,R4);
not not1349(N1317,R6);
not not1350(N1318,R7);
not not1351(N1331,R4);
not not1352(N1332,R6);
not not1353(N1333,R7);
not not1354(N1347,R5);
not not1355(N1348,R7);
not not1356(N1362,R5);
not not1357(N1363,R7);
not not1358(N1376,R3);
not not1359(N1377,R6);
not not1360(N1378,R7);
not not1361(N1392,R3);
not not1362(N1393,R6);
not not1363(N1406,R4);
not not1364(N1407,R6);
not not1365(N1408,R7);
not not1366(N1422,R5);
not not1367(N1423,R6);
not not1368(N1436,R4);
not not1369(N1437,R5);
not not1370(N1451,R5);
not not1371(N1463,R5);
not not1372(N1464,R6);
not not1373(N1465,R7);
not not1374(N1477,R5);
not not1375(N1478,R6);
not not1376(N1479,R7);
not not1377(N1490,R4);
not not1378(N1491,R5);
not not1379(N1492,R6);
not not1380(N1493,R7);
not not1381(N1507,R5);
not not1382(N1520,R5);
not not1383(N1521,R7);
not not1384(N1533,R4);
not not1385(N1534,R5);
not not1386(N1535,R6);
not not1387(N1547,R4);
not not1388(N1548,R5);
not not1389(N1549,R7);
not not1390(N1560,R3);
not not1391(N1561,R5);
not not1392(N1562,R6);
not not1393(N1563,R7);
not not1394(N1574,R4);
not not1395(N1575,R5);
not not1396(N1576,R6);
not not1397(N1577,R7);
not not1398(N1589,R5);
not not1399(N1590,R6);
not not1400(N1591,R7);
not not1401(N1603,R4);
not not1402(N1604,R6);
not not1403(N1605,R7);
not not1404(N1619,R5);
not not1405(N1632,R4);
not not1406(N1633,R7);
not not1407(N1645,R4);
not not1408(N1646,R6);
not not1409(N1647,R7);
not not1410(N1660,R4);
not not1411(N1661,R6);
not not1412(N1673,R4);
not not1413(N1674,R5);
not not1414(N1675,R7);
not not1415(N1688,R4);
not not1416(N1689,R6);
not not1417(N1702,R4);
not not1418(N1703,R7);
not not1419(N1716,R4);
not not1420(N1717,R5);
not not1421(N1730,R4);
not not1422(N1731,R5);
not not1423(N1744,R4);
not not1424(N1745,R5);
not not1425(N1759,R5);
not not1426(N1772,R6);
not not1427(N1773,R7);
not not1428(N1786,R4);
not not1429(N1787,R6);
not not1430(N1800,R3);
not not1431(N1801,R6);
not not1432(N1815,R7);
not not1433(N1828,R5);
not not1434(N1829,R7);
not not1435(N1843,R5);
not not1436(N1854,R3);
not not1437(N1855,R4);
not not1438(N1856,R6);
not not1439(N1857,R7);
not not1440(N1871,R5);
not not1441(N1883,R4);
not not1442(N1884,R5);
not not1443(N1885,R6);
not not1444(N1898,R3);
not not1445(N1899,R7);
not not1446(N1912,R5);
not not1447(N1913,R7);
not not1448(N1927,R5);
not not1449(N1941,R7);
not not1450(N1955,R6);
not not1451(N1969,R5);
not not1452(N1995,R4);
not not1453(N1996,R5);
not not1454(N1997,R6);
not not1455(N2009,R4);
not not1456(N2010,R5);
not not1457(N2011,R6);
not not1458(N2023,R4);
not not1459(N2024,R5);
not not1460(N2025,R6);
not not1461(N2038,R4);
not not1462(N2039,R6);
not not1463(N2052,R5);
not not1464(N2053,R6);
not not1465(N2065,R4);
not not1466(N2066,R5);
not not1467(N2067,R6);
not not1468(N2081,R5);
not not1469(N2093,R4);
not not1470(N2094,R6);
not not1471(N2095,R7);
not not1472(N2108,R6);
not not1473(N2109,R7);
not not1474(N2119,R4);
not not1475(N2120,R5);
not not1476(N2121,R6);
not not1477(N2122,R7);
not not1478(N2133,R5);
not not1479(N2134,R6);
not not1480(N2135,R7);
not not1481(N2146,R5);
not not1482(N2147,R6);
not not1483(N2148,R7);
not not1484(N2160,R4);
not not1485(N2161,R6);
not not1486(N2174,R6);
not not1487(N2186,R5);
not not1488(N2187,R7);
not not1489(N2199,R4);
not not1490(N2200,R5);
not not1491(N2212,R4);
not not1492(N2213,R6);
not not1493(N2225,R4);
not not1494(N2226,R6);
not not1495(N2238,R5);
not not1496(N2239,R7);
not not1497(N2250,R4);
not not1498(N2251,R5);
not not1499(N2252,R7);
not not1500(N2265,R7);
not not1501(N2278,R6);
not not1502(N2290,R4);
not not1503(N2291,R5);
not not1504(N2302,R4);
not not1505(N2303,R5);
not not1506(N2304,R6);
not not1507(N2316,R6);
not not1508(N2317,R7);
not not1509(N2329,R5);
not not1510(N2330,R7);
not not1511(N2343,R7);
not not1512(N2356,R7);
not not1513(N2368,R4);
not not1514(N2369,R6);
not not1515(N2382,R6);
not not1516(N2394,R4);
not not1517(N2395,R7);
not not1518(N2407,R6);
not not1519(N2408,R7);
not not1520(N2420,R5);
not not1521(N2421,R7);
not not1522(N2433,R5);
not not1523(N2434,R7);
not not1524(N2446,R5);
not not1525(N2447,R7);
not not1526(N2459,R5);
not not1527(N2460,R7);
not not1528(N2473,R6);
not not1529(N2486,R6);
not not1530(N2498,R5);
not not1531(N2499,R6);
not not1532(N2512,R3);
not not1533(N2524,R6);
not not1534(N2525,R7);
not not1535(N2536,R4);
not not1536(N2537,R5);
not not1537(N2538,R6);
not not1538(N2551,R6);
not not1539(N2564,R6);
not not1540(N2577,R3);
not not1541(N2589,R5);
not not1542(N2590,R6);
not not1543(N2603,R4);
not not1544(N2614,R4);
not not1545(N2615,R6);
not not1546(N2627,R4);
not not1547(N2638,R4);
not not1548(N2639,R5);
not not1549(N2650,R4);
not not1550(N2651,R7);
not not1551(N2662,R4);
not not1552(N2663,R5);
not not1553(N2674,R5);
not not1554(N2675,R6);
not not1555(N2687,R6);
not not1556(N2699,R6);
not not1557(N2710,R4);
not not1558(N2711,R6);
not not1559(N2723,R7);
not not1560(N2735,R6);
not not1561(N2747,R5);
not not1562(N2759,R5);
not not1563(N2771,R7);
not not1564(N2783,R5);
not not1565(N2794,R5);
not not1566(N2795,R6);
not not1567(N2806,R4);
not not1568(N2807,R6);
not not1569(N2818,R4);
not not1570(N2819,R5);
not not1571(N2831,R6);
not not1572(N2843,R6);
not not1573(N2867,R7);
not not1574(N2878,R3);
not not1575(N2879,R7);
not not1576(N2914,R5);
not not1577(N2915,R6);
not not1578(N2939,R5);
not not1579(N2951,R7);
not not1580(N2963,R3);
not not1581(N2975,R3);
not not1582(N2987,R7);
not not1583(N3011,R5);
not not1584(N3021,R4);
not not1585(N3022,R5);
not not1586(N3023,R6);
not not1587(N3035,R6);
not not1588(N3046,R6);
not not1589(N3047,R7);
not not1590(N3058,R6);
not not1591(N3059,R7);
not not1592(N3071,R5);
not not1593(N3082,R3);
not not1594(N3083,R4);
not not1595(N3094,R6);
not not1596(N3104,R4);
not not1597(N3105,R6);
not not1598(N3116,R6);
not not1599(N3127,R7);
not not1600(N3137,R5);
not not1601(N3138,R7);
not not1602(N3148,R5);
not not1603(N3149,R6);
not not1604(N3159,R4);
not not1605(N3160,R5);
not not1606(N3182,R7);
not not1607(N3193,R7);
not not1608(N3225,R3);
not not1609(N3226,R6);
not not1610(N3270,R6);
not not1611(N3271,R7);
not not1612(N3287,R7);
not not1613(N3302,R6);
not not1614(N3303,R7);
not not1615(N3318,R6);
not not1616(N3319,R7);
not not1617(N3334,R6);
not not1618(N3335,R7);
not not1619(N3350,R6);
not not1620(N3351,R7);
not not1621(N3367,R7);
not not1622(N3382,R6);
not not1623(N3396,R6);
not not1624(N3397,R7);
not not1625(N3411,R6);
not not1626(N3412,R7);
not not1627(N3426,R5);
not not1628(N3427,R6);
not not1629(N3442,R7);
not not1630(N3456,R6);
not not1631(N3457,R7);
not not1632(N3471,R6);
not not1633(N3472,R7);
not not1634(N3486,R5);
not not1635(N3487,R6);
not not1636(N3502,R6);
not not1637(N3516,R6);
not not1638(N3517,R7);
not not1639(N3531,R6);
not not1640(N3544,R6);
not not1641(N3545,R7);
not not1642(N3558,R6);
not not1643(N3559,R7);
not not1644(N3572,R6);
not not1645(N3573,R7);
not not1646(N3586,R5);
not not1647(N3587,R6);
not not1648(N3601,R6);
not not1649(N3614,R6);
not not1650(N3615,R7);
not not1651(N3629,R7);
not not1652(N3642,R6);
not not1653(N3643,R7);
not not1654(N3657,R7);
not not1655(N3670,R5);
not not1656(N3671,R6);
not not1657(N3684,R5);
not not1658(N3685,R6);
not not1659(N3699,R7);
not not1660(N3713,R7);
not not1661(N3726,R6);
not not1662(N3727,R7);
not not1663(N3741,R7);
not not1664(N3755,R6);
not not1665(N3768,R6);
not not1666(N3769,R7);
not not1667(N3782,R6);
not not1668(N3783,R7);
not not1669(N3797,R6);
not not1670(N3811,R7);
not not1671(N3824,R5);
not not1672(N3825,R6);
not not1673(N3838,R6);
not not1674(N3839,R7);
not not1675(N3853,R6);
not not1676(N3867,R6);
not not1677(N3881,R7);
not not1678(N3893,R6);
not not1679(N3894,R7);
not not1680(N3906,R6);
not not1681(N3907,R7);
not not1682(N3919,R6);
not not1683(N3920,R7);
not not1684(N3932,R6);
not not1685(N3933,R7);
not not1686(N3945,R5);
not not1687(N3946,R6);
not not1688(N3958,R6);
not not1689(N3959,R7);
not not1690(N3972,R4);
not not1691(N3984,R6);
not not1692(N3985,R7);
not not1693(N3998,R5);
not not1694(N4011,R7);
not not1695(N4023,R6);
not not1696(N4024,R7);
not not1697(N4037,R7);
not not1698(N4049,R6);
not not1699(N4050,R7);
not not1700(N4063,R7);
not not1701(N4076,R6);
not not1702(N4089,R6);
not not1703(N4102,R6);
not not1704(N4128,R6);
not not1705(N4141,R6);
not not1706(N4154,R6);
not not1707(N4167,R6);
not not1708(N4180,R7);
not not1709(N4193,R7);
not not1710(N4206,R6);
not not1711(N4219,R6);
not not1712(N4231,R6);
not not1713(N4232,R7);
not not1714(N4244,R6);
not not1715(N4245,R7);
not not1716(N4257,R6);
not not1717(N4258,R7);
not not1718(N4271,R7);
not not1719(N4296,R4);
not not1720(N4297,R6);
not not1721(N4310,R5);
not not1722(N4323,R6);
not not1723(N4336,R5);
not not1724(N4349,R6);
not not1725(N4361,R6);
not not1726(N4362,R7);
not not1727(N4374,R6);
not not1728(N4375,R7);
not not1729(N4388,R6);
not not1730(N4400,R6);
not not1731(N4401,R7);
not not1732(N4414,R6);
not not1733(N4427,R5);
not not1734(N4440,R6);
not not1735(N4452,R6);
not not1736(N4453,R7);
not not1737(N4466,R6);
not not1738(N4478,R4);
not not1739(N4479,R5);
not not1740(N4492,R6);
not not1741(N4503,R6);
not not1742(N4504,R7);
not not1743(N4516,R7);
not not1744(N4527,R6);
not not1745(N4528,R7);
not not1746(N4540,R7);
not not1747(N4552,R6);
not not1748(N4564,R7);
not not1749(N4576,R6);
not not1750(N4588,R7);
not not1751(N4600,R6);
not not1752(N4611,R6);
not not1753(N4612,R7);
not not1754(N4624,R7);
not not1755(N4636,R7);
not not1756(N4648,R6);
not not1757(N4660,R6);
not not1758(N4672,R7);
not not1759(N4684,R7);
not not1760(N4696,R6);
not not1761(N4720,R7);
not not1762(N4732,R5);
not not1763(N4744,R5);
not not1764(N4756,R5);
not not1765(N4768,R6);
not not1766(N4780,R6);
not not1767(N4791,R6);
not not1768(N4792,R7);
not not1769(N4803,R6);
not not1770(N4804,R7);
not not1771(N4815,R6);
not not1772(N4816,R7);
not not1773(N4828,R5);
not not1774(N4840,R7);
not not1775(N4852,R7);
not not1776(N4888,R7);
not not1777(N4911,R6);
not not1778(N4912,R7);
not not1779(N4924,R5);
not not1780(N4935,R6);
not not1781(N4936,R7);
not not1782(N4948,R6);
not not1783(N4960,R7);
not not1784(N4972,R5);
not not1785(N4982,R6);
not not1786(N4983,R7);
not not1787(N4993,R5);
not not1788(N4994,R6);
not not1789(N5004,R5);
not not1790(N5005,R6);
not not1791(N5016,R7);
not not1792(N5027,R6);
not not1793(N5049,R6);
not not1794(N5060,R6);
not not1795(N5082,R7);
not not1796(N5093,R7);
not not1797(N5103,R6);
not not1798(N5104,R7);
not not1799(N5115,R6);
not not1800(N5137,R6);
not not1801(N5148,R7);
not not1802(N5170,R6);
not not1803(N5191,R7);
not not1804(N5211,R7);
not not1805(N5240,R5);
not not1806(N5241,R7);
not not1807(N5940,in0);
not not1808(N5941,in2);
not not1809(N5942,R0);
not not1810(N5943,R2);
not not1811(N5944,R3);
not not1812(N5958,in0);
not not1813(N5959,in1);
not not1814(N5960,in2);
not not1815(N5961,R0);
not not1816(N5962,R1);
not not1817(N5976,in0);
not not1818(N5977,in1);
not not1819(N5978,in2);
not not1820(N5979,R0);
not not1821(N5980,R1);
not not1822(N5981,R2);
not not1823(N5994,in1);
not not1824(N5995,in2);
not not1825(N5996,R1);
not not1826(N5997,R2);
not not1827(N5998,R3);
not not1828(N6011,in0);
not not1829(N6012,in1);
not not1830(N6013,in2);
not not1831(N6014,R1);
not not1832(N6028,in0);
not not1833(N6029,in1);
not not1834(N6030,in2);
not not1835(N6031,R0);
not not1836(N6032,R1);
not not1837(N6033,R2);
not not1838(N6045,in1);
not not1839(N6046,in2);
not not1840(N6047,R0);
not not1841(N6048,R2);
not not1842(N6049,R3);
not not1843(N6062,in0);
not not1844(N6063,R0);
not not1845(N6064,R2);
not not1846(N6078,in1);
not not1847(N6079,in2);
not not1848(N6080,R1);
not not1849(N6081,R3);
not not1850(N6094,in2);
not not1851(N6095,R0);
not not1852(N6096,R1);
not not1853(N6097,R2);
not not1854(N6110,in0);
not not1855(N6111,in2);
not not1856(N6112,R0);
not not1857(N6113,R1);
not not1858(N6126,in1);
not not1859(N6127,in2);
not not1860(N6128,R1);
not not1861(N6129,R3);
not not1862(N6142,in1);
not not1863(N6143,R0);
not not1864(N6144,R3);
not not1865(N6158,in1);
not not1866(N6159,R0);
not not1867(N6160,R1);
not not1868(N6161,R3);
not not1869(N6174,in1);
not not1870(N6175,in2);
not not1871(N6176,R1);
not not1872(N6177,R2);
not not1873(N6190,in0);
not not1874(N6191,R0);
not not1875(N6192,R1);
not not1876(N6193,R2);
not not1877(N6194,R3);
not not1878(N6206,in1);
not not1879(N6207,in2);
not not1880(N6208,R0);
not not1881(N6209,R1);
not not1882(N6210,R2);
not not1883(N6222,in0);
not not1884(N6223,in2);
not not1885(N6224,R0);
not not1886(N6225,R1);
not not1887(N6226,R2);
not not1888(N6238,in0);
not not1889(N6239,in1);
not not1890(N6240,in2);
not not1891(N6241,R0);
not not1892(N6242,R3);
not not1893(N6254,in0);
not not1894(N6255,in2);
not not1895(N6256,R0);
not not1896(N6257,R1);
not not1897(N6258,R2);
not not1898(N6270,in0);
not not1899(N6271,R0);
not not1900(N6272,R1);
not not1901(N6273,R2);
not not1902(N6286,in0);
not not1903(N6287,in1);
not not1904(N6288,in2);
not not1905(N6289,R1);
not not1906(N6302,in0);
not not1907(N6303,R0);
not not1908(N6304,R1);
not not1909(N6317,in1);
not not1910(N6318,in2);
not not1911(N6332,in1);
not not1912(N6333,in2);
not not1913(N6334,R3);
not not1914(N6347,in0);
not not1915(N6348,in2);
not not1916(N6349,R0);
not not1917(N6350,R2);
not not1918(N6362,in0);
not not1919(N6363,in2);
not not1920(N6364,R1);
not not1921(N6365,R2);
not not1922(N6377,in0);
not not1923(N6378,in1);
not not1924(N6379,R0);
not not1925(N6380,R2);
not not1926(N6392,in0);
not not1927(N6393,in2);
not not1928(N6394,R0);
not not1929(N6395,R2);
not not1930(N6396,R3);
not not1931(N6407,in0);
not not1932(N6408,in1);
not not1933(N6409,in2);
not not1934(N6410,R0);
not not1935(N6422,in0);
not not1936(N6423,R2);
not not1937(N6424,R3);
not not1938(N6437,in1);
not not1939(N6438,R2);
not not1940(N6439,R3);
not not1941(N6452,in1);
not not1942(N6453,R0);
not not1943(N6454,R1);
not not1944(N6455,R2);
not not1945(N6467,in2);
not not1946(N6468,R0);
not not1947(N6469,R1);
not not1948(N6470,R2);
not not1949(N6482,in0);
not not1950(N6483,in1);
not not1951(N6484,in2);
not not1952(N6485,R0);
not not1953(N6486,R1);
not not1954(N6497,in0);
not not1955(N6498,in1);
not not1956(N6499,R0);
not not1957(N6500,R1);
not not1958(N6512,in2);
not not1959(N6513,R1);
not not1960(N6514,R3);
not not1961(N6527,in0);
not not1962(N6528,in1);
not not1963(N6529,in2);
not not1964(N6530,R1);
not not1965(N6531,R2);
not not1966(N6542,in0);
not not1967(N6543,R0);
not not1968(N6544,R2);
not not1969(N6557,in0);
not not1970(N6558,in2);
not not1971(N6559,R0);
not not1972(N6560,R1);
not not1973(N6572,in1);
not not1974(N6573,in2);
not not1975(N6574,R0);
not not1976(N6575,R1);
not not1977(N6576,R3);
not not1978(N6587,in2);
not not1979(N6588,R0);
not not1980(N6589,R3);
not not1981(N6602,R0);
not not1982(N6603,R1);
not not1983(N6604,R2);
not not1984(N6617,in0);
not not1985(N6618,R0);
not not1986(N6619,R2);
not not1987(N6632,in0);
not not1988(N6633,in1);
not not1989(N6634,R0);
not not1990(N6635,R1);
not not1991(N6647,in0);
not not1992(N6648,in1);
not not1993(N6649,R1);
not not1994(N6662,in1);
not not1995(N6663,in2);
not not1996(N6664,R2);
not not1997(N6665,R3);
not not1998(N6677,in0);
not not1999(N6678,in1);
not not2000(N6679,R0);
not not2001(N6680,R1);
not not2002(N6692,in0);
not not2003(N6693,in1);
not not2004(N6694,R0);
not not2005(N6707,in0);
not not2006(N6708,R0);
not not2007(N6721,in2);
not not2008(N6722,R1);
not not2009(N6723,R2);
not not2010(N6735,in1);
not not2011(N6736,R1);
not not2012(N6749,in1);
not not2013(N6750,R2);
not not2014(N6751,R3);
not not2015(N6763,in0);
not not2016(N6764,in2);
not not2017(N6765,R3);
not not2018(N6777,in1);
not not2019(N6778,R1);
not not2020(N6779,R2);
not not2021(N6791,in0);
not not2022(N6792,R0);
not not2023(N6793,R1);
not not2024(N6805,in0);
not not2025(N6806,in1);
not not2026(N6807,in2);
not not2027(N6808,R2);
not not2028(N6819,in0);
not not2029(N6820,R0);
not not2030(N6821,R2);
not not2031(N6833,in0);
not not2032(N6834,in2);
not not2033(N6835,R2);
not not2034(N6847,in0);
not not2035(N6848,in1);
not not2036(N6849,R2);
not not2037(N6861,in0);
not not2038(N6862,in2);
not not2039(N6863,R2);
not not2040(N6875,in1);
not not2041(N6889,R0);
not not2042(N6890,R1);
not not2043(N6903,R0);
not not2044(N6904,R3);
not not2045(N6917,in1);
not not2046(N6918,R0);
not not2047(N6931,R1);
not not2048(N6932,R2);
not not2049(N6933,R3);
not not2050(N6945,R0);
not not2051(N6946,R1);
not not2052(N6947,R2);
not not2053(N6959,R1);
not not2054(N6960,R3);
not not2055(N6973,in2);
not not2056(N6974,R1);
not not2057(N6975,R3);
not not2058(N6987,in0);
not not2059(N6988,in2);
not not2060(N6989,R1);
not not2061(N7001,in1);
not not2062(N7002,in2);
not not2063(N7003,R2);
not not2064(N7015,in1);
not not2065(N7016,R0);
not not2066(N7017,R2);
not not2067(N7029,in0);
not not2068(N7030,R2);
not not2069(N7031,R3);
not not2070(N7043,in2);
not not2071(N7044,R0);
not not2072(N7057,in2);
not not2073(N7058,R0);
not not2074(N7071,in2);
not not2075(N7072,R2);
not not2076(N7085,in0);
not not2077(N7086,in1);
not not2078(N7099,in0);
not not2079(N7100,in2);
not not2080(N7101,R2);
not not2081(N7113,in2);
not not2082(N7114,R1);
not not2083(N7115,R2);
not not2084(N7127,in0);
not not2085(N7140,in1);
not not2086(N7166,R3);
not not2087(N7179,R2);
not not2088(N7192,R1);
not not2089(N7205,in1);
not not2090(N7206,in2);
not not2091(N7218,in0);
not not2092(N7219,R0);
not not2093(N7231,in0);
not not2094(N7232,R0);
not not2095(N7233,R2);
not not2096(N7244,in1);
not not2097(N7245,in2);
not not2098(N7246,R2);
not not2099(N7257,in1);
not not2100(N7258,R1);
not not2101(N7259,R2);
not not2102(N7270,in2);
not not2103(N7271,R1);
not not2104(N7272,R2);
not not2105(N7283,in1);
not not2106(N7284,in2);
not not2107(N7285,R3);
not not2108(N7296,in0);
not not2109(N7297,in1);
not not2110(N7298,R3);
not not2111(N7309,in2);
not not2112(N7310,R0);
not not2113(N7322,in0);
not not2114(N7323,in1);
not not2115(N7324,in2);
not not2116(N7325,R2);
not not2117(N7335,in0);
not not2118(N7336,in1);
not not2119(N7337,R2);
not not2120(N7348,in1);
not not2121(N7349,R1);
not not2122(N7350,R3);
not not2123(N7361,in2);
not not2124(N7362,R1);
not not2125(N7363,R3);
not not2126(N7374,in1);
not not2127(N7375,in2);
not not2128(N7376,R1);
not not2129(N7387,in1);
not not2130(N7388,in2);
not not2131(N7389,R3);
not not2132(N7400,in0);
not not2133(N7401,in1);
not not2134(N7402,R3);
not not2135(N7413,in0);
not not2136(N7414,in2);
not not2137(N7415,R3);
not not2138(N7426,in1);
not not2139(N7427,R0);
not not2140(N7428,R3);
not not2141(N7439,R0);
not not2142(N7440,R1);
not not2143(N7441,R3);
not not2144(N7452,in0);
not not2145(N7453,in1);
not not2146(N7454,R1);
not not2147(N7465,in0);
not not2148(N7466,R1);
not not2149(N7478,in1);
not not2150(N7479,in2);
not not2151(N7480,R0);
not not2152(N7481,R2);
not not2153(N7491,in0);
not not2154(N7492,in2);
not not2155(N7493,R2);
not not2156(N7504,in0);
not not2157(N7505,R0);
not not2158(N7506,R3);
not not2159(N7517,in1);
not not2160(N7518,R0);
not not2161(N7519,R3);
not not2162(N7530,in0);
not not2163(N7543,R0);
not not2164(N7544,R1);
not not2165(N7556,R1);
not not2166(N7557,R2);
not not2167(N7569,in0);
not not2168(N7570,R2);
not not2169(N7582,R3);
not not2170(N7595,in0);
not not2171(N7596,in2);
not not2172(N7608,in0);
not not2173(N7609,R2);
not not2174(N7633,in0);
not not2175(N7634,R2);
not not2176(N7645,in1);
not not2177(N7646,R2);
not not2178(N7657,R2);
not not2179(N7669,in2);
not not2180(N7670,R2);
not not2181(N7681,in0);
not not2182(N7682,in2);
not not2183(N7693,R1);
not not2184(N7705,in0);
not not2185(N7706,R0);
not not2186(N7717,in1);
not not2187(N7718,R0);
not not2188(N7719,R1);
not not2189(N7729,R0);
not not2190(N7730,R2);
not not2191(N7741,in0);
not not2192(N7742,R2);
not not2193(N7753,in1);
not not2194(N7754,in2);
not not2195(N7765,in0);
not not2196(N7766,in2);
not not2197(N7777,in0);
not not2198(N7778,R2);
not not2199(N7789,in1);
not not2200(N7801,in1);
not not2201(N7802,R2);
not not2202(N7813,R2);
not not2203(N7825,in2);
not not2204(N7826,R0);
not not2205(N7827,R2);
not not2206(N7837,in0);
not not2207(N7838,in1);
not not2208(N7839,in2);
not not2209(N7849,in2);
not not2210(N7850,R0);
not not2211(N7861,in2);
not not2212(N7862,R0);
not not2213(N7873,in0);
not not2214(N7885,R3);
not not2215(N7897,in0);
not not2216(N7898,R1);
not not2217(N7909,in1);
not not2218(N7910,R2);
not not2219(N7920,R0);
not not2220(N7921,R3);
not not2221(N7942,in2);
not not2222(N7953,R1);
not not2223(N7975,R1);
not not2224(N7986,in2);
not not2225(N7997,R0);
not not2226(N8008,in1);
not not2227(N8019,in0);
not not2228(N8020,R1);
not not2229(N8030,R3);
not not2230(N8041,R2);
not not2231(N8051,in2);
not not2232(N8071,in0);
not not2233(N8091,in1);
not not2234(N8101,R1);
not not2235(N8129,in1);
not not2236(N8130,in2);
not not2237(N8131,R0);
not not2238(N8132,R1);
not not2239(N8133,R2);
not not2240(N8134,R3);
not not2241(N8135,R5);
not not2242(N8145,in0);
not not2243(N8146,in2);
not not2244(N8147,R0);
not not2245(N8148,R1);
not not2246(N8149,R2);
not not2247(N8150,R3);
not not2248(N8161,in0);
not not2249(N8162,R0);
not not2250(N8163,R1);
not not2251(N8164,R2);
not not2252(N8165,R3);
not not2253(N8176,in0);
not not2254(N8177,in1);
not not2255(N8178,in2);
not not2256(N8179,R1);
not not2257(N8180,R2);
not not2258(N8181,R4);
not not2259(N8191,in2);
not not2260(N8192,R0);
not not2261(N8193,R2);
not not2262(N8194,R4);
not not2263(N8195,R5);
not not2264(N8206,R0);
not not2265(N8207,R1);
not not2266(N8208,R2);
not not2267(N8209,R3);
not not2268(N8210,R4);
not not2269(N8221,R0);
not not2270(N8222,R1);
not not2271(N8223,R2);
not not2272(N8224,R3);
not not2273(N8225,R4);
not not2274(N8226,R5);
not not2275(N8236,in0);
not not2276(N8237,in2);
not not2277(N8238,R0);
not not2278(N8239,R2);
not not2279(N8240,R3);
not not2280(N8241,R4);
not not2281(N8251,in1);
not not2282(N8252,in2);
not not2283(N8253,R0);
not not2284(N8254,R2);
not not2285(N8255,R3);
not not2286(N8266,in0);
not not2287(N8267,R0);
not not2288(N8268,R1);
not not2289(N8269,R2);
not not2290(N8270,R3);
not not2291(N8281,in2);
not not2292(N8282,R0);
not not2293(N8283,R1);
not not2294(N8284,R3);
not not2295(N8285,R4);
not not2296(N8296,in0);
not not2297(N8297,in1);
not not2298(N8298,R2);
not not2299(N8299,R3);
not not2300(N8300,R4);
not not2301(N8301,R5);
not not2302(N8311,in0);
not not2303(N8312,in1);
not not2304(N8313,R1);
not not2305(N8314,R2);
not not2306(N8315,R3);
not not2307(N8326,in2);
not not2308(N8327,R0);
not not2309(N8328,R2);
not not2310(N8329,R4);
not not2311(N8330,R5);
not not2312(N8341,in1);
not not2313(N8342,in2);
not not2314(N8343,R1);
not not2315(N8344,R2);
not not2316(N8345,R4);
not not2317(N8356,in1);
not not2318(N8357,in2);
not not2319(N8358,R1);
not not2320(N8359,R2);
not not2321(N8360,R3);
not not2322(N8361,R5);
not not2323(N8371,in1);
not not2324(N8372,R0);
not not2325(N8373,R1);
not not2326(N8374,R3);
not not2327(N8385,in1);
not not2328(N8386,R0);
not not2329(N8387,R1);
not not2330(N8388,R2);
not not2331(N8389,R5);
not not2332(N8399,R0);
not not2333(N8400,R1);
not not2334(N8401,R2);
not not2335(N8402,R3);
not not2336(N8403,R5);
not not2337(N8413,R0);
not not2338(N8414,R1);
not not2339(N8415,R2);
not not2340(N8416,R3);
not not2341(N8417,R5);
not not2342(N8427,in2);
not not2343(N8428,R0);
not not2344(N8429,R1);
not not2345(N8430,R5);
not not2346(N8441,in1);
not not2347(N8442,in2);
not not2348(N8443,R0);
not not2349(N8444,R5);
not not2350(N8455,in0);
not not2351(N8456,R0);
not not2352(N8457,R1);
not not2353(N8458,R4);
not not2354(N8459,R5);
not not2355(N8469,in1);
not not2356(N8470,in2);
not not2357(N8471,R2);
not not2358(N8472,R3);
not not2359(N8473,R4);
not not2360(N8483,in1);
not not2361(N8484,R0);
not not2362(N8485,R1);
not not2363(N8486,R4);
not not2364(N8497,in0);
not not2365(N8498,in1);
not not2366(N8499,R0);
not not2367(N8500,R2);
not not2368(N8501,R3);
not not2369(N8511,in0);
not not2370(N8512,in2);
not not2371(N8513,R4);
not not2372(N8514,R5);
not not2373(N8525,in1);
not not2374(N8526,R2);
not not2375(N8527,R4);
not not2376(N8528,R5);
not not2377(N8539,in0);
not not2378(N8540,in1);
not not2379(N8541,R1);
not not2380(N8542,R4);
not not2381(N8543,R5);
not not2382(N8553,R0);
not not2383(N8554,R1);
not not2384(N8555,R2);
not not2385(N8556,R3);
not not2386(N8557,R5);
not not2387(N8567,in0);
not not2388(N8568,in2);
not not2389(N8569,R1);
not not2390(N8570,R3);
not not2391(N8571,R5);
not not2392(N8581,in0);
not not2393(N8582,in1);
not not2394(N8583,R1);
not not2395(N8584,R3);
not not2396(N8585,R5);
not not2397(N8595,in1);
not not2398(N8596,R1);
not not2399(N8597,R3);
not not2400(N8598,R4);
not not2401(N8609,in0);
not not2402(N8610,R3);
not not2403(N8611,R4);
not not2404(N8612,R5);
not not2405(N8623,in2);
not not2406(N8624,R3);
not not2407(N8625,R4);
not not2408(N8626,R5);
not not2409(N8637,in1);
not not2410(N8638,R1);
not not2411(N8639,R2);
not not2412(N8640,R3);
not not2413(N8651,in0);
not not2414(N8652,in2);
not not2415(N8653,R0);
not not2416(N8654,R2);
not not2417(N8655,R4);
not not2418(N8665,in0);
not not2419(N8666,in1);
not not2420(N8667,R0);
not not2421(N8668,R2);
not not2422(N8669,R4);
not not2423(N8679,in1);
not not2424(N8680,in2);
not not2425(N8681,R1);
not not2426(N8682,R2);
not not2427(N8683,R4);
not not2428(N8693,in1);
not not2429(N8694,R1);
not not2430(N8695,R2);
not not2431(N8696,R4);
not not2432(N8707,in1);
not not2433(N8708,R0);
not not2434(N8709,R1);
not not2435(N8710,R3);
not not2436(N8721,in0);
not not2437(N8722,R1);
not not2438(N8723,R2);
not not2439(N8724,R3);
not not2440(N8725,R5);
not not2441(N8735,in1);
not not2442(N8736,in2);
not not2443(N8737,R2);
not not2444(N8738,R5);
not not2445(N8749,in0);
not not2446(N8750,in1);
not not2447(N8751,R0);
not not2448(N8752,R3);
not not2449(N8753,R5);
not not2450(N8763,in2);
not not2451(N8764,R0);
not not2452(N8765,R2);
not not2453(N8766,R4);
not not2454(N8767,R5);
not not2455(N8777,in0);
not not2456(N8778,in1);
not not2457(N8779,R0);
not not2458(N8780,R3);
not not2459(N8781,R5);
not not2460(N8791,in1);
not not2461(N8792,in2);
not not2462(N8793,R2);
not not2463(N8794,R4);
not not2464(N8795,R5);
not not2465(N8805,R1);
not not2466(N8806,R2);
not not2467(N8807,R3);
not not2468(N8808,R4);
not not2469(N8819,in1);
not not2470(N8820,in2);
not not2471(N8821,R0);
not not2472(N8822,R1);
not not2473(N8823,R3);
not not2474(N8833,in0);
not not2475(N8834,in2);
not not2476(N8835,R3);
not not2477(N8836,R4);
not not2478(N8847,in0);
not not2479(N8848,R1);
not not2480(N8849,R4);
not not2481(N8850,R5);
not not2482(N8861,in1);
not not2483(N8862,in2);
not not2484(N8863,R1);
not not2485(N8864,R5);
not not2486(N8875,R0);
not not2487(N8876,R1);
not not2488(N8877,R3);
not not2489(N8878,R4);
not not2490(N8889,in1);
not not2491(N8890,in2);
not not2492(N8891,R0);
not not2493(N8892,R2);
not not2494(N8893,R5);
not not2495(N8903,R0);
not not2496(N8904,R4);
not not2497(N8905,R5);
not not2498(N8916,in2);
not not2499(N8917,R0);
not not2500(N8918,R2);
not not2501(N8919,R4);
not not2502(N8920,R5);
not not2503(N8929,in1);
not not2504(N8930,R0);
not not2505(N8931,R2);
not not2506(N8942,in2);
not not2507(N8943,R2);
not not2508(N8944,R3);
not not2509(N8945,R5);
not not2510(N8955,in1);
not not2511(N8956,R0);
not not2512(N8957,R5);
not not2513(N8968,R0);
not not2514(N8969,R2);
not not2515(N8970,R5);
not not2516(N8981,R0);
not not2517(N8982,R1);
not not2518(N8983,R2);
not not2519(N8994,in0);
not not2520(N8995,in1);
not not2521(N8996,R1);
not not2522(N8997,R4);
not not2523(N9007,in2);
not not2524(N9008,R0);
not not2525(N9009,R2);
not not2526(N9010,R3);
not not2527(N9011,R5);
not not2528(N9020,R2);
not not2529(N9021,R4);
not not2530(N9022,R5);
not not2531(N9033,in1);
not not2532(N9034,R0);
not not2533(N9035,R2);
not not2534(N9036,R3);
not not2535(N9046,in0);
not not2536(N9047,R2);
not not2537(N9048,R4);
not not2538(N9049,R5);
not not2539(N9059,R1);
not not2540(N9060,R3);
not not2541(N9061,R4);
not not2542(N9062,R5);
not not2543(N9072,R1);
not not2544(N9073,R3);
not not2545(N9074,R4);
not not2546(N9075,R5);
not not2547(N9085,in1);
not not2548(N9086,in2);
not not2549(N9087,R3);
not not2550(N9088,R4);
not not2551(N9089,R5);
not not2552(N9098,in1);
not not2553(N9099,in2);
not not2554(N9100,R0);
not not2555(N9101,R4);
not not2556(N9111,in1);
not not2557(N9112,R0);
not not2558(N9113,R3);
not not2559(N9114,R4);
not not2560(N9124,R0);
not not2561(N9125,R1);
not not2562(N9126,R3);
not not2563(N9127,R5);
not not2564(N9137,in2);
not not2565(N9138,R1);
not not2566(N9139,R2);
not not2567(N9140,R5);
not not2568(N9150,in2);
not not2569(N9151,R0);
not not2570(N9152,R2);
not not2571(N9153,R5);
not not2572(N9163,in1);
not not2573(N9164,R0);
not not2574(N9165,R2);
not not2575(N9166,R5);
not not2576(N9176,in2);
not not2577(N9177,R0);
not not2578(N9178,R2);
not not2579(N9179,R4);
not not2580(N9189,R0);
not not2581(N9190,R2);
not not2582(N9191,R3);
not not2583(N9202,in1);
not not2584(N9203,R0);
not not2585(N9204,R3);
not not2586(N9215,in2);
not not2587(N9216,R0);
not not2588(N9217,R2);
not not2589(N9228,in0);
not not2590(N9229,R1);
not not2591(N9230,R2);
not not2592(N9231,R4);
not not2593(N9241,in1);
not not2594(N9242,in2);
not not2595(N9243,R2);
not not2596(N9244,R3);
not not2597(N9254,R2);
not not2598(N9255,R3);
not not2599(N9256,R5);
not not2600(N9267,R2);
not not2601(N9268,R3);
not not2602(N9269,R5);
not not2603(N9280,in0);
not not2604(N9281,in1);
not not2605(N9282,R0);
not not2606(N9283,R5);
not not2607(N9293,in0);
not not2608(N9294,R1);
not not2609(N9295,R2);
not not2610(N9296,R4);
not not2611(N9306,R1);
not not2612(N9307,R2);
not not2613(N9308,R4);
not not2614(N9309,R5);
not not2615(N9319,R1);
not not2616(N9320,R2);
not not2617(N9321,R4);
not not2618(N9322,R5);
not not2619(N9332,in1);
not not2620(N9333,in2);
not not2621(N9334,R2);
not not2622(N9335,R3);
not not2623(N9336,R5);
not not2624(N9345,in1);
not not2625(N9346,in2);
not not2626(N9347,R2);
not not2627(N9348,R3);
not not2628(N9358,in0);
not not2629(N9359,R1);
not not2630(N9360,R3);
not not2631(N9371,R1);
not not2632(N9372,R2);
not not2633(N9373,R3);
not not2634(N9384,R1);
not not2635(N9385,R2);
not not2636(N9386,R3);
not not2637(N9397,in0);
not not2638(N9398,in2);
not not2639(N9399,R0);
not not2640(N9400,R5);
not not2641(N9410,in0);
not not2642(N9411,R0);
not not2643(N9412,R1);
not not2644(N9413,R4);
not not2645(N9423,in1);
not not2646(N9424,R0);
not not2647(N9425,R1);
not not2648(N9426,R4);
not not2649(N9436,in0);
not not2650(N9437,in1);
not not2651(N9438,R4);
not not2652(N9449,in0);
not not2653(N9450,R1);
not not2654(N9451,R3);
not not2655(N9452,R4);
not not2656(N9462,in0);
not not2657(N9463,in1);
not not2658(N9464,R3);
not not2659(N9465,R4);
not not2660(N9475,in0);
not not2661(N9476,in1);
not not2662(N9477,R3);
not not2663(N9478,R5);
not not2664(N9488,in2);
not not2665(N9489,R1);
not not2666(N9490,R2);
not not2667(N9501,in0);
not not2668(N9502,in2);
not not2669(N9503,R0);
not not2670(N9504,R1);
not not2671(N9514,in1);
not not2672(N9515,R4);
not not2673(N9516,R5);
not not2674(N9527,R0);
not not2675(N9528,R1);
not not2676(N9529,R5);
not not2677(N9540,in0);
not not2678(N9541,in1);
not not2679(N9542,R0);
not not2680(N9543,R3);
not not2681(N9553,R3);
not not2682(N9554,R4);
not not2683(N9555,R5);
not not2684(N9566,in0);
not not2685(N9567,in2);
not not2686(N9568,R0);
not not2687(N9569,R2);
not not2688(N9579,in2);
not not2689(N9580,R2);
not not2690(N9581,R5);
not not2691(N9592,in1);
not not2692(N9593,R2);
not not2693(N9594,R3);
not not2694(N9605,in0);
not not2695(N9606,R0);
not not2696(N9607,R2);
not not2697(N9608,R3);
not not2698(N9618,in1);
not not2699(N9619,in2);
not not2700(N9620,R2);
not not2701(N9621,R4);
not not2702(N9631,in0);
not not2703(N9632,in1);
not not2704(N9633,R1);
not not2705(N9634,R2);
not not2706(N9644,R1);
not not2707(N9645,R3);
not not2708(N9646,R5);
not not2709(N9656,in0);
not not2710(N9657,in1);
not not2711(N9658,R1);
not not2712(N9668,R2);
not not2713(N9669,R3);
not not2714(N9670,R4);
not not2715(N9680,in0);
not not2716(N9681,R0);
not not2717(N9682,R1);
not not2718(N9692,in1);
not not2719(N9693,in2);
not not2720(N9694,R0);
not not2721(N9704,in1);
not not2722(N9705,in2);
not not2723(N9706,R5);
not not2724(N9716,R0);
not not2725(N9717,R3);
not not2726(N9718,R4);
not not2727(N9728,R1);
not not2728(N9729,R2);
not not2729(N9730,R4);
not not2730(N9740,in2);
not not2731(N9741,R0);
not not2732(N9742,R4);
not not2733(N9752,in2);
not not2734(N9753,R1);
not not2735(N9754,R4);
not not2736(N9755,R5);
not not2737(N9764,in1);
not not2738(N9765,R0);
not not2739(N9766,R1);
not not2740(N9776,in0);
not not2741(N9777,R0);
not not2742(N9778,R4);
not not2743(N9788,in1);
not not2744(N9789,R0);
not not2745(N9790,R2);
not not2746(N9791,R4);
not not2747(N9800,R0);
not not2748(N9801,R2);
not not2749(N9802,R4);
not not2750(N9812,in1);
not not2751(N9813,R2);
not not2752(N9814,R4);
not not2753(N9824,R1);
not not2754(N9825,R3);
not not2755(N9836,in1);
not not2756(N9837,R0);
not not2757(N9838,R1);
not not2758(N9839,R5);
not not2759(N9848,in0);
not not2760(N9849,R2);
not not2761(N9850,R3);
not not2762(N9860,in1);
not not2763(N9861,R2);
not not2764(N9872,in1);
not not2765(N9873,in2);
not not2766(N9874,R3);
not not2767(N9884,in2);
not not2768(N9885,R0);
not not2769(N9886,R5);
not not2770(N9896,in2);
not not2771(N9897,R0);
not not2772(N9898,R3);
not not2773(N9899,R5);
not not2774(N9908,R0);
not not2775(N9909,R1);
not not2776(N9910,R4);
not not2777(N9911,R5);
not not2778(N9920,R0);
not not2779(N9921,R4);
not not2780(N9922,R5);
not not2781(N9932,R0);
not not2782(N9933,R4);
not not2783(N9934,R5);
not not2784(N9944,in1);
not not2785(N9945,R1);
not not2786(N9946,R5);
not not2787(N9956,R1);
not not2788(N9957,R4);
not not2789(N9958,R5);
not not2790(N9968,R2);
not not2791(N9969,R4);
not not2792(N9970,R5);
not not2793(N9980,in0);
not not2794(N9981,R1);
not not2795(N9982,R3);
not not2796(N9992,in1);
not not2797(N9993,R1);
not not2798(N9994,R3);
not not2799(N10004,in1);
not not2800(N10005,R4);
not not2801(N10006,R5);
not not2802(N10016,in1);
not not2803(N10017,in2);
not not2804(N10018,R0);
not not2805(N10019,R3);
not not2806(N10028,in1);
not not2807(N10029,R1);
not not2808(N10030,R3);
not not2809(N10040,R0);
not not2810(N10041,R1);
not not2811(N10042,R3);
not not2812(N10052,in1);
not not2813(N10053,R1);
not not2814(N10054,R3);
not not2815(N10064,R0);
not not2816(N10065,R1);
not not2817(N10066,R3);
not not2818(N10076,in1);
not not2819(N10077,in2);
not not2820(N10078,R2);
not not2821(N10088,R0);
not not2822(N10089,R1);
not not2823(N10090,R5);
not not2824(N10100,R0);
not not2825(N10101,R2);
not not2826(N10102,R3);
not not2827(N10112,R1);
not not2828(N10113,R2);
not not2829(N10114,R4);
not not2830(N10124,in1);
not not2831(N10125,R3);
not not2832(N10126,R4);
not not2833(N10127,R5);
not not2834(N10136,in2);
not not2835(N10137,R3);
not not2836(N10138,R4);
not not2837(N10139,R5);
not not2838(N10148,in1);
not not2839(N10149,R3);
not not2840(N10150,R5);
not not2841(N10160,R0);
not not2842(N10161,R2);
not not2843(N10162,R5);
not not2844(N10172,R0);
not not2845(N10173,R1);
not not2846(N10174,R4);
not not2847(N10184,in1);
not not2848(N10185,R4);
not not2849(N10196,in0);
not not2850(N10197,R0);
not not2851(N10198,R1);
not not2852(N10208,in2);
not not2853(N10219,in1);
not not2854(N10220,R0);
not not2855(N10230,R2);
not not2856(N10241,R0);
not not2857(N10242,R2);
not not2858(N10243,R5);
not not2859(N10252,R2);
not not2860(N10253,R4);
not not2861(N10263,in2);
not not2862(N10264,R2);
not not2863(N10274,in0);
not not2864(N10275,in2);
not not2865(N10276,R1);
not not2866(N10285,R0);
not not2867(N10286,R4);
not not2868(N10296,R1);
not not2869(N10297,R2);
not not2870(N10307,R0);
not not2871(N10318,in0);
not not2872(N10319,R3);
not not2873(N10329,R0);
not not2874(N10330,R2);
not not2875(N10340,R1);
not not2876(N10341,R2);
not not2877(N10351,R1);
not not2878(N10352,R5);
not not2879(N10362,in0);
not not2880(N10363,R5);
not not2881(N10373,in1);
not not2882(N10374,R0);
not not2883(N10384,R0);
not not2884(N10385,R5);
not not2885(N10395,R0);
not not2886(N10396,R5);
not not2887(N10406,R0);
not not2888(N10407,R3);
not not2889(N10417,in2);
not not2890(N10418,R0);
not not2891(N10419,R4);
not not2892(N10428,R2);
not not2893(N10429,R3);
not not2894(N10430,R5);
not not2895(N10439,R2);
not not2896(N10440,R3);
not not2897(N10441,R5);
not not2898(N10450,R2);
not not2899(N10451,R3);
not not2900(N10461,R2);
not not2901(N10462,R3);
not not2902(N10472,R2);
not not2903(N10473,R3);
not not2904(N10483,in1);
not not2905(N10484,in2);
not not2906(N10494,in1);
not not2907(N10495,R0);
not not2908(N10505,R2);
not not2909(N10516,R0);
not not2910(N10517,R3);
not not2911(N10527,in2);
not not2912(N10538,in1);
not not2913(N10539,R3);
not not2914(N10549,in2);
not not2915(N10560,in2);
not not2916(N10561,R1);
not not2917(N10571,R0);
not not2918(N10572,R1);
not not2919(N10582,R3);
not not2920(N10583,R4);
not not2921(N10593,in0);
not not2922(N10594,R2);
not not2923(N10604,R1);
not not2924(N10605,R3);
not not2925(N10615,in1);
not not2926(N10616,R0);
not not2927(N10617,R4);
not not2928(N10626,in1);
not not2929(N10627,R0);
not not2930(N10628,R2);
not not2931(N10637,in2);
not not2932(N10638,R0);
not not2933(N10648,in0);
not not2934(N10649,R2);
not not2935(N10659,in2);
not not2936(N10660,R2);
not not2937(N10670,R0);
not not2938(N10671,R4);
not not2939(N10681,R5);
not not2940(N10691,R4);
not not2941(N10692,R5);
not not2942(N10701,R3);
not not2943(N10711,in1);
not not2944(N10712,R5);
not not2945(N10721,in2);
not not2946(N10722,R5);
not not2947(N10731,in1);
not not2948(N10741,R5);
not not2949(N10751,in2);
not not2950(N10752,R1);
not not2951(N10761,R1);
not not2952(N10762,R5);
not not2953(N10771,in1);
not not2954(N10781,R3);
not not2955(N10791,in1);
not not2956(N10792,R3);
not not2957(N10801,in2);
not not2958(N10802,R0);
not not2959(N10811,in2);
not not2960(N10812,R0);
not not2961(N10821,in1);
not not2962(N10831,in1);
not not2963(N10832,R3);
not not2964(N10841,in0);
not not2965(N10842,R3);
not not2966(N10851,in1);
not not2967(N10852,R3);
not not2968(N10861,in1);
not not2969(N10862,R1);
not not2970(N10871,in1);
not not2971(N10872,in2);
not not2972(N10881,in2);
not not2973(N10891,R0);
not not2974(N10901,R3);
not not2975(N10911,R2);
not not2976(N10912,R5);
not not2977(N10931,R0);
not not2978(N10940,R1);
not not2979(N10949,R3);
not not2980(N10958,R3);
not not2981(N10967,R2);
not not2982(N10975,in1);
not not2983(N10976,in2);
not not2984(N10977,R2);
not not2985(N10978,R5);
not not2986(N10979,R6);
not not2987(N10980,R7);
not not2988(N10988,R0);
not not2989(N10989,R1);
not not2990(N10990,R2);
not not2991(N10991,R3);
not not2992(N10992,R6);
not not2993(N10993,R7);
not not2994(N11001,R1);
not not2995(N11002,R2);
not not2996(N11003,R3);
not not2997(N11004,R4);
not not2998(N11005,R6);
not not2999(N11006,R7);
not not3000(N11014,in2);
not not3001(N11015,R0);
not not3002(N11016,R5);
not not3003(N11017,R6);
not not3004(N11018,R7);
not not3005(N11026,in2);
not not3006(N11027,R0);
not not3007(N11028,R3);
not not3008(N11029,R6);
not not3009(N11030,R7);
not not3010(N11038,R1);
not not3011(N11039,R3);
not not3012(N11040,R4);
not not3013(N11041,R5);
not not3014(N11042,R6);
not not3015(N11050,R2);
not not3016(N11051,R3);
not not3017(N11052,R4);
not not3018(N11053,R5);
not not3019(N11054,R6);
not not3020(N11062,R2);
not not3021(N11063,R3);
not not3022(N11064,R4);
not not3023(N11065,R5);
not not3024(N11066,R6);
not not3025(N11074,R0);
not not3026(N11075,R1);
not not3027(N11076,R3);
not not3028(N11077,R5);
not not3029(N11078,R7);
not not3030(N11086,in1);
not not3031(N11087,in2);
not not3032(N11088,R0);
not not3033(N11089,R5);
not not3034(N11090,R6);
not not3035(N11098,in1);
not not3036(N11099,in2);
not not3037(N11100,R1);
not not3038(N11101,R4);
not not3039(N11102,R6);
not not3040(N11110,in0);
not not3041(N11111,in1);
not not3042(N11112,in2);
not not3043(N11113,R1);
not not3044(N11114,R6);
not not3045(N11122,R1);
not not3046(N11123,R4);
not not3047(N11124,R5);
not not3048(N11125,R7);
not not3049(N11133,in2);
not not3050(N11134,R3);
not not3051(N11135,R4);
not not3052(N11136,R6);
not not3053(N11144,R2);
not not3054(N11145,R4);
not not3055(N11146,R5);
not not3056(N11147,R7);
not not3057(N11155,in1);
not not3058(N11156,R1);
not not3059(N11157,R4);
not not3060(N11158,R5);
not not3061(N11166,R0);
not not3062(N11167,R3);
not not3063(N11168,R4);
not not3064(N11169,R6);
not not3065(N11177,R1);
not not3066(N11178,R2);
not not3067(N11179,R4);
not not3068(N11180,R7);
not not3069(N11188,R1);
not not3070(N11189,R2);
not not3071(N11190,R4);
not not3072(N11191,R7);
not not3073(N11199,in1);
not not3074(N11200,R0);
not not3075(N11201,R4);
not not3076(N11202,R5);
not not3077(N11210,R0);
not not3078(N11211,R2);
not not3079(N11212,R4);
not not3080(N11213,R5);
not not3081(N11221,in1);
not not3082(N11222,R1);
not not3083(N11223,R5);
not not3084(N11224,R7);
not not3085(N11232,in2);
not not3086(N11233,R4);
not not3087(N11234,R6);
not not3088(N11235,R7);
not not3089(N11243,R0);
not not3090(N11244,R3);
not not3091(N11245,R6);
not not3092(N11246,R7);
not not3093(N11254,in1);
not not3094(N11255,R3);
not not3095(N11256,R4);
not not3096(N11257,R6);
not not3097(N11265,in2);
not not3098(N11266,R0);
not not3099(N11267,R5);
not not3100(N11268,R6);
not not3101(N11276,in1);
not not3102(N11277,R2);
not not3103(N11278,R4);
not not3104(N11286,in1);
not not3105(N11287,R1);
not not3106(N11288,R7);
not not3107(N11296,R3);
not not3108(N11297,R4);
not not3109(N11298,R7);
not not3110(N11306,R0);
not not3111(N11307,R1);
not not3112(N11308,R6);
not not3113(N11316,R0);
not not3114(N11317,R1);
not not3115(N11318,R5);
not not3116(N11326,R0);
not not3117(N11327,R1);
not not3118(N11328,R5);
not not3119(N11336,in2);
not not3120(N11337,R3);
not not3121(N11338,R7);
not not3122(N11346,R1);
not not3123(N11347,R4);
not not3124(N11348,R6);
not not3125(N11356,R1);
not not3126(N11357,R4);
not not3127(N11358,R6);
not not3128(N11366,R4);
not not3129(N11367,R5);
not not3130(N11368,R6);
not not3131(N11376,in2);
not not3132(N11377,R4);
not not3133(N11378,R7);
not not3134(N11386,in2);
not not3135(N11387,R1);
not not3136(N11388,R7);
not not3137(N11396,R0);
not not3138(N11397,R4);
not not3139(N11398,R5);
not not3140(N11406,R5);
not not3141(N11407,R6);
not not3142(N11414,in1);
not not3143(N11415,R0);
not not3144(N11416,R2);
not not3145(N11417,R4);
not not3146(N11418,R5);
not not3147(N11419,R7);
not not3148(N11426,R1);
not not3149(N11427,R4);
not not3150(N11428,R5);
not not3151(N11429,R7);
not not3152(N5945,R4);
not not3153(N5946,R5);
not not3154(N5947,R6);
not not3155(N5948,R7);
not not3156(N5963,R3);
not not3157(N5964,R5);
not not3158(N5965,R6);
not not3159(N5966,R7);
not not3160(N5982,R4);
not not3161(N5983,R5);
not not3162(N5984,R6);
not not3163(N5999,R4);
not not3164(N6000,R6);
not not3165(N6001,R7);
not not3166(N6015,R4);
not not3167(N6016,R5);
not not3168(N6017,R6);
not not3169(N6018,R7);
not not3170(N6034,R6);
not not3171(N6035,R7);
not not3172(N6050,R5);
not not3173(N6051,R6);
not not3174(N6052,R7);
not not3175(N6065,R4);
not not3176(N6066,R5);
not not3177(N6067,R6);
not not3178(N6068,R7);
not not3179(N6082,R4);
not not3180(N6083,R5);
not not3181(N6084,R7);
not not3182(N6098,R4);
not not3183(N6099,R5);
not not3184(N6100,R6);
not not3185(N6114,R5);
not not3186(N6115,R6);
not not3187(N6116,R7);
not not3188(N6130,R4);
not not3189(N6131,R5);
not not3190(N6132,R6);
not not3191(N6145,R4);
not not3192(N6146,R5);
not not3193(N6147,R6);
not not3194(N6148,R7);
not not3195(N6162,R4);
not not3196(N6163,R5);
not not3197(N6164,R6);
not not3198(N6178,R4);
not not3199(N6179,R5);
not not3200(N6180,R6);
not not3201(N6195,R5);
not not3202(N6196,R7);
not not3203(N6211,R5);
not not3204(N6212,R7);
not not3205(N6227,R5);
not not3206(N6228,R6);
not not3207(N6243,R4);
not not3208(N6244,R7);
not not3209(N6259,R4);
not not3210(N6260,R6);
not not3211(N6274,R5);
not not3212(N6275,R6);
not not3213(N6276,R7);
not not3214(N6290,R4);
not not3215(N6291,R5);
not not3216(N6292,R6);
not not3217(N6305,R5);
not not3218(N6306,R6);
not not3219(N6307,R7);
not not3220(N6319,R4);
not not3221(N6320,R5);
not not3222(N6321,R6);
not not3223(N6322,R7);
not not3224(N6335,R5);
not not3225(N6336,R6);
not not3226(N6337,R7);
not not3227(N6351,R6);
not not3228(N6352,R7);
not not3229(N6366,R5);
not not3230(N6367,R7);
not not3231(N6381,R6);
not not3232(N6382,R7);
not not3233(N6397,R5);
not not3234(N6411,R4);
not not3235(N6412,R5);
not not3236(N6425,R4);
not not3237(N6426,R6);
not not3238(N6427,R7);
not not3239(N6440,R4);
not not3240(N6441,R6);
not not3241(N6442,R7);
not not3242(N6456,R4);
not not3243(N6457,R5);
not not3244(N6471,R4);
not not3245(N6472,R5);
not not3246(N6487,R7);
not not3247(N6501,R3);
not not3248(N6502,R6);
not not3249(N6515,R5);
not not3250(N6516,R6);
not not3251(N6517,R7);
not not3252(N6532,R5);
not not3253(N6545,R5);
not not3254(N6546,R6);
not not3255(N6547,R7);
not not3256(N6561,R4);
not not3257(N6562,R7);
not not3258(N6577,R5);
not not3259(N6590,R4);
not not3260(N6591,R5);
not not3261(N6592,R7);
not not3262(N6605,R4);
not not3263(N6606,R5);
not not3264(N6607,R6);
not not3265(N6620,R3);
not not3266(N6621,R4);
not not3267(N6622,R5);
not not3268(N6636,R4);
not not3269(N6637,R5);
not not3270(N6650,R4);
not not3271(N6651,R6);
not not3272(N6652,R7);
not not3273(N6666,R6);
not not3274(N6667,R7);
not not3275(N6681,R3);
not not3276(N6682,R5);
not not3277(N6695,R3);
not not3278(N6696,R4);
not not3279(N6697,R7);
not not3280(N6709,R5);
not not3281(N6710,R6);
not not3282(N6711,R7);
not not3283(N6724,R4);
not not3284(N6725,R6);
not not3285(N6737,R5);
not not3286(N6738,R6);
not not3287(N6739,R7);
not not3288(N6752,R5);
not not3289(N6753,R6);
not not3290(N6766,R4);
not not3291(N6767,R7);
not not3292(N6780,R5);
not not3293(N6781,R7);
not not3294(N6794,R6);
not not3295(N6795,R7);
not not3296(N6809,R6);
not not3297(N6822,R5);
not not3298(N6823,R7);
not not3299(N6836,R4);
not not3300(N6837,R7);
not not3301(N6850,R5);
not not3302(N6851,R6);
not not3303(N6864,R5);
not not3304(N6865,R6);
not not3305(N6876,R3);
not not3306(N6877,R5);
not not3307(N6878,R6);
not not3308(N6879,R7);
not not3309(N6891,R4);
not not3310(N6892,R6);
not not3311(N6893,R7);
not not3312(N6905,R5);
not not3313(N6906,R6);
not not3314(N6907,R7);
not not3315(N6919,R3);
not not3316(N6920,R5);
not not3317(N6921,R6);
not not3318(N6934,R5);
not not3319(N6935,R7);
not not3320(N6948,R5);
not not3321(N6949,R7);
not not3322(N6961,R5);
not not3323(N6962,R6);
not not3324(N6963,R7);
not not3325(N6976,R6);
not not3326(N6977,R7);
not not3327(N6990,R4);
not not3328(N6991,R7);
not not3329(N7004,R5);
not not3330(N7005,R7);
not not3331(N7018,R3);
not not3332(N7019,R5);
not not3333(N7032,R4);
not not3334(N7033,R5);
not not3335(N7045,R3);
not not3336(N7046,R4);
not not3337(N7047,R5);
not not3338(N7059,R4);
not not3339(N7060,R5);
not not3340(N7061,R6);
not not3341(N7073,R4);
not not3342(N7074,R6);
not not3343(N7075,R7);
not not3344(N7087,R3);
not not3345(N7088,R6);
not not3346(N7089,R7);
not not3347(N7102,R3);
not not3348(N7103,R6);
not not3349(N7116,R5);
not not3350(N7117,R6);
not not3351(N7128,R5);
not not3352(N7129,R6);
not not3353(N7130,R7);
not not3354(N7141,R5);
not not3355(N7142,R6);
not not3356(N7143,R7);
not not3357(N7153,R4);
not not3358(N7154,R5);
not not3359(N7155,R6);
not not3360(N7156,R7);
not not3361(N7167,R5);
not not3362(N7168,R6);
not not3363(N7169,R7);
not not3364(N7180,R5);
not not3365(N7181,R6);
not not3366(N7182,R7);
not not3367(N7193,R5);
not not3368(N7194,R6);
not not3369(N7195,R7);
not not3370(N7207,R4);
not not3371(N7208,R6);
not not3372(N7220,R4);
not not3373(N7221,R5);
not not3374(N7234,R5);
not not3375(N7247,R6);
not not3376(N7260,R7);
not not3377(N7273,R7);
not not3378(N7286,R7);
not not3379(N7299,R6);
not not3380(N7311,R6);
not not3381(N7312,R7);
not not3382(N7338,R5);
not not3383(N7351,R5);
not not3384(N7364,R5);
not not3385(N7377,R5);
not not3386(N7390,R4);
not not3387(N7403,R7);
not not3388(N7416,R7);
not not3389(N7429,R5);
not not3390(N7442,R5);
not not3391(N7455,R5);
not not3392(N7467,R4);
not not3393(N7468,R5);
not not3394(N7494,R7);
not not3395(N7507,R6);
not not3396(N7520,R6);
not not3397(N7531,R3);
not not3398(N7532,R4);
not not3399(N7533,R6);
not not3400(N7545,R5);
not not3401(N7546,R7);
not not3402(N7558,R6);
not not3403(N7559,R7);
not not3404(N7571,R4);
not not3405(N7572,R5);
not not3406(N7583,R4);
not not3407(N7584,R6);
not not3408(N7585,R7);
not not3409(N7597,R6);
not not3410(N7598,R7);
not not3411(N7610,R5);
not not3412(N7611,R6);
not not3413(N7621,R5);
not not3414(N7622,R6);
not not3415(N7623,R7);
not not3416(N7635,R6);
not not3417(N7647,R6);
not not3418(N7658,R4);
not not3419(N7659,R7);
not not3420(N7671,R7);
not not3421(N7683,R5);
not not3422(N7694,R4);
not not3423(N7695,R7);
not not3424(N7707,R6);
not not3425(N7731,R4);
not not3426(N7743,R4);
not not3427(N7755,R4);
not not3428(N7767,R4);
not not3429(N7779,R5);
not not3430(N7790,R4);
not not3431(N7791,R5);
not not3432(N7803,R7);
not not3433(N7814,R5);
not not3434(N7815,R7);
not not3435(N7851,R7);
not not3436(N7863,R3);
not not3437(N7874,R6);
not not3438(N7875,R7);
not not3439(N7886,R6);
not not3440(N7887,R7);
not not3441(N7899,R6);
not not3442(N7931,R4);
not not3443(N7932,R6);
not not3444(N7943,R4);
not not3445(N7954,R7);
not not3446(N7964,R4);
not not3447(N7965,R7);
not not3448(N7976,R4);
not not3449(N7987,R7);
not not3450(N7998,R7);
not not3451(N8009,R4);
not not3452(N8031,R5);
not not3453(N8061,R6);
not not3454(N8081,R4);
not not3455(N8111,R5);
not not3456(N8136,R6);
not not3457(N8151,R5);
not not3458(N8152,R6);
not not3459(N8166,R6);
not not3460(N8167,R7);
not not3461(N8182,R7);
not not3462(N8196,R6);
not not3463(N8197,R7);
not not3464(N8211,R5);
not not3465(N8212,R7);
not not3466(N8227,R7);
not not3467(N8242,R5);
not not3468(N8256,R6);
not not3469(N8257,R7);
not not3470(N8271,R5);
not not3471(N8272,R6);
not not3472(N8286,R6);
not not3473(N8287,R7);
not not3474(N8302,R6);
not not3475(N8316,R5);
not not3476(N8317,R6);
not not3477(N8331,R6);
not not3478(N8332,R7);
not not3479(N8346,R5);
not not3480(N8347,R7);
not not3481(N8362,R6);
not not3482(N8375,R6);
not not3483(N8376,R7);
not not3484(N8390,R6);
not not3485(N8404,R6);
not not3486(N8418,R6);
not not3487(N8431,R6);
not not3488(N8432,R7);
not not3489(N8445,R6);
not not3490(N8446,R7);
not not3491(N8460,R7);
not not3492(N8474,R7);
not not3493(N8487,R6);
not not3494(N8488,R7);
not not3495(N8502,R5);
not not3496(N8515,R6);
not not3497(N8516,R7);
not not3498(N8529,R6);
not not3499(N8530,R7);
not not3500(N8544,R7);
not not3501(N8558,R7);
not not3502(N8572,R7);
not not3503(N8586,R7);
not not3504(N8599,R5);
not not3505(N8600,R6);
not not3506(N8613,R6);
not not3507(N8614,R7);
not not3508(N8627,R6);
not not3509(N8628,R7);
not not3510(N8641,R6);
not not3511(N8642,R7);
not not3512(N8656,R7);
not not3513(N8670,R7);
not not3514(N8684,R6);
not not3515(N8697,R6);
not not3516(N8698,R7);
not not3517(N8711,R5);
not not3518(N8712,R7);
not not3519(N8726,R6);
not not3520(N8739,R6);
not not3521(N8740,R7);
not not3522(N8754,R6);
not not3523(N8768,R6);
not not3524(N8782,R6);
not not3525(N8796,R7);
not not3526(N8809,R6);
not not3527(N8810,R7);
not not3528(N8824,R6);
not not3529(N8837,R6);
not not3530(N8838,R7);
not not3531(N8851,R6);
not not3532(N8852,R7);
not not3533(N8865,R6);
not not3534(N8866,R7);
not not3535(N8879,R6);
not not3536(N8880,R7);
not not3537(N8894,R7);
not not3538(N8906,R6);
not not3539(N8907,R7);
not not3540(N8932,R6);
not not3541(N8933,R7);
not not3542(N8946,R6);
not not3543(N8958,R6);
not not3544(N8959,R7);
not not3545(N8971,R6);
not not3546(N8972,R7);
not not3547(N8984,R6);
not not3548(N8985,R7);
not not3549(N8998,R6);
not not3550(N9023,R6);
not not3551(N9024,R7);
not not3552(N9037,R7);
not not3553(N9050,R7);
not not3554(N9063,R7);
not not3555(N9076,R7);
not not3556(N9102,R6);
not not3557(N9115,R6);
not not3558(N9128,R7);
not not3559(N9141,R7);
not not3560(N9154,R7);
not not3561(N9167,R7);
not not3562(N9180,R7);
not not3563(N9192,R6);
not not3564(N9193,R7);
not not3565(N9205,R6);
not not3566(N9206,R7);
not not3567(N9218,R6);
not not3568(N9219,R7);
not not3569(N9232,R6);
not not3570(N9245,R7);
not not3571(N9257,R6);
not not3572(N9258,R7);
not not3573(N9270,R6);
not not3574(N9271,R7);
not not3575(N9284,R6);
not not3576(N9297,R7);
not not3577(N9310,R6);
not not3578(N9323,R6);
not not3579(N9349,R6);
not not3580(N9361,R5);
not not3581(N9362,R7);
not not3582(N9374,R5);
not not3583(N9375,R6);
not not3584(N9387,R5);
not not3585(N9388,R6);
not not3586(N9401,R6);
not not3587(N9414,R6);
not not3588(N9427,R6);
not not3589(N9439,R6);
not not3590(N9440,R7);
not not3591(N9453,R6);
not not3592(N9466,R5);
not not3593(N9479,R7);
not not3594(N9491,R6);
not not3595(N9492,R7);
not not3596(N9505,R6);
not not3597(N9517,R6);
not not3598(N9518,R7);
not not3599(N9530,R6);
not not3600(N9531,R7);
not not3601(N9544,R5);
not not3602(N9556,R6);
not not3603(N9557,R7);
not not3604(N9570,R5);
not not3605(N9582,R6);
not not3606(N9583,R7);
not not3607(N9595,R5);
not not3608(N9596,R7);
not not3609(N9609,R5);
not not3610(N9622,R7);
not not3611(N9635,R6);
not not3612(N9647,R7);
not not3613(N9659,R7);
not not3614(N9671,R7);
not not3615(N9683,R7);
not not3616(N9695,R6);
not not3617(N9707,R7);
not not3618(N9719,R7);
not not3619(N9731,R6);
not not3620(N9743,R6);
not not3621(N9767,R6);
not not3622(N9779,R6);
not not3623(N9803,R7);
not not3624(N9815,R7);
not not3625(N9826,R6);
not not3626(N9827,R7);
not not3627(N9851,R7);
not not3628(N9862,R5);
not not3629(N9863,R6);
not not3630(N9875,R6);
not not3631(N9887,R7);
not not3632(N9923,R6);
not not3633(N9935,R6);
not not3634(N9947,R6);
not not3635(N9959,R6);
not not3636(N9971,R7);
not not3637(N9983,R6);
not not3638(N9995,R6);
not not3639(N10007,R6);
not not3640(N10031,R7);
not not3641(N10043,R6);
not not3642(N10055,R6);
not not3643(N10067,R6);
not not3644(N10079,R5);
not not3645(N10091,R6);
not not3646(N10103,R7);
not not3647(N10115,R5);
not not3648(N10151,R7);
not not3649(N10163,R7);
not not3650(N10175,R6);
not not3651(N10186,R6);
not not3652(N10187,R7);
not not3653(N10199,R6);
not not3654(N10209,R5);
not not3655(N10210,R7);
not not3656(N10221,R6);
not not3657(N10231,R6);
not not3658(N10232,R7);
not not3659(N10254,R6);
not not3660(N10265,R6);
not not3661(N10287,R5);
not not3662(N10298,R6);
not not3663(N10308,R6);
not not3664(N10309,R7);
not not3665(N10320,R7);
not not3666(N10331,R6);
not not3667(N10342,R5);
not not3668(N10353,R7);
not not3669(N10364,R6);
not not3670(N10375,R5);
not not3671(N10386,R6);
not not3672(N10397,R6);
not not3673(N10408,R5);
not not3674(N10452,R6);
not not3675(N10463,R6);
not not3676(N10474,R6);
not not3677(N10485,R7);
not not3678(N10496,R7);
not not3679(N10506,R6);
not not3680(N10507,R7);
not not3681(N10518,R7);
not not3682(N10528,R6);
not not3683(N10529,R7);
not not3684(N10540,R7);
not not3685(N10550,R6);
not not3686(N10551,R7);
not not3687(N10562,R6);
not not3688(N10573,R7);
not not3689(N10584,R6);
not not3690(N10595,R7);
not not3691(N10606,R7);
not not3692(N10639,R6);
not not3693(N10650,R6);
not not3694(N10661,R4);
not not3695(N10672,R7);
not not3696(N10682,R6);
not not3697(N10702,R6);
not not3698(N10732,R5);
not not3699(N10742,R7);
not not3700(N10772,R7);
not not3701(N10782,R7);
not not3702(N10822,R6);
not not3703(N10882,R5);
not not3704(N10892,R7);
not not3705(N10902,R6);
not not3706(N10921,R6);
not not3707(N10922,R7);
not not3708(N11891,in1);
not not3709(N11892,R0);
not not3710(N11893,R1);
not not3711(N11894,R2);
not not3712(N11895,R3);
not not3713(N11909,in1);
not not3714(N11910,in2);
not not3715(N11911,R0);
not not3716(N11912,R1);
not not3717(N11913,R2);
not not3718(N11914,R3);
not not3719(N11927,in1);
not not3720(N11928,in2);
not not3721(N11929,R0);
not not3722(N11930,R1);
not not3723(N11931,R2);
not not3724(N11944,in0);
not not3725(N11945,in1);
not not3726(N11946,in2);
not not3727(N11947,R1);
not not3728(N11948,R3);
not not3729(N11961,in0);
not not3730(N11962,in2);
not not3731(N11963,R0);
not not3732(N11964,R1);
not not3733(N11965,R2);
not not3734(N11978,in0);
not not3735(N11979,in1);
not not3736(N11980,in2);
not not3737(N11981,R0);
not not3738(N11982,R2);
not not3739(N11995,R0);
not not3740(N11996,R2);
not not3741(N11997,R3);
not not3742(N12011,in0);
not not3743(N12012,R0);
not not3744(N12013,R1);
not not3745(N12014,R2);
not not3746(N12015,R3);
not not3747(N12027,in0);
not not3748(N12028,in2);
not not3749(N12029,R0);
not not3750(N12030,R2);
not not3751(N12043,in0);
not not3752(N12044,in1);
not not3753(N12045,in2);
not not3754(N12046,R1);
not not3755(N12047,R2);
not not3756(N12059,in0);
not not3757(N12060,in1);
not not3758(N12061,in2);
not not3759(N12062,R0);
not not3760(N12063,R1);
not not3761(N12075,in0);
not not3762(N12076,in1);
not not3763(N12077,in2);
not not3764(N12078,R0);
not not3765(N12079,R2);
not not3766(N12091,in0);
not not3767(N12092,in2);
not not3768(N12093,R1);
not not3769(N12094,R2);
not not3770(N12095,R3);
not not3771(N12107,in0);
not not3772(N12108,in1);
not not3773(N12109,R0);
not not3774(N12110,R2);
not not3775(N12123,in0);
not not3776(N12124,in1);
not not3777(N12125,in2);
not not3778(N12126,R0);
not not3779(N12127,R2);
not not3780(N12139,in0);
not not3781(N12140,in1);
not not3782(N12141,R1);
not not3783(N12142,R2);
not not3784(N12155,in0);
not not3785(N12156,in1);
not not3786(N12157,in2);
not not3787(N12158,R3);
not not3788(N12171,in0);
not not3789(N12172,in1);
not not3790(N12173,R1);
not not3791(N12174,R2);
not not3792(N12187,in0);
not not3793(N12188,in2);
not not3794(N12189,R0);
not not3795(N12190,R1);
not not3796(N12203,in1);
not not3797(N12204,in2);
not not3798(N12205,R0);
not not3799(N12218,in0);
not not3800(N12219,in1);
not not3801(N12220,R0);
not not3802(N12233,in1);
not not3803(N12234,in2);
not not3804(N12235,R2);
not not3805(N12248,R0);
not not3806(N12249,R1);
not not3807(N12250,R2);
not not3808(N12263,in0);
not not3809(N12264,in2);
not not3810(N12265,R0);
not not3811(N12266,R2);
not not3812(N12278,in2);
not not3813(N12279,R1);
not not3814(N12280,R3);
not not3815(N12293,in0);
not not3816(N12294,in1);
not not3817(N12295,R1);
not not3818(N12308,in1);
not not3819(N12309,R0);
not not3820(N12310,R1);
not not3821(N12311,R2);
not not3822(N12323,in0);
not not3823(N12324,R0);
not not3824(N12325,R1);
not not3825(N12326,R2);
not not3826(N12338,in2);
not not3827(N12339,R0);
not not3828(N12340,R1);
not not3829(N12341,R2);
not not3830(N12353,in0);
not not3831(N12354,in1);
not not3832(N12355,R2);
not not3833(N12368,R0);
not not3834(N12369,R1);
not not3835(N12370,R3);
not not3836(N12383,R0);
not not3837(N12384,R1);
not not3838(N12398,in2);
not not3839(N12399,R1);
not not3840(N12400,R2);
not not3841(N12413,in1);
not not3842(N12414,R0);
not not3843(N12415,R1);
not not3844(N12428,in2);
not not3845(N12429,R0);
not not3846(N12430,R1);
not not3847(N12443,in0);
not not3848(N12444,R0);
not not3849(N12445,R1);
not not3850(N12458,in1);
not not3851(N12459,in2);
not not3852(N12460,R0);
not not3853(N12461,R1);
not not3854(N12473,in0);
not not3855(N12474,in1);
not not3856(N12475,in2);
not not3857(N12476,R0);
not not3858(N12488,in0);
not not3859(N12489,in1);
not not3860(N12490,in2);
not not3861(N12491,R1);
not not3862(N12503,in2);
not not3863(N12504,R0);
not not3864(N12505,R1);
not not3865(N12506,R2);
not not3866(N12518,in1);
not not3867(N12519,in2);
not not3868(N12520,R0);
not not3869(N12521,R1);
not not3870(N12533,in0);
not not3871(N12534,in1);
not not3872(N12535,R0);
not not3873(N12536,R2);
not not3874(N12548,in0);
not not3875(N12549,R1);
not not3876(N12550,R2);
not not3877(N12551,R3);
not not3878(N12563,in1);
not not3879(N12564,in2);
not not3880(N12565,R1);
not not3881(N12566,R2);
not not3882(N12578,in0);
not not3883(N12579,in2);
not not3884(N12580,R1);
not not3885(N12593,in1);
not not3886(N12594,R0);
not not3887(N12595,R1);
not not3888(N12596,R2);
not not3889(N12608,in0);
not not3890(N12609,R1);
not not3891(N12610,R2);
not not3892(N12611,R3);
not not3893(N12623,in2);
not not3894(N12624,R1);
not not3895(N12625,R2);
not not3896(N12626,R3);
not not3897(N12638,in0);
not not3898(N12639,in1);
not not3899(N12640,in2);
not not3900(N12641,R3);
not not3901(N12653,in1);
not not3902(N12654,R1);
not not3903(N12655,R2);
not not3904(N12668,in0);
not not3905(N12669,in1);
not not3906(N12670,R2);
not not3907(N12683,in0);
not not3908(N12684,in1);
not not3909(N12685,R0);
not not3910(N12686,R2);
not not3911(N12698,in2);
not not3912(N12699,R1);
not not3913(N12700,R2);
not not3914(N12713,in2);
not not3915(N12714,R0);
not not3916(N12715,R2);
not not3917(N12728,in0);
not not3918(N12729,in1);
not not3919(N12730,R3);
not not3920(N12743,in2);
not not3921(N12744,R0);
not not3922(N12745,R3);
not not3923(N12758,in2);
not not3924(N12759,R1);
not not3925(N12760,R2);
not not3926(N12772,in0);
not not3927(N12773,R1);
not not3928(N12774,R3);
not not3929(N12786,in2);
not not3930(N12787,R1);
not not3931(N12788,R3);
not not3932(N12800,in1);
not not3933(N12801,R1);
not not3934(N12802,R2);
not not3935(N12814,R1);
not not3936(N12815,R2);
not not3937(N12828,in0);
not not3938(N12829,R0);
not not3939(N12830,R2);
not not3940(N12842,in0);
not not3941(N12843,in1);
not not3942(N12844,R2);
not not3943(N12856,in0);
not not3944(N12857,in1);
not not3945(N12858,in2);
not not3946(N12859,R1);
not not3947(N12870,in0);
not not3948(N12871,in2);
not not3949(N12872,R2);
not not3950(N12884,in0);
not not3951(N12885,in1);
not not3952(N12886,R2);
not not3953(N12898,in1);
not not3954(N12899,R0);
not not3955(N12900,R1);
not not3956(N12912,R1);
not not3957(N12913,R2);
not not3958(N12926,in0);
not not3959(N12927,R1);
not not3960(N12928,R2);
not not3961(N12940,in2);
not not3962(N12941,R0);
not not3963(N12942,R1);
not not3964(N12943,R3);
not not3965(N12954,in0);
not not3966(N12955,R0);
not not3967(N12956,R1);
not not3968(N12957,R3);
not not3969(N12968,R1);
not not3970(N12969,R2);
not not3971(N12970,R3);
not not3972(N12982,in0);
not not3973(N12983,R1);
not not3974(N12984,R2);
not not3975(N12996,R0);
not not3976(N12997,R1);
not not3977(N12998,R2);
not not3978(N13010,in2);
not not3979(N13011,R0);
not not3980(N13012,R1);
not not3981(N13013,R2);
not not3982(N13024,in1);
not not3983(N13025,R0);
not not3984(N13038,in0);
not not3985(N13039,R1);
not not3986(N13052,in0);
not not3987(N13053,in2);
not not3988(N13054,R0);
not not3989(N13066,in0);
not not3990(N13067,R2);
not not3991(N13068,R3);
not not3992(N13080,in1);
not not3993(N13081,in2);
not not3994(N13082,R0);
not not3995(N13083,R3);
not not3996(N13094,in0);
not not3997(N13095,in1);
not not3998(N13096,R0);
not not3999(N13097,R1);
not not4000(N13108,R0);
not not4001(N13109,R2);
not not4002(N13110,R3);
not not4003(N13122,in0);
not not4004(N13123,R0);
not not4005(N13124,R2);
not not4006(N13136,R0);
not not4007(N13137,R3);
not not4008(N13150,in1);
not not4009(N13151,in2);
not not4010(N13152,R1);
not not4011(N13164,in0);
not not4012(N13165,in1);
not not4013(N13166,R1);
not not4014(N13178,in0);
not not4015(N13179,in1);
not not4016(N13180,R0);
not not4017(N13181,R3);
not not4018(N13192,in0);
not not4019(N13193,R2);
not not4020(N13206,in2);
not not4021(N13207,R0);
not not4022(N13208,R3);
not not4023(N13220,in1);
not not4024(N13221,in2);
not not4025(N13222,R1);
not not4026(N13234,in1);
not not4027(N13235,in2);
not not4028(N13236,R0);
not not4029(N13237,R1);
not not4030(N13248,in0);
not not4031(N13249,in2);
not not4032(N13250,R0);
not not4033(N13251,R1);
not not4034(N13262,in0);
not not4035(N13263,in1);
not not4036(N13264,R1);
not not4037(N13265,R2);
not not4038(N13276,in0);
not not4039(N13277,in2);
not not4040(N13278,R2);
not not4041(N13290,in2);
not not4042(N13291,R1);
not not4043(N13292,R3);
not not4044(N13304,in0);
not not4045(N13305,in2);
not not4046(N13306,R1);
not not4047(N13318,in2);
not not4048(N13319,R0);
not not4049(N13320,R1);
not not4050(N13332,R0);
not not4051(N13345,R2);
not not4052(N13358,R1);
not not4053(N13359,R2);
not not4054(N13371,R1);
not not4055(N13384,in2);
not not4056(N13385,R1);
not not4057(N13397,in0);
not not4058(N13398,R0);
not not4059(N13410,R1);
not not4060(N13423,R0);
not not4061(N13424,R1);
not not4062(N13449,in2);
not not4063(N13450,R1);
not not4064(N13451,R2);
not not4065(N13462,R0);
not not4066(N13463,R1);
not not4067(N13475,in2);
not not4068(N13476,R0);
not not4069(N13488,R2);
not not4070(N13489,R3);
not not4071(N13501,in2);
not not4072(N13502,R0);
not not4073(N13514,R0);
not not4074(N13515,R3);
not not4075(N13527,in2);
not not4076(N13528,R0);
not not4077(N13540,R0);
not not4078(N13541,R2);
not not4079(N13542,R3);
not not4080(N13553,in2);
not not4081(N13554,R0);
not not4082(N13555,R1);
not not4083(N13566,in0);
not not4084(N13567,R1);
not not4085(N13579,in0);
not not4086(N13580,in2);
not not4087(N13581,R2);
not not4088(N13592,in1);
not not4089(N13593,in2);
not not4090(N13605,R1);
not not4091(N13606,R2);
not not4092(N13618,in1);
not not4093(N13619,R3);
not not4094(N13631,in0);
not not4095(N13644,in1);
not not4096(N13645,R2);
not not4097(N13646,R3);
not not4098(N13657,R1);
not not4099(N13658,R2);
not not4100(N13670,in1);
not not4101(N13671,in2);
not not4102(N13683,in1);
not not4103(N13684,R1);
not not4104(N13696,in0);
not not4105(N13697,in2);
not not4106(N13709,in2);
not not4107(N13710,R0);
not not4108(N13711,R1);
not not4109(N13722,in1);
not not4110(N13723,in2);
not not4111(N13724,R0);
not not4112(N13735,in0);
not not4113(N13736,in1);
not not4114(N13737,R0);
not not4115(N13738,R2);
not not4116(N13748,in2);
not not4117(N13761,in0);
not not4118(N13762,R1);
not not4119(N13774,R0);
not not4120(N13787,in1);
not not4121(N13788,R1);
not not4122(N13800,in2);
not not4123(N13813,in0);
not not4124(N13814,R3);
not not4125(N13826,R0);
not not4126(N13827,R1);
not not4127(N13839,in2);
not not4128(N13840,R1);
not not4129(N13852,in0);
not not4130(N13853,R1);
not not4131(N13865,in0);
not not4132(N13866,in2);
not not4133(N13878,in0);
not not4134(N13879,R2);
not not4135(N13891,in1);
not not4136(N13892,R1);
not not4137(N13904,R0);
not not4138(N13905,R1);
not not4139(N13917,in0);
not not4140(N13918,R1);
not not4141(N13930,in2);
not not4142(N13931,R0);
not not4143(N13942,R0);
not not4144(N13954,R0);
not not4145(N13966,R3);
not not4146(N13990,in1);
not not4147(N13991,R3);
not not4148(N14002,R1);
not not4149(N14003,R2);
not not4150(N14014,in0);
not not4151(N14026,in2);
not not4152(N14038,in1);
not not4153(N14039,in2);
not not4154(N14050,in2);
not not4155(N14051,R0);
not not4156(N14052,R1);
not not4157(N14062,in1);
not not4158(N14063,in2);
not not4159(N14074,in1);
not not4160(N14075,in2);
not not4161(N14076,R3);
not not4162(N14086,in1);
not not4163(N14098,in0);
not not4164(N14099,R0);
not not4165(N14110,in2);
not not4166(N14111,R0);
not not4167(N14122,in1);
not not4168(N14134,R2);
not not4169(N14146,in1);
not not4170(N14147,R3);
not not4171(N14158,in2);
not not4172(N14159,R3);
not not4173(N14170,R1);
not not4174(N14171,R3);
not not4175(N14182,in2);
not not4176(N14183,R1);
not not4177(N14194,in2);
not not4178(N14195,R1);
not not4179(N14206,in2);
not not4180(N14207,R0);
not not4181(N14208,R2);
not not4182(N14218,in2);
not not4183(N14219,R0);
not not4184(N14230,R2);
not not4185(N14242,in0);
not not4186(N14243,R0);
not not4187(N14254,in0);
not not4188(N14255,in1);
not not4189(N14277,R0);
not not4190(N14299,R1);
not not4191(N14321,R0);
not not4192(N14322,R1);
not not4193(N14332,R1);
not not4194(N14365,in1);
not not4195(N14376,R2);
not not4196(N14387,R1);
not not4197(N14398,in0);
not not4198(N14409,in2);
not not4199(N14410,R1);
not not4200(N14431,R1);
not not4201(N14452,in1);
not not4202(N14462,R3);
not not4203(N14482,in0);
not not4204(N14510,in2);
not not4205(N14511,R0);
not not4206(N14512,R2);
not not4207(N14513,R3);
not not4208(N14514,R4);
not not4209(N14515,R5);
not not4210(N14526,in2);
not not4211(N14527,R0);
not not4212(N14528,R2);
not not4213(N14529,R3);
not not4214(N14530,R4);
not not4215(N14531,R5);
not not4216(N14542,in0);
not not4217(N14543,in1);
not not4218(N14544,in2);
not not4219(N14545,R2);
not not4220(N14546,R4);
not not4221(N14547,R5);
not not4222(N14558,in1);
not not4223(N14559,R0);
not not4224(N14560,R1);
not not4225(N14561,R2);
not not4226(N14562,R3);
not not4227(N14563,R5);
not not4228(N14573,in1);
not not4229(N14574,R0);
not not4230(N14575,R1);
not not4231(N14576,R2);
not not4232(N14577,R4);
not not4233(N14578,R5);
not not4234(N14588,in1);
not not4235(N14589,in2);
not not4236(N14590,R0);
not not4237(N14591,R2);
not not4238(N14592,R4);
not not4239(N14593,R5);
not not4240(N14603,in0);
not not4241(N14604,in1);
not not4242(N14605,R2);
not not4243(N14606,R3);
not not4244(N14607,R5);
not not4245(N14618,in0);
not not4246(N14619,in1);
not not4247(N14620,R0);
not not4248(N14621,R1);
not not4249(N14622,R3);
not not4250(N14623,R5);
not not4251(N14633,in0);
not not4252(N14634,in2);
not not4253(N14635,R0);
not not4254(N14636,R2);
not not4255(N14637,R3);
not not4256(N14648,in1);
not not4257(N14649,in2);
not not4258(N14650,R1);
not not4259(N14651,R2);
not not4260(N14652,R4);
not not4261(N14663,in1);
not not4262(N14664,in2);
not not4263(N14665,R1);
not not4264(N14666,R2);
not not4265(N14667,R3);
not not4266(N14678,in1);
not not4267(N14679,in2);
not not4268(N14680,R0);
not not4269(N14681,R2);
not not4270(N14682,R5);
not not4271(N14693,in0);
not not4272(N14694,in1);
not not4273(N14695,in2);
not not4274(N14696,R0);
not not4275(N14697,R3);
not not4276(N14708,in1);
not not4277(N14709,R1);
not not4278(N14710,R2);
not not4279(N14711,R3);
not not4280(N14722,in2);
not not4281(N14723,R1);
not not4282(N14724,R2);
not not4283(N14725,R3);
not not4284(N14726,R5);
not not4285(N14736,in0);
not not4286(N14737,in1);
not not4287(N14738,in2);
not not4288(N14739,R1);
not not4289(N14740,R2);
not not4290(N14750,in1);
not not4291(N14751,R1);
not not4292(N14752,R3);
not not4293(N14753,R4);
not not4294(N14754,R5);
not not4295(N14764,in1);
not not4296(N14765,R1);
not not4297(N14766,R3);
not not4298(N14767,R4);
not not4299(N14768,R5);
not not4300(N14778,in0);
not not4301(N14779,in2);
not not4302(N14780,R4);
not not4303(N14781,R5);
not not4304(N14792,in1);
not not4305(N14793,in2);
not not4306(N14794,R1);
not not4307(N14795,R2);
not not4308(N14796,R4);
not not4309(N14806,R0);
not not4310(N14807,R1);
not not4311(N14808,R2);
not not4312(N14809,R3);
not not4313(N14820,R0);
not not4314(N14821,R1);
not not4315(N14822,R2);
not not4316(N14823,R4);
not not4317(N14824,R5);
not not4318(N14834,in0);
not not4319(N14835,in2);
not not4320(N14836,R0);
not not4321(N14837,R3);
not not4322(N14838,R4);
not not4323(N14848,in0);
not not4324(N14849,in1);
not not4325(N14850,R0);
not not4326(N14851,R3);
not not4327(N14852,R4);
not not4328(N14862,in1);
not not4329(N14863,R2);
not not4330(N14864,R4);
not not4331(N14865,R5);
not not4332(N14876,in1);
not not4333(N14877,R1);
not not4334(N14878,R3);
not not4335(N14879,R4);
not not4336(N14880,R5);
not not4337(N14890,in0);
not not4338(N14891,R2);
not not4339(N14892,R4);
not not4340(N14893,R5);
not not4341(N14904,R0);
not not4342(N14905,R1);
not not4343(N14906,R2);
not not4344(N14907,R3);
not not4345(N14908,R5);
not not4346(N14918,in1);
not not4347(N14919,R3);
not not4348(N14920,R4);
not not4349(N14921,R5);
not not4350(N14932,in0);
not not4351(N14933,R0);
not not4352(N14934,R2);
not not4353(N14935,R4);
not not4354(N14946,in0);
not not4355(N14947,in1);
not not4356(N14948,R1);
not not4357(N14949,R2);
not not4358(N14950,R4);
not not4359(N14960,in0);
not not4360(N14961,R0);
not not4361(N14962,R1);
not not4362(N14963,R5);
not not4363(N14974,in1);
not not4364(N14975,in2);
not not4365(N14976,R3);
not not4366(N14977,R5);
not not4367(N14988,in1);
not not4368(N14989,R1);
not not4369(N14990,R2);
not not4370(N14991,R4);
not not4371(N14992,R5);
not not4372(N15002,in1);
not not4373(N15003,in2);
not not4374(N15004,R0);
not not4375(N15005,R4);
not not4376(N15006,R5);
not not4377(N15016,in2);
not not4378(N15017,R0);
not not4379(N15018,R2);
not not4380(N15019,R4);
not not4381(N15030,in1);
not not4382(N15031,in2);
not not4383(N15032,R0);
not not4384(N15033,R2);
not not4385(N15034,R4);
not not4386(N15044,in0);
not not4387(N15045,in2);
not not4388(N15046,R0);
not not4389(N15047,R4);
not not4390(N15048,R5);
not not4391(N15058,in0);
not not4392(N15059,R1);
not not4393(N15060,R2);
not not4394(N15061,R4);
not not4395(N15072,in0);
not not4396(N15073,in1);
not not4397(N15074,in2);
not not4398(N15075,R1);
not not4399(N15076,R5);
not not4400(N15086,in2);
not not4401(N15087,R1);
not not4402(N15088,R4);
not not4403(N15089,R5);
not not4404(N15100,in2);
not not4405(N15101,R1);
not not4406(N15102,R3);
not not4407(N15103,R4);
not not4408(N15104,R5);
not not4409(N15114,in0);
not not4410(N15115,R0);
not not4411(N15116,R1);
not not4412(N15117,R3);
not not4413(N15118,R5);
not not4414(N15128,in1);
not not4415(N15129,in2);
not not4416(N15130,R1);
not not4417(N15131,R5);
not not4418(N15142,in0);
not not4419(N15143,in2);
not not4420(N15144,R0);
not not4421(N15145,R2);
not not4422(N15146,R3);
not not4423(N15156,in0);
not not4424(N15157,R0);
not not4425(N15158,R2);
not not4426(N15159,R3);
not not4427(N15170,in0);
not not4428(N15171,R0);
not not4429(N15172,R2);
not not4430(N15173,R5);
not not4431(N15184,R1);
not not4432(N15185,R2);
not not4433(N15186,R3);
not not4434(N15187,R4);
not not4435(N15198,in0);
not not4436(N15199,in2);
not not4437(N15200,R5);
not not4438(N15211,R0);
not not4439(N15212,R2);
not not4440(N15213,R5);
not not4441(N15224,in2);
not not4442(N15225,R1);
not not4443(N15226,R4);
not not4444(N15227,R5);
not not4445(N15237,R0);
not not4446(N15238,R1);
not not4447(N15239,R5);
not not4448(N15250,in0);
not not4449(N15251,in2);
not not4450(N15252,R0);
not not4451(N15253,R3);
not not4452(N15254,R5);
not not4453(N15263,R0);
not not4454(N15264,R4);
not not4455(N15265,R5);
not not4456(N15276,in2);
not not4457(N15277,R0);
not not4458(N15278,R5);
not not4459(N15289,in0);
not not4460(N15290,in1);
not not4461(N15291,R0);
not not4462(N15302,in0);
not not4463(N15303,R1);
not not4464(N15304,R2);
not not4465(N15305,R4);
not not4466(N15315,R0);
not not4467(N15316,R1);
not not4468(N15317,R4);
not not4469(N15318,R5);
not not4470(N15328,in0);
not not4471(N15329,in2);
not not4472(N15330,R5);
not not4473(N15341,R0);
not not4474(N15342,R2);
not not4475(N15343,R4);
not not4476(N15344,R5);
not not4477(N15354,in2);
not not4478(N15355,R0);
not not4479(N15356,R2);
not not4480(N15357,R4);
not not4481(N15367,in2);
not not4482(N15368,R2);
not not4483(N15369,R5);
not not4484(N15380,in1);
not not4485(N15381,in2);
not not4486(N15382,R0);
not not4487(N15383,R3);
not not4488(N15393,in1);
not not4489(N15394,R1);
not not4490(N15395,R2);
not not4491(N15396,R4);
not not4492(N15406,in1);
not not4493(N15407,R0);
not not4494(N15408,R2);
not not4495(N15409,R5);
not not4496(N15419,in2);
not not4497(N15420,R3);
not not4498(N15421,R5);
not not4499(N15432,in1);
not not4500(N15433,R3);
not not4501(N15434,R5);
not not4502(N15445,in0);
not not4503(N15446,R2);
not not4504(N15447,R3);
not not4505(N15448,R4);
not not4506(N15458,in2);
not not4507(N15459,R0);
not not4508(N15460,R2);
not not4509(N15461,R4);
not not4510(N15471,in2);
not not4511(N15472,R1);
not not4512(N15473,R2);
not not4513(N15474,R4);
not not4514(N15484,in0);
not not4515(N15485,in1);
not not4516(N15486,R4);
not not4517(N15497,R2);
not not4518(N15498,R3);
not not4519(N15499,R5);
not not4520(N15510,in2);
not not4521(N15511,R1);
not not4522(N15512,R2);
not not4523(N15513,R4);
not not4524(N15523,in0);
not not4525(N15524,R0);
not not4526(N15525,R3);
not not4527(N15526,R5);
not not4528(N15536,in1);
not not4529(N15537,in2);
not not4530(N15538,R2);
not not4531(N15539,R3);
not not4532(N15540,R5);
not not4533(N15549,in2);
not not4534(N15550,R0);
not not4535(N15551,R2);
not not4536(N15552,R3);
not not4537(N15562,in0);
not not4538(N15563,R3);
not not4539(N15564,R5);
not not4540(N15575,in1);
not not4541(N15576,R2);
not not4542(N15577,R3);
not not4543(N15588,in2);
not not4544(N15589,R0);
not not4545(N15590,R1);
not not4546(N15591,R4);
not not4547(N15601,in0);
not not4548(N15602,R1);
not not4549(N15603,R3);
not not4550(N15604,R4);
not not4551(N15614,in1);
not not4552(N15615,R2);
not not4553(N15616,R4);
not not4554(N15617,R5);
not not4555(N15627,in0);
not not4556(N15628,in1);
not not4557(N15629,in2);
not not4558(N15630,R5);
not not4559(N15640,in1);
not not4560(N15641,in2);
not not4561(N15642,R3);
not not4562(N15653,in1);
not not4563(N15654,in2);
not not4564(N15655,R1);
not not4565(N15656,R3);
not not4566(N15666,in0);
not not4567(N15667,in1);
not not4568(N15668,R0);
not not4569(N15669,R3);
not not4570(N15670,R5);
not not4571(N15679,in0);
not not4572(N15680,in1);
not not4573(N15681,R3);
not not4574(N15682,R4);
not not4575(N15692,in2);
not not4576(N15693,R0);
not not4577(N15694,R2);
not not4578(N15705,R1);
not not4579(N15706,R2);
not not4580(N15707,R4);
not not4581(N15708,R5);
not not4582(N15718,in1);
not not4583(N15719,R1);
not not4584(N15720,R4);
not not4585(N15721,R5);
not not4586(N15731,in0);
not not4587(N15732,in1);
not not4588(N15733,R3);
not not4589(N15744,in1);
not not4590(N15745,in2);
not not4591(N15746,R4);
not not4592(N15747,R5);
not not4593(N15757,in0);
not not4594(N15758,in2);
not not4595(N15759,R4);
not not4596(N15760,R5);
not not4597(N15770,in1);
not not4598(N15771,in2);
not not4599(N15772,R3);
not not4600(N15783,in0);
not not4601(N15784,in1);
not not4602(N15785,R3);
not not4603(N15796,in0);
not not4604(N15797,in1);
not not4605(N15798,in2);
not not4606(N15799,R2);
not not4607(N15800,R5);
not not4608(N15809,in1);
not not4609(N15810,in2);
not not4610(N15811,R0);
not not4611(N15812,R1);
not not4612(N15822,in1);
not not4613(N15823,R0);
not not4614(N15824,R2);
not not4615(N15825,R4);
not not4616(N15834,R0);
not not4617(N15835,R3);
not not4618(N15846,R1);
not not4619(N15847,R3);
not not4620(N15848,R4);
not not4621(N15858,R2);
not not4622(N15859,R3);
not not4623(N15860,R5);
not not4624(N15870,in1);
not not4625(N15871,R1);
not not4626(N15872,R3);
not not4627(N15882,R0);
not not4628(N15883,R2);
not not4629(N15884,R4);
not not4630(N15894,R0);
not not4631(N15895,R2);
not not4632(N15896,R3);
not not4633(N15897,R5);
not not4634(N15906,R0);
not not4635(N15907,R2);
not not4636(N15908,R3);
not not4637(N15909,R5);
not not4638(N15918,in1);
not not4639(N15919,R3);
not not4640(N15920,R4);
not not4641(N15930,in2);
not not4642(N15931,R3);
not not4643(N15932,R4);
not not4644(N15942,in1);
not not4645(N15943,R3);
not not4646(N15944,R4);
not not4647(N15954,R4);
not not4648(N15955,R5);
not not4649(N15966,in1);
not not4650(N15967,in2);
not not4651(N15968,R4);
not not4652(N15978,in0);
not not4653(N15979,R0);
not not4654(N15980,R4);
not not4655(N15990,in2);
not not4656(N15991,R3);
not not4657(N15992,R4);
not not4658(N15993,R5);
not not4659(N16002,R1);
not not4660(N16003,R3);
not not4661(N16004,R4);
not not4662(N16005,R5);
not not4663(N16014,in1);
not not4664(N16015,R0);
not not4665(N16016,R4);
not not4666(N16026,in2);
not not4667(N16027,R0);
not not4668(N16028,R2);
not not4669(N16029,R4);
not not4670(N16038,R0);
not not4671(N16039,R3);
not not4672(N16040,R4);
not not4673(N16050,in0);
not not4674(N16051,R0);
not not4675(N16052,R4);
not not4676(N16062,in1);
not not4677(N16063,R0);
not not4678(N16064,R2);
not not4679(N16065,R4);
not not4680(N16074,R1);
not not4681(N16075,R3);
not not4682(N16086,R0);
not not4683(N16087,R4);
not not4684(N16098,in0);
not not4685(N16099,in2);
not not4686(N16100,R4);
not not4687(N16110,in0);
not not4688(N16111,in1);
not not4689(N16112,R2);
not not4690(N16122,in0);
not not4691(N16123,R0);
not not4692(N16124,R2);
not not4693(N16134,in1);
not not4694(N16135,R1);
not not4695(N16136,R3);
not not4696(N16137,R5);
not not4697(N16146,R0);
not not4698(N16147,R1);
not not4699(N16148,R3);
not not4700(N16149,R5);
not not4701(N16158,R0);
not not4702(N16159,R1);
not not4703(N16160,R3);
not not4704(N16161,R5);
not not4705(N16170,R0);
not not4706(N16171,R3);
not not4707(N16172,R4);
not not4708(N16182,in1);
not not4709(N16183,R0);
not not4710(N16184,R3);
not not4711(N16194,in0);
not not4712(N16195,in1);
not not4713(N16196,R0);
not not4714(N16206,R1);
not not4715(N16207,R3);
not not4716(N16218,in0);
not not4717(N16219,in1);
not not4718(N16220,in2);
not not4719(N16221,R2);
not not4720(N16230,in0);
not not4721(N16231,R2);
not not4722(N16242,R3);
not not4723(N16243,R4);
not not4724(N16244,R5);
not not4725(N16254,in0);
not not4726(N16255,R1);
not not4727(N16256,R3);
not not4728(N16266,in2);
not not4729(N16267,R2);
not not4730(N16278,R0);
not not4731(N16279,R1);
not not4732(N16280,R3);
not not4733(N16290,in0);
not not4734(N16291,R1);
not not4735(N16292,R4);
not not4736(N16302,in2);
not not4737(N16303,R3);
not not4738(N16304,R4);
not not4739(N16314,in2);
not not4740(N16315,R1);
not not4741(N16316,R4);
not not4742(N16317,R5);
not not4743(N16326,R2);
not not4744(N16327,R3);
not not4745(N16328,R4);
not not4746(N16338,in0);
not not4747(N16339,in2);
not not4748(N16350,R0);
not not4749(N16351,R2);
not not4750(N16352,R5);
not not4751(N16362,in2);
not not4752(N16363,R2);
not not4753(N16364,R3);
not not4754(N16365,R5);
not not4755(N16374,R2);
not not4756(N16375,R4);
not not4757(N16376,R5);
not not4758(N16386,in1);
not not4759(N16387,R1);
not not4760(N16388,R3);
not not4761(N16398,in2);
not not4762(N16399,R1);
not not4763(N16400,R3);
not not4764(N16410,in0);
not not4765(N16411,R2);
not not4766(N16422,in2);
not not4767(N16423,R4);
not not4768(N16434,in2);
not not4769(N16435,R3);
not not4770(N16446,in1);
not not4771(N16447,in2);
not not4772(N16448,R0);
not not4773(N16458,R0);
not not4774(N16459,R2);
not not4775(N16460,R5);
not not4776(N16469,in2);
not not4777(N16480,in0);
not not4778(N16491,R0);
not not4779(N16492,R2);
not not4780(N16502,in1);
not not4781(N16503,R4);
not not4782(N16513,in1);
not not4783(N16514,R0);
not not4784(N16515,R5);
not not4785(N16524,R2);
not not4786(N16525,R4);
not not4787(N16535,in2);
not not4788(N16536,R2);
not not4789(N16546,in1);
not not4790(N16547,R1);
not not4791(N16557,R1);
not not4792(N16558,R2);
not not4793(N16568,R1);
not not4794(N16569,R2);
not not4795(N16579,in1);
not not4796(N16580,R2);
not not4797(N16581,R5);
not not4798(N16590,in1);
not not4799(N16591,R1);
not not4800(N16601,in2);
not not4801(N16602,R1);
not not4802(N16612,R0);
not not4803(N16613,R3);
not not4804(N16623,in1);
not not4805(N16624,R0);
not not4806(N16634,in1);
not not4807(N16635,in2);
not not4808(N16636,R1);
not not4809(N16645,R0);
not not4810(N16646,R4);
not not4811(N16656,R1);
not not4812(N16657,R4);
not not4813(N16658,R5);
not not4814(N16667,in1);
not not4815(N16668,R0);
not not4816(N16678,in1);
not not4817(N16679,R3);
not not4818(N16689,in1);
not not4819(N16690,R0);
not not4820(N16700,R3);
not not4821(N16701,R4);
not not4822(N16702,R5);
not not4823(N16711,in1);
not not4824(N16712,R0);
not not4825(N16713,R2);
not not4826(N16722,R0);
not not4827(N16723,R2);
not not4828(N16733,in1);
not not4829(N16734,R0);
not not4830(N16735,R3);
not not4831(N16744,R2);
not not4832(N16745,R4);
not not4833(N16755,in1);
not not4834(N16756,R1);
not not4835(N16766,in0);
not not4836(N16767,R2);
not not4837(N16768,R4);
not not4838(N16777,in0);
not not4839(N16778,in2);
not not4840(N16788,R2);
not not4841(N16789,R5);
not not4842(N16799,R3);
not not4843(N16800,R4);
not not4844(N16810,R0);
not not4845(N16811,R2);
not not4846(N16812,R4);
not not4847(N16821,in2);
not not4848(N16822,R3);
not not4849(N16832,R2);
not not4850(N16833,R3);
not not4851(N16843,R1);
not not4852(N16844,R3);
not not4853(N16845,R5);
not not4854(N16854,in1);
not not4855(N16855,R1);
not not4856(N16856,R5);
not not4857(N16865,in1);
not not4858(N16876,in2);
not not4859(N16887,in1);
not not4860(N16888,R3);
not not4861(N16889,R5);
not not4862(N16898,R5);
not not4863(N16908,in1);
not not4864(N16909,R0);
not not4865(N16918,in0);
not not4866(N16919,in1);
not not4867(N16928,R4);
not not4868(N16938,in0);
not not4869(N16939,in1);
not not4870(N16948,in1);
not not4871(N16949,R0);
not not4872(N16958,in1);
not not4873(N16968,R5);
not not4874(N16978,in2);
not not4875(N16988,R3);
not not4876(N16998,R4);
not not4877(N17008,in2);
not not4878(N17009,R4);
not not4879(N17018,R3);
not not4880(N17019,R5);
not not4881(N17028,R0);
not not4882(N17029,R3);
not not4883(N17038,in2);
not not4884(N17048,in1);
not not4885(N17049,R4);
not not4886(N17058,R3);
not not4887(N17068,R2);
not not4888(N17077,R2);
not not4889(N17086,R2);
not not4890(N17095,R1);
not not4891(N17104,R1);
not not4892(N17113,in2);
not not4893(N17122,R2);
not not4894(N17131,R4);
not not4895(N17140,R0);
not not4896(N17149,in2);
not not4897(N17165,in2);
not not4898(N17166,R0);
not not4899(N17167,R1);
not not4900(N17168,R2);
not not4901(N17169,R3);
not not4902(N17170,R6);
not not4903(N17171,R7);
not not4904(N17179,in1);
not not4905(N17180,R0);
not not4906(N17181,R1);
not not4907(N17182,R3);
not not4908(N17183,R4);
not not4909(N17184,R6);
not not4910(N17185,R7);
not not4911(N17193,in1);
not not4912(N17194,R1);
not not4913(N17195,R2);
not not4914(N17196,R3);
not not4915(N17197,R4);
not not4916(N17198,R6);
not not4917(N17199,R7);
not not4918(N17207,in2);
not not4919(N17208,R1);
not not4920(N17209,R2);
not not4921(N17210,R3);
not not4922(N17211,R4);
not not4923(N17212,R6);
not not4924(N17213,R7);
not not4925(N17221,in1);
not not4926(N17222,R0);
not not4927(N17223,R1);
not not4928(N17224,R5);
not not4929(N17225,R6);
not not4930(N17226,R7);
not not4931(N17234,in1);
not not4932(N17235,R0);
not not4933(N17236,R4);
not not4934(N17237,R5);
not not4935(N17238,R6);
not not4936(N17239,R7);
not not4937(N17247,in1);
not not4938(N17248,R1);
not not4939(N17249,R4);
not not4940(N17250,R5);
not not4941(N17251,R6);
not not4942(N17252,R7);
not not4943(N17260,R0);
not not4944(N17261,R2);
not not4945(N17262,R4);
not not4946(N17263,R5);
not not4947(N17264,R6);
not not4948(N17265,R7);
not not4949(N17273,R0);
not not4950(N17274,R1);
not not4951(N17275,R3);
not not4952(N17276,R4);
not not4953(N17277,R6);
not not4954(N17278,R7);
not not4955(N17286,R2);
not not4956(N17287,R3);
not not4957(N17288,R4);
not not4958(N17289,R5);
not not4959(N17290,R6);
not not4960(N17298,in1);
not not4961(N17299,R0);
not not4962(N17300,R3);
not not4963(N17301,R4);
not not4964(N17302,R6);
not not4965(N17310,R0);
not not4966(N17311,R1);
not not4967(N17312,R3);
not not4968(N17313,R5);
not not4969(N17314,R7);
not not4970(N17322,in1);
not not4971(N17323,R0);
not not4972(N17324,R2);
not not4973(N17325,R6);
not not4974(N17326,R7);
not not4975(N17334,in1);
not not4976(N17335,R0);
not not4977(N17336,R5);
not not4978(N17337,R6);
not not4979(N17338,R7);
not not4980(N17346,in0);
not not4981(N17347,in1);
not not4982(N17348,R2);
not not4983(N17349,R3);
not not4984(N17350,R6);
not not4985(N17358,R0);
not not4986(N17359,R2);
not not4987(N17360,R4);
not not4988(N17361,R5);
not not4989(N17362,R6);
not not4990(N17370,in2);
not not4991(N17371,R2);
not not4992(N17372,R4);
not not4993(N17373,R5);
not not4994(N17374,R7);
not not4995(N17382,in2);
not not4996(N17383,R0);
not not4997(N17384,R2);
not not4998(N17385,R6);
not not4999(N17386,R7);
not not5000(N17394,in1);
not not5001(N17395,R5);
not not5002(N17396,R6);
not not5003(N17397,R7);
not not5004(N17405,R0);
not not5005(N17406,R3);
not not5006(N17407,R6);
not not5007(N17408,R7);
not not5008(N17416,R2);
not not5009(N17417,R3);
not not5010(N17418,R4);
not not5011(N17419,R7);
not not5012(N17427,in1);
not not5013(N17428,R0);
not not5014(N17429,R3);
not not5015(N17430,R7);
not not5016(N17438,in1);
not not5017(N17439,R1);
not not5018(N17440,R4);
not not5019(N17441,R5);
not not5020(N17449,R1);
not not5021(N17450,R2);
not not5022(N17451,R4);
not not5023(N17452,R7);
not not5024(N17460,in1);
not not5025(N17461,R0);
not not5026(N17462,R1);
not not5027(N17463,R5);
not not5028(N17471,in1);
not not5029(N17472,R0);
not not5030(N17473,R5);
not not5031(N17474,R6);
not not5032(N17482,in2);
not not5033(N17483,R0);
not not5034(N17484,R4);
not not5035(N17485,R5);
not not5036(N17493,in2);
not not5037(N17494,R2);
not not5038(N17495,R4);
not not5039(N17496,R7);
not not5040(N17504,in1);
not not5041(N17505,R1);
not not5042(N17506,R4);
not not5043(N17507,R6);
not not5044(N17515,in1);
not not5045(N17516,in2);
not not5046(N17517,R2);
not not5047(N17518,R6);
not not5048(N17526,in1);
not not5049(N17527,R4);
not not5050(N17528,R6);
not not5051(N17529,R7);
not not5052(N17537,in1);
not not5053(N17538,R2);
not not5054(N17539,R3);
not not5055(N17540,R7);
not not5056(N17548,in2);
not not5057(N17549,R0);
not not5058(N17550,R4);
not not5059(N17551,R5);
not not5060(N17559,in2);
not not5061(N17560,R0);
not not5062(N17561,R5);
not not5063(N17562,R6);
not not5064(N17570,in2);
not not5065(N17571,R1);
not not5066(N17572,R4);
not not5067(N17573,R6);
not not5068(N17581,in1);
not not5069(N17582,R2);
not not5070(N17583,R4);
not not5071(N17591,in1);
not not5072(N17592,R4);
not not5073(N17593,R7);
not not5074(N17601,in2);
not not5075(N17602,R2);
not not5076(N17603,R7);
not not5077(N17611,R2);
not not5078(N17612,R3);
not not5079(N17613,R6);
not not5080(N17621,in2);
not not5081(N17622,R2);
not not5082(N17623,R5);
not not5083(N17631,R0);
not not5084(N17632,R1);
not not5085(N17633,R5);
not not5086(N17641,in1);
not not5087(N17642,R2);
not not5088(N17643,R6);
not not5089(N11896,R4);
not not5090(N11897,R5);
not not5091(N11898,R6);
not not5092(N11899,R7);
not not5093(N11915,R4);
not not5094(N11916,R5);
not not5095(N11917,R7);
not not5096(N11932,R4);
not not5097(N11933,R5);
not not5098(N11934,R6);
not not5099(N11949,R4);
not not5100(N11950,R5);
not not5101(N11951,R6);
not not5102(N11966,R5);
not not5103(N11967,R6);
not not5104(N11968,R7);
not not5105(N11983,R3);
not not5106(N11984,R4);
not not5107(N11985,R5);
not not5108(N11998,R4);
not not5109(N11999,R5);
not not5110(N12000,R6);
not not5111(N12001,R7);
not not5112(N12016,R5);
not not5113(N12017,R6);
not not5114(N12031,R4);
not not5115(N12032,R5);
not not5116(N12033,R7);
not not5117(N12048,R4);
not not5118(N12049,R6);
not not5119(N12064,R4);
not not5120(N12065,R6);
not not5121(N12080,R4);
not not5122(N12081,R5);
not not5123(N12096,R5);
not not5124(N12097,R7);
not not5125(N12111,R4);
not not5126(N12112,R6);
not not5127(N12113,R7);
not not5128(N12128,R4);
not not5129(N12129,R7);
not not5130(N12143,R3);
not not5131(N12144,R5);
not not5132(N12145,R6);
not not5133(N12159,R4);
not not5134(N12160,R5);
not not5135(N12161,R7);
not not5136(N12175,R3);
not not5137(N12176,R5);
not not5138(N12177,R7);
not not5139(N12191,R4);
not not5140(N12192,R5);
not not5141(N12193,R6);
not not5142(N12206,R5);
not not5143(N12207,R6);
not not5144(N12208,R7);
not not5145(N12221,R5);
not not5146(N12222,R6);
not not5147(N12223,R7);
not not5148(N12236,R5);
not not5149(N12237,R6);
not not5150(N12238,R7);
not not5151(N12251,R4);
not not5152(N12252,R5);
not not5153(N12253,R6);
not not5154(N12267,R6);
not not5155(N12268,R7);
not not5156(N12281,R4);
not not5157(N12282,R5);
not not5158(N12283,R6);
not not5159(N12296,R4);
not not5160(N12297,R5);
not not5161(N12298,R7);
not not5162(N12312,R6);
not not5163(N12313,R7);
not not5164(N12327,R6);
not not5165(N12328,R7);
not not5166(N12342,R6);
not not5167(N12343,R7);
not not5168(N12356,R4);
not not5169(N12357,R5);
not not5170(N12358,R6);
not not5171(N12371,R4);
not not5172(N12372,R5);
not not5173(N12373,R6);
not not5174(N12385,R4);
not not5175(N12386,R5);
not not5176(N12387,R6);
not not5177(N12388,R7);
not not5178(N12401,R4);
not not5179(N12402,R5);
not not5180(N12403,R6);
not not5181(N12416,R4);
not not5182(N12417,R6);
not not5183(N12418,R7);
not not5184(N12431,R4);
not not5185(N12432,R6);
not not5186(N12433,R7);
not not5187(N12446,R4);
not not5188(N12447,R6);
not not5189(N12448,R7);
not not5190(N12462,R4);
not not5191(N12463,R7);
not not5192(N12477,R4);
not not5193(N12478,R6);
not not5194(N12492,R4);
not not5195(N12493,R6);
not not5196(N12507,R4);
not not5197(N12508,R5);
not not5198(N12522,R6);
not not5199(N12523,R7);
not not5200(N12537,R4);
not not5201(N12538,R6);
not not5202(N12552,R5);
not not5203(N12553,R6);
not not5204(N12567,R5);
not not5205(N12568,R7);
not not5206(N12581,R5);
not not5207(N12582,R6);
not not5208(N12583,R7);
not not5209(N12597,R5);
not not5210(N12598,R6);
not not5211(N12612,R6);
not not5212(N12613,R7);
not not5213(N12627,R6);
not not5214(N12628,R7);
not not5215(N12642,R5);
not not5216(N12643,R7);
not not5217(N12656,R5);
not not5218(N12657,R6);
not not5219(N12658,R7);
not not5220(N12671,R5);
not not5221(N12672,R6);
not not5222(N12673,R7);
not not5223(N12687,R5);
not not5224(N12688,R6);
not not5225(N12701,R3);
not not5226(N12702,R5);
not not5227(N12703,R7);
not not5228(N12716,R3);
not not5229(N12717,R4);
not not5230(N12718,R5);
not not5231(N12731,R4);
not not5232(N12732,R6);
not not5233(N12733,R7);
not not5234(N12746,R4);
not not5235(N12747,R6);
not not5236(N12748,R7);
not not5237(N12761,R5);
not not5238(N12762,R7);
not not5239(N12775,R5);
not not5240(N12776,R7);
not not5241(N12789,R5);
not not5242(N12790,R7);
not not5243(N12803,R5);
not not5244(N12804,R7);
not not5245(N12816,R4);
not not5246(N12817,R5);
not not5247(N12818,R7);
not not5248(N12831,R5);
not not5249(N12832,R7);
not not5250(N12845,R4);
not not5251(N12846,R7);
not not5252(N12860,R7);
not not5253(N12873,R4);
not not5254(N12874,R6);
not not5255(N12887,R4);
not not5256(N12888,R6);
not not5257(N12901,R4);
not not5258(N12902,R6);
not not5259(N12914,R3);
not not5260(N12915,R5);
not not5261(N12916,R7);
not not5262(N12929,R4);
not not5263(N12930,R5);
not not5264(N12944,R6);
not not5265(N12958,R6);
not not5266(N12971,R5);
not not5267(N12972,R6);
not not5268(N12985,R5);
not not5269(N12986,R7);
not not5270(N12999,R5);
not not5271(N13000,R6);
not not5272(N13014,R5);
not not5273(N13026,R4);
not not5274(N13027,R5);
not not5275(N13028,R6);
not not5276(N13040,R5);
not not5277(N13041,R6);
not not5278(N13042,R7);
not not5279(N13055,R5);
not not5280(N13056,R7);
not not5281(N13069,R4);
not not5282(N13070,R5);
not not5283(N13084,R5);
not not5284(N13098,R5);
not not5285(N13111,R5);
not not5286(N13112,R7);
not not5287(N13125,R3);
not not5288(N13126,R7);
not not5289(N13138,R4);
not not5290(N13139,R5);
not not5291(N13140,R6);
not not5292(N13153,R5);
not not5293(N13154,R6);
not not5294(N13167,R5);
not not5295(N13168,R6);
not not5296(N13182,R6);
not not5297(N13194,R3);
not not5298(N13195,R5);
not not5299(N13196,R7);
not not5300(N13209,R5);
not not5301(N13210,R7);
not not5302(N13223,R3);
not not5303(N13224,R7);
not not5304(N13238,R7);
not not5305(N13252,R7);
not not5306(N13266,R6);
not not5307(N13279,R3);
not not5308(N13280,R6);
not not5309(N13293,R5);
not not5310(N13294,R6);
not not5311(N13307,R5);
not not5312(N13308,R6);
not not5313(N13321,R5);
not not5314(N13322,R6);
not not5315(N13333,R5);
not not5316(N13334,R6);
not not5317(N13335,R7);
not not5318(N13346,R5);
not not5319(N13347,R6);
not not5320(N13348,R7);
not not5321(N13360,R4);
not not5322(N13361,R6);
not not5323(N13372,R5);
not not5324(N13373,R6);
not not5325(N13374,R7);
not not5326(N13386,R5);
not not5327(N13387,R6);
not not5328(N13399,R4);
not not5329(N13400,R5);
not not5330(N13411,R4);
not not5331(N13412,R5);
not not5332(N13413,R7);
not not5333(N13425,R6);
not not5334(N13426,R7);
not not5335(N13436,R3);
not not5336(N13437,R5);
not not5337(N13438,R6);
not not5338(N13439,R7);
not not5339(N13452,R6);
not not5340(N13464,R4);
not not5341(N13465,R7);
not not5342(N13477,R4);
not not5343(N13478,R6);
not not5344(N13490,R4);
not not5345(N13491,R6);
not not5346(N13503,R6);
not not5347(N13504,R7);
not not5348(N13516,R4);
not not5349(N13517,R7);
not not5350(N13529,R3);
not not5351(N13530,R7);
not not5352(N13543,R7);
not not5353(N13556,R6);
not not5354(N13568,R6);
not not5355(N13569,R7);
not not5356(N13582,R7);
not not5357(N13594,R6);
not not5358(N13595,R7);
not not5359(N13607,R5);
not not5360(N13608,R7);
not not5361(N13620,R5);
not not5362(N13621,R7);
not not5363(N13632,R4);
not not5364(N13633,R5);
not not5365(N13634,R6);
not not5366(N13647,R5);
not not5367(N13659,R6);
not not5368(N13660,R7);
not not5369(N13672,R5);
not not5370(N13673,R7);
not not5371(N13685,R5);
not not5372(N13686,R7);
not not5373(N13698,R3);
not not5374(N13699,R6);
not not5375(N13712,R5);
not not5376(N13725,R7);
not not5377(N13749,R4);
not not5378(N13750,R5);
not not5379(N13751,R6);
not not5380(N13763,R4);
not not5381(N13764,R6);
not not5382(N13775,R4);
not not5383(N13776,R5);
not not5384(N13777,R6);
not not5385(N13789,R5);
not not5386(N13790,R6);
not not5387(N13801,R3);
not not5388(N13802,R5);
not not5389(N13803,R6);
not not5390(N13815,R5);
not not5391(N13816,R7);
not not5392(N13828,R5);
not not5393(N13829,R7);
not not5394(N13841,R5);
not not5395(N13842,R7);
not not5396(N13854,R5);
not not5397(N13855,R7);
not not5398(N13867,R6);
not not5399(N13868,R7);
not not5400(N13880,R3);
not not5401(N13881,R7);
not not5402(N13893,R6);
not not5403(N13894,R7);
not not5404(N13906,R5);
not not5405(N13907,R6);
not not5406(N13919,R5);
not not5407(N13920,R6);
not not5408(N13932,R3);
not not5409(N13943,R4);
not not5410(N13944,R5);
not not5411(N13955,R5);
not not5412(N13956,R7);
not not5413(N13967,R5);
not not5414(N13968,R7);
not not5415(N13978,R4);
not not5416(N13979,R5);
not not5417(N13980,R7);
not not5418(N13992,R7);
not not5419(N14004,R5);
not not5420(N14015,R5);
not not5421(N14016,R6);
not not5422(N14027,R5);
not not5423(N14028,R6);
not not5424(N14040,R5);
not not5425(N14064,R4);
not not5426(N14087,R4);
not not5427(N14088,R5);
not not5428(N14100,R5);
not not5429(N14112,R7);
not not5430(N14123,R5);
not not5431(N14124,R7);
not not5432(N14135,R5);
not not5433(N14136,R7);
not not5434(N14148,R4);
not not5435(N14160,R4);
not not5436(N14172,R7);
not not5437(N14184,R7);
not not5438(N14196,R5);
not not5439(N14220,R5);
not not5440(N14231,R6);
not not5441(N14232,R7);
not not5442(N14244,R4);
not not5443(N14256,R3);
not not5444(N14266,R5);
not not5445(N14267,R7);
not not5446(N14278,R6);
not not5447(N14288,R4);
not not5448(N14289,R6);
not not5449(N14300,R7);
not not5450(N14310,R4);
not not5451(N14311,R7);
not not5452(N14333,R6);
not not5453(N14343,R6);
not not5454(N14344,R7);
not not5455(N14354,R6);
not not5456(N14355,R7);
not not5457(N14366,R6);
not not5458(N14377,R5);
not not5459(N14388,R5);
not not5460(N14399,R3);
not not5461(N14420,R3);
not not5462(N14421,R7);
not not5463(N14432,R7);
not not5464(N14442,R5);
not not5465(N14472,R4);
not not5466(N14492,R5);
not not5467(N14516,R6);
not not5468(N14517,R7);
not not5469(N14532,R6);
not not5470(N14533,R7);
not not5471(N14548,R6);
not not5472(N14549,R7);
not not5473(N14564,R6);
not not5474(N14579,R7);
not not5475(N14594,R7);
not not5476(N14608,R6);
not not5477(N14609,R7);
not not5478(N14624,R7);
not not5479(N14638,R6);
not not5480(N14639,R7);
not not5481(N14653,R6);
not not5482(N14654,R7);
not not5483(N14668,R5);
not not5484(N14669,R6);
not not5485(N14683,R6);
not not5486(N14684,R7);
not not5487(N14698,R6);
not not5488(N14699,R7);
not not5489(N14712,R6);
not not5490(N14713,R7);
not not5491(N14727,R6);
not not5492(N14741,R5);
not not5493(N14755,R6);
not not5494(N14769,R6);
not not5495(N14782,R6);
not not5496(N14783,R7);
not not5497(N14797,R7);
not not5498(N14810,R5);
not not5499(N14811,R6);
not not5500(N14825,R7);
not not5501(N14839,R5);
not not5502(N14853,R5);
not not5503(N14866,R6);
not not5504(N14867,R7);
not not5505(N14881,R7);
not not5506(N14894,R6);
not not5507(N14895,R7);
not not5508(N14909,R7);
not not5509(N14922,R6);
not not5510(N14923,R7);
not not5511(N14936,R6);
not not5512(N14937,R7);
not not5513(N14951,R6);
not not5514(N14964,R6);
not not5515(N14965,R7);
not not5516(N14978,R6);
not not5517(N14979,R7);
not not5518(N14993,R6);
not not5519(N15007,R6);
not not5520(N15020,R5);
not not5521(N15021,R6);
not not5522(N15035,R5);
not not5523(N15049,R6);
not not5524(N15062,R5);
not not5525(N15063,R6);
not not5526(N15077,R6);
not not5527(N15090,R6);
not not5528(N15091,R7);
not not5529(N15105,R7);
not not5530(N15119,R7);
not not5531(N15132,R6);
not not5532(N15133,R7);
not not5533(N15147,R7);
not not5534(N15160,R6);
not not5535(N15161,R7);
not not5536(N15174,R6);
not not5537(N15175,R7);
not not5538(N15188,R6);
not not5539(N15189,R7);
not not5540(N15201,R6);
not not5541(N15202,R7);
not not5542(N15214,R6);
not not5543(N15215,R7);
not not5544(N15228,R7);
not not5545(N15240,R6);
not not5546(N15241,R7);
not not5547(N15266,R6);
not not5548(N15267,R7);
not not5549(N15279,R6);
not not5550(N15280,R7);
not not5551(N15292,R6);
not not5552(N15293,R7);
not not5553(N15306,R7);
not not5554(N15319,R7);
not not5555(N15331,R6);
not not5556(N15332,R7);
not not5557(N15345,R7);
not not5558(N15358,R7);
not not5559(N15370,R6);
not not5560(N15371,R7);
not not5561(N15384,R7);
not not5562(N15397,R6);
not not5563(N15410,R7);
not not5564(N15422,R6);
not not5565(N15423,R7);
not not5566(N15435,R6);
not not5567(N15436,R7);
not not5568(N15449,R7);
not not5569(N15462,R7);
not not5570(N15475,R6);
not not5571(N15487,R6);
not not5572(N15488,R7);
not not5573(N15500,R6);
not not5574(N15501,R7);
not not5575(N15514,R7);
not not5576(N15527,R6);
not not5577(N15553,R5);
not not5578(N15565,R6);
not not5579(N15566,R7);
not not5580(N15578,R5);
not not5581(N15579,R7);
not not5582(N15592,R6);
not not5583(N15605,R6);
not not5584(N15618,R7);
not not5585(N15631,R6);
not not5586(N15643,R6);
not not5587(N15644,R7);
not not5588(N15657,R6);
not not5589(N15683,R5);
not not5590(N15695,R5);
not not5591(N15696,R7);
not not5592(N15709,R6);
not not5593(N15722,R6);
not not5594(N15734,R5);
not not5595(N15735,R6);
not not5596(N15748,R6);
not not5597(N15761,R6);
not not5598(N15773,R5);
not not5599(N15774,R7);
not not5600(N15786,R6);
not not5601(N15787,R7);
not not5602(N15813,R6);
not not5603(N15836,R6);
not not5604(N15837,R7);
not not5605(N15849,R5);
not not5606(N15861,R6);
not not5607(N15873,R5);
not not5608(N15885,R7);
not not5609(N15921,R6);
not not5610(N15933,R7);
not not5611(N15945,R7);
not not5612(N15956,R6);
not not5613(N15957,R7);
not not5614(N15969,R7);
not not5615(N15981,R6);
not not5616(N16017,R6);
not not5617(N16041,R6);
not not5618(N16053,R6);
not not5619(N16076,R4);
not not5620(N16077,R6);
not not5621(N16088,R6);
not not5622(N16089,R7);
not not5623(N16101,R6);
not not5624(N16113,R7);
not not5625(N16125,R5);
not not5626(N16173,R5);
not not5627(N16185,R5);
not not5628(N16197,R6);
not not5629(N16208,R6);
not not5630(N16209,R7);
not not5631(N16232,R6);
not not5632(N16233,R7);
not not5633(N16245,R6);
not not5634(N16257,R7);
not not5635(N16268,R6);
not not5636(N16269,R7);
not not5637(N16281,R6);
not not5638(N16293,R7);
not not5639(N16305,R6);
not not5640(N16329,R7);
not not5641(N16340,R5);
not not5642(N16341,R7);
not not5643(N16353,R6);
not not5644(N16377,R7);
not not5645(N16389,R6);
not not5646(N16401,R6);
not not5647(N16412,R6);
not not5648(N16413,R7);
not not5649(N16424,R6);
not not5650(N16425,R7);
not not5651(N16436,R6);
not not5652(N16437,R7);
not not5653(N16449,R4);
not not5654(N16470,R5);
not not5655(N16471,R7);
not not5656(N16481,R5);
not not5657(N16482,R7);
not not5658(N16493,R6);
not not5659(N16504,R6);
not not5660(N16526,R6);
not not5661(N16537,R4);
not not5662(N16548,R7);
not not5663(N16559,R7);
not not5664(N16570,R7);
not not5665(N16592,R7);
not not5666(N16603,R7);
not not5667(N16614,R5);
not not5668(N16625,R6);
not not5669(N16647,R6);
not not5670(N16669,R6);
not not5671(N16680,R6);
not not5672(N16691,R5);
not not5673(N16724,R6);
not not5674(N16746,R7);
not not5675(N16757,R6);
not not5676(N16779,R7);
not not5677(N16790,R6);
not not5678(N16801,R7);
not not5679(N16823,R7);
not not5680(N16834,R7);
not not5681(N16866,R6);
not not5682(N16867,R7);
not not5683(N16877,R6);
not not5684(N16878,R7);
not not5685(N16899,R6);
not not5686(N16929,R6);
not not5687(N16959,R7);
not not5688(N16969,R6);
not not5689(N16979,R6);
not not5690(N16989,R6);
not not5691(N16999,R6);
not not5692(N17039,R5);
not not5693(N17059,R6);
not not5694(N18119,in0);
not not5695(N18120,in2);
not not5696(N18121,R0);
not not5697(N18122,R2);
not not5698(N18123,R3);
not not5699(N18137,in1);
not not5700(N18138,in2);
not not5701(N18139,R1);
not not5702(N18140,R2);
not not5703(N18141,R3);
not not5704(N18154,in0);
not not5705(N18155,R0);
not not5706(N18156,R1);
not not5707(N18157,R2);
not not5708(N18158,R3);
not not5709(N18171,in0);
not not5710(N18172,in1);
not not5711(N18173,R0);
not not5712(N18174,R1);
not not5713(N18175,R3);
not not5714(N18188,in1);
not not5715(N18189,R0);
not not5716(N18190,R1);
not not5717(N18191,R2);
not not5718(N18192,R3);
not not5719(N18205,in0);
not not5720(N18206,in1);
not not5721(N18207,in2);
not not5722(N18208,R0);
not not5723(N18209,R1);
not not5724(N18210,R2);
not not5725(N18222,in0);
not not5726(N18223,in1);
not not5727(N18224,in2);
not not5728(N18225,R1);
not not5729(N18226,R2);
not not5730(N18239,in0);
not not5731(N18240,R0);
not not5732(N18241,R2);
not not5733(N18255,in1);
not not5734(N18256,R0);
not not5735(N18257,R1);
not not5736(N18258,R2);
not not5737(N18259,R3);
not not5738(N18271,in0);
not not5739(N18272,R0);
not not5740(N18273,R1);
not not5741(N18274,R2);
not not5742(N18287,in2);
not not5743(N18288,R0);
not not5744(N18289,R1);
not not5745(N18290,R3);
not not5746(N18303,in1);
not not5747(N18304,R0);
not not5748(N18305,R1);
not not5749(N18306,R3);
not not5750(N18319,in1);
not not5751(N18320,in2);
not not5752(N18321,R0);
not not5753(N18322,R2);
not not5754(N18335,in0);
not not5755(N18336,in1);
not not5756(N18337,in2);
not not5757(N18338,R3);
not not5758(N18351,in0);
not not5759(N18352,in1);
not not5760(N18353,in2);
not not5761(N18354,R0);
not not5762(N18367,in0);
not not5763(N18368,in1);
not not5764(N18369,in2);
not not5765(N18370,R0);
not not5766(N18371,R3);
not not5767(N18383,in0);
not not5768(N18384,R0);
not not5769(N18385,R2);
not not5770(N18386,R3);
not not5771(N18399,in0);
not not5772(N18400,in1);
not not5773(N18401,R1);
not not5774(N18415,in0);
not not5775(N18416,R1);
not not5776(N18417,R3);
not not5777(N18431,in0);
not not5778(N18432,in1);
not not5779(N18433,in2);
not not5780(N18434,R1);
not not5781(N18447,in0);
not not5782(N18448,in2);
not not5783(N18449,R2);
not not5784(N18450,R3);
not not5785(N18463,in1);
not not5786(N18464,R0);
not not5787(N18465,R1);
not not5788(N18466,R2);
not not5789(N18479,in0);
not not5790(N18480,in1);
not not5791(N18481,R1);
not not5792(N18482,R3);
not not5793(N18495,in0);
not not5794(N18496,in2);
not not5795(N18497,R1);
not not5796(N18498,R2);
not not5797(N18511,in1);
not not5798(N18512,in2);
not not5799(N18513,R0);
not not5800(N18514,R2);
not not5801(N18527,in0);
not not5802(N18528,in1);
not not5803(N18529,R0);
not not5804(N18530,R2);
not not5805(N18543,in0);
not not5806(N18544,in1);
not not5807(N18545,in2);
not not5808(N18546,R1);
not not5809(N18547,R3);
not not5810(N18559,in1);
not not5811(N18560,in2);
not not5812(N18561,R2);
not not5813(N18562,R3);
not not5814(N18574,in0);
not not5815(N18575,in1);
not not5816(N18589,in1);
not not5817(N18590,in2);
not not5818(N18591,R1);
not not5819(N18604,in1);
not not5820(N18605,R3);
not not5821(N18619,in1);
not not5822(N18620,in2);
not not5823(N18621,R0);
not not5824(N18622,R2);
not not5825(N18634,in2);
not not5826(N18635,R0);
not not5827(N18636,R1);
not not5828(N18649,in0);
not not5829(N18650,R2);
not not5830(N18651,R3);
not not5831(N18664,in1);
not not5832(N18665,R2);
not not5833(N18666,R3);
not not5834(N18679,in0);
not not5835(N18680,in2);
not not5836(N18681,R0);
not not5837(N18682,R1);
not not5838(N18694,in0);
not not5839(N18695,in1);
not not5840(N18696,R0);
not not5841(N18709,in0);
not not5842(N18710,in1);
not not5843(N18711,in2);
not not5844(N18712,R3);
not not5845(N18724,in1);
not not5846(N18725,in2);
not not5847(N18726,R0);
not not5848(N18727,R2);
not not5849(N18739,in0);
not not5850(N18740,R3);
not not5851(N18754,in2);
not not5852(N18755,R3);
not not5853(N18769,in2);
not not5854(N18770,R1);
not not5855(N18784,in1);
not not5856(N18785,R0);
not not5857(N18786,R1);
not not5858(N18787,R2);
not not5859(N18799,in2);
not not5860(N18800,R0);
not not5861(N18801,R1);
not not5862(N18802,R2);
not not5863(N18814,in0);
not not5864(N18815,R0);
not not5865(N18816,R2);
not not5866(N18817,R3);
not not5867(N18829,R0);
not not5868(N18830,R2);
not not5869(N18831,R3);
not not5870(N18844,in1);
not not5871(N18845,in2);
not not5872(N18846,R1);
not not5873(N18859,in0);
not not5874(N18860,in1);
not not5875(N18861,in2);
not not5876(N18862,R2);
not not5877(N18874,in0);
not not5878(N18875,R2);
not not5879(N18876,R3);
not not5880(N18889,in0);
not not5881(N18890,in1);
not not5882(N18891,in2);
not not5883(N18904,in1);
not not5884(N18905,in2);
not not5885(N18906,R2);
not not5886(N18907,R3);
not not5887(N18919,in1);
not not5888(N18920,R0);
not not5889(N18933,in2);
not not5890(N18934,R3);
not not5891(N18947,R1);
not not5892(N18948,R3);
not not5893(N18961,R1);
not not5894(N18962,R2);
not not5895(N18975,in0);
not not5896(N18976,in1);
not not5897(N18989,in2);
not not5898(N18990,R0);
not not5899(N18991,R2);
not not5900(N19003,in1);
not not5901(N19004,R0);
not not5902(N19005,R2);
not not5903(N19017,R0);
not not5904(N19018,R2);
not not5905(N19031,in2);
not not5906(N19032,R0);
not not5907(N19033,R2);
not not5908(N19045,in0);
not not5909(N19046,R2);
not not5910(N19047,R3);
not not5911(N19059,in1);
not not5912(N19060,R2);
not not5913(N19061,R3);
not not5914(N19073,in2);
not not5915(N19074,R0);
not not5916(N19075,R3);
not not5917(N19087,in0);
not not5918(N19088,R0);
not not5919(N19089,R1);
not not5920(N19101,in0);
not not5921(N19102,in1);
not not5922(N19103,in2);
not not5923(N19104,R2);
not not5924(N19115,in0);
not not5925(N19116,in1);
not not5926(N19117,R2);
not not5927(N19129,R0);
not not5928(N19130,R1);
not not5929(N19131,R3);
not not5930(N19143,in2);
not not5931(N19144,R0);
not not5932(N19145,R3);
not not5933(N19157,in1);
not not5934(N19158,in2);
not not5935(N19159,R1);
not not5936(N19160,R3);
not not5937(N19171,R0);
not not5938(N19172,R1);
not not5939(N19185,in0);
not not5940(N19186,R0);
not not5941(N19199,in1);
not not5942(N19200,R3);
not not5943(N19213,in1);
not not5944(N19214,R0);
not not5945(N19215,R2);
not not5946(N19216,R3);
not not5947(N19227,R0);
not not5948(N19228,R1);
not not5949(N19229,R2);
not not5950(N19241,in2);
not not5951(N19242,R1);
not not5952(N19243,R2);
not not5953(N19255,in0);
not not5954(N19256,in2);
not not5955(N19257,R1);
not not5956(N19269,in1);
not not5957(N19270,R0);
not not5958(N19271,R2);
not not5959(N19283,in1);
not not5960(N19284,in2);
not not5961(N19285,R0);
not not5962(N19297,in2);
not not5963(N19298,R0);
not not5964(N19299,R2);
not not5965(N19311,in2);
not not5966(N19312,R0);
not not5967(N19313,R1);
not not5968(N19314,R3);
not not5969(N19325,in2);
not not5970(N19326,R0);
not not5971(N19327,R1);
not not5972(N19339,R1);
not not5973(N19340,R2);
not not5974(N19341,R3);
not not5975(N19353,in1);
not not5976(N19354,R1);
not not5977(N19355,R2);
not not5978(N19367,in0);
not not5979(N19368,R3);
not not5980(N19381,R0);
not not5981(N19382,R1);
not not5982(N19383,R2);
not not5983(N19395,in0);
not not5984(N19396,in1);
not not5985(N19397,in2);
not not5986(N19409,in0);
not not5987(N19410,in1);
not not5988(N19411,in2);
not not5989(N19412,R3);
not not5990(N19423,in1);
not not5991(N19424,in2);
not not5992(N19425,R0);
not not5993(N19426,R3);
not not5994(N19437,in0);
not not5995(N19438,in2);
not not5996(N19439,R0);
not not5997(N19440,R1);
not not5998(N19451,in0);
not not5999(N19452,R0);
not not6000(N19465,in0);
not not6001(N19466,R0);
not not6002(N19479,in1);
not not6003(N19480,in2);
not not6004(N19481,R2);
not not6005(N19493,in2);
not not6006(N19494,R2);
not not6007(N19507,in0);
not not6008(N19508,in2);
not not6009(N19509,R1);
not not6010(N19521,in1);
not not6011(N19522,in2);
not not6012(N19523,R1);
not not6013(N19535,in0);
not not6014(N19536,in1);
not not6015(N19537,R1);
not not6016(N19549,in0);
not not6017(N19550,in1);
not not6018(N19551,R0);
not not6019(N19563,in0);
not not6020(N19564,in2);
not not6021(N19565,R1);
not not6022(N19566,R2);
not not6023(N19577,in0);
not not6024(N19578,in1);
not not6025(N19579,R2);
not not6026(N19591,in0);
not not6027(N19592,in1);
not not6028(N19605,in0);
not not6029(N19606,in1);
not not6030(N19607,R2);
not not6031(N19619,in0);
not not6032(N19620,in1);
not not6033(N19621,in2);
not not6034(N19622,R0);
not not6035(N19633,in2);
not not6036(N19634,R0);
not not6037(N19635,R1);
not not6038(N19647,in0);
not not6039(N19648,R0);
not not6040(N19661,in2);
not not6041(N19662,R3);
not not6042(N19675,in1);
not not6043(N19676,in2);
not not6044(N19677,R1);
not not6045(N19678,R2);
not not6046(N19689,in1);
not not6047(N19690,R0);
not not6048(N19691,R1);
not not6049(N19703,in0);
not not6050(N19704,in1);
not not6051(N19705,R0);
not not6052(N19717,in2);
not not6053(N19718,R0);
not not6054(N19719,R1);
not not6055(N19731,R0);
not not6056(N19732,R2);
not not6057(N19744,R2);
not not6058(N19757,in0);
not not6059(N19758,R2);
not not6060(N19770,in1);
not not6061(N19771,in2);
not not6062(N19772,R0);
not not6063(N19773,R3);
not not6064(N19783,R1);
not not6065(N19784,R2);
not not6066(N19796,in0);
not not6067(N19797,R1);
not not6068(N19809,R1);
not not6069(N19822,in2);
not not6070(N19823,R1);
not not6071(N19835,in0);
not not6072(N19836,R1);
not not6073(N19848,in0);
not not6074(N19849,in2);
not not6075(N19850,R1);
not not6076(N19861,R0);
not not6077(N19874,in1);
not not6078(N19875,R1);
not not6079(N19876,R2);
not not6080(N19887,in0);
not not6081(N19888,in1);
not not6082(N19889,R3);
not not6083(N19900,in0);
not not6084(N19901,R1);
not not6085(N19902,R2);
not not6086(N19913,in1);
not not6087(N19914,R0);
not not6088(N19926,in0);
not not6089(N19927,R0);
not not6090(N19939,R0);
not not6091(N19940,R3);
not not6092(N19952,in0);
not not6093(N19953,in1);
not not6094(N19954,R2);
not not6095(N19965,in0);
not not6096(N19966,R0);
not not6097(N19967,R2);
not not6098(N19978,in0);
not not6099(N19979,in1);
not not6100(N19980,R3);
not not6101(N19991,in0);
not not6102(N19992,in1);
not not6103(N20004,R0);
not not6104(N20005,R1);
not not6105(N20006,R2);
not not6106(N20017,in0);
not not6107(N20018,R0);
not not6108(N20019,R1);
not not6109(N20030,R1);
not not6110(N20031,R2);
not not6111(N20043,in0);
not not6112(N20044,R0);
not not6113(N20056,in1);
not not6114(N20057,R0);
not not6115(N20069,in2);
not not6116(N20070,R2);
not not6117(N20082,in1);
not not6118(N20083,R2);
not not6119(N20095,in0);
not not6120(N20096,in1);
not not6121(N20097,in2);
not not6122(N20108,in0);
not not6123(N20109,R3);
not not6124(N20121,in0);
not not6125(N20122,in2);
not not6126(N20123,R0);
not not6127(N20134,in0);
not not6128(N20135,R0);
not not6129(N20136,R3);
not not6130(N20147,in1);
not not6131(N20148,R2);
not not6132(N20160,in0);
not not6133(N20161,in1);
not not6134(N20162,in2);
not not6135(N20173,in0);
not not6136(N20174,R0);
not not6137(N20175,R1);
not not6138(N20186,in0);
not not6139(N20187,in2);
not not6140(N20199,in1);
not not6141(N20200,R3);
not not6142(N20212,in2);
not not6143(N20213,R3);
not not6144(N20225,in0);
not not6145(N20226,in1);
not not6146(N20227,in2);
not not6147(N20238,R1);
not not6148(N20239,R2);
not not6149(N20251,R2);
not not6150(N20263,R2);
not not6151(N20275,in2);
not not6152(N20276,R0);
not not6153(N20287,in0);
not not6154(N20288,R0);
not not6155(N20299,R2);
not not6156(N20311,R0);
not not6157(N20312,R2);
not not6158(N20323,R3);
not not6159(N20335,in0);
not not6160(N20347,in2);
not not6161(N20348,R1);
not not6162(N20359,R1);
not not6163(N20371,in0);
not not6164(N20372,R3);
not not6165(N20383,in2);
not not6166(N20407,in2);
not not6167(N20419,R0);
not not6168(N20420,R2);
not not6169(N20431,in2);
not not6170(N20432,R2);
not not6171(N20443,in1);
not not6172(N20467,in0);
not not6173(N20479,in1);
not not6174(N20480,R1);
not not6175(N20491,in0);
not not6176(N20492,in1);
not not6177(N20493,R2);
not not6178(N20503,in1);
not not6179(N20515,R3);
not not6180(N20527,in1);
not not6181(N20528,R0);
not not6182(N20529,R2);
not not6183(N20539,in1);
not not6184(N20540,R1);
not not6185(N20551,in2);
not not6186(N20552,R1);
not not6187(N20563,R0);
not not6188(N20564,R2);
not not6189(N20575,in0);
not not6190(N20576,R0);
not not6191(N20577,R2);
not not6192(N20587,in2);
not not6193(N20588,R2);
not not6194(N20599,in0);
not not6195(N20600,in1);
not not6196(N20611,R0);
not not6197(N20612,R1);
not not6198(N20623,R3);
not not6199(N20635,in2);
not not6200(N20647,R1);
not not6201(N20659,R0);
not not6202(N20682,R2);
not not6203(N20693,R2);
not not6204(N20704,R0);
not not6205(N20715,in0);
not not6206(N20716,R0);
not not6207(N20726,in0);
not not6208(N20747,R2);
not not6209(N20757,R0);
not not6210(N20777,R1);
not not6211(N20827,R2);
not not6212(N20847,R1);
not not6213(N20856,in0);
not not6214(N20857,R0);
not not6215(N20858,R2);
not not6216(N20859,R3);
not not6217(N20860,R4);
not not6218(N20861,R5);
not not6219(N20872,in0);
not not6220(N20873,in2);
not not6221(N20874,R0);
not not6222(N20875,R1);
not not6223(N20876,R2);
not not6224(N20877,R3);
not not6225(N20888,in0);
not not6226(N20889,in2);
not not6227(N20890,R1);
not not6228(N20891,R2);
not not6229(N20892,R3);
not not6230(N20903,in0);
not not6231(N20904,in1);
not not6232(N20905,in2);
not not6233(N20906,R1);
not not6234(N20907,R2);
not not6235(N20908,R5);
not not6236(N20918,in0);
not not6237(N20919,in2);
not not6238(N20920,R1);
not not6239(N20921,R2);
not not6240(N20922,R4);
not not6241(N20933,in0);
not not6242(N20934,in2);
not not6243(N20935,R1);
not not6244(N20936,R3);
not not6245(N20937,R4);
not not6246(N20938,R5);
not not6247(N20948,in0);
not not6248(N20949,in1);
not not6249(N20950,R0);
not not6250(N20951,R1);
not not6251(N20952,R3);
not not6252(N20953,R5);
not not6253(N20963,in1);
not not6254(N20964,in2);
not not6255(N20965,R3);
not not6256(N20966,R4);
not not6257(N20967,R5);
not not6258(N20978,in2);
not not6259(N20979,R0);
not not6260(N20980,R1);
not not6261(N20981,R2);
not not6262(N20982,R3);
not not6263(N20993,in0);
not not6264(N20994,in2);
not not6265(N20995,R0);
not not6266(N20996,R2);
not not6267(N20997,R4);
not not6268(N21008,in1);
not not6269(N21009,in2);
not not6270(N21010,R1);
not not6271(N21011,R2);
not not6272(N21012,R4);
not not6273(N21023,in1);
not not6274(N21024,R1);
not not6275(N21025,R2);
not not6276(N21026,R3);
not not6277(N21027,R4);
not not6278(N21038,in2);
not not6279(N21039,R1);
not not6280(N21040,R2);
not not6281(N21041,R3);
not not6282(N21042,R4);
not not6283(N21053,in0);
not not6284(N21054,in2);
not not6285(N21055,R0);
not not6286(N21056,R1);
not not6287(N21057,R3);
not not6288(N21058,R5);
not not6289(N21068,in0);
not not6290(N21069,R0);
not not6291(N21070,R1);
not not6292(N21071,R2);
not not6293(N21072,R3);
not not6294(N21083,in1);
not not6295(N21084,in2);
not not6296(N21085,R0);
not not6297(N21086,R5);
not not6298(N21097,in2);
not not6299(N21098,R0);
not not6300(N21099,R4);
not not6301(N21100,R5);
not not6302(N21111,in1);
not not6303(N21112,R0);
not not6304(N21113,R4);
not not6305(N21114,R5);
not not6306(N21125,in1);
not not6307(N21126,in2);
not not6308(N21127,R0);
not not6309(N21128,R3);
not not6310(N21139,in2);
not not6311(N21140,R1);
not not6312(N21141,R3);
not not6313(N21142,R4);
not not6314(N21143,R5);
not not6315(N21153,in1);
not not6316(N21154,R1);
not not6317(N21155,R3);
not not6318(N21156,R4);
not not6319(N21157,R5);
not not6320(N21167,in0);
not not6321(N21168,R0);
not not6322(N21169,R1);
not not6323(N21170,R4);
not not6324(N21181,in2);
not not6325(N21182,R0);
not not6326(N21183,R1);
not not6327(N21184,R4);
not not6328(N21195,in1);
not not6329(N21196,R0);
not not6330(N21197,R2);
not not6331(N21198,R4);
not not6332(N21199,R5);
not not6333(N21209,in1);
not not6334(N21210,R1);
not not6335(N21211,R3);
not not6336(N21212,R4);
not not6337(N21213,R5);
not not6338(N21223,in1);
not not6339(N21224,in2);
not not6340(N21225,R1);
not not6341(N21226,R2);
not not6342(N21227,R4);
not not6343(N21237,in0);
not not6344(N21238,in1);
not not6345(N21239,in2);
not not6346(N21240,R0);
not not6347(N21241,R4);
not not6348(N21251,R0);
not not6349(N21252,R1);
not not6350(N21253,R2);
not not6351(N21254,R3);
not not6352(N21255,R5);
not not6353(N21265,in1);
not not6354(N21266,in2);
not not6355(N21267,R0);
not not6356(N21268,R2);
not not6357(N21279,in2);
not not6358(N21280,R2);
not not6359(N21281,R3);
not not6360(N21282,R5);
not not6361(N21293,in2);
not not6362(N21294,R2);
not not6363(N21295,R3);
not not6364(N21296,R5);
not not6365(N21307,in2);
not not6366(N21308,R1);
not not6367(N21309,R2);
not not6368(N21310,R5);
not not6369(N21321,in0);
not not6370(N21322,in1);
not not6371(N21323,R0);
not not6372(N21324,R2);
not not6373(N21325,R3);
not not6374(N21335,in0);
not not6375(N21336,in1);
not not6376(N21337,R0);
not not6377(N21338,R2);
not not6378(N21339,R5);
not not6379(N21349,in0);
not not6380(N21350,in1);
not not6381(N21351,R2);
not not6382(N21352,R3);
not not6383(N21363,in2);
not not6384(N21364,R1);
not not6385(N21365,R2);
not not6386(N21366,R3);
not not6387(N21377,in1);
not not6388(N21378,R2);
not not6389(N21379,R4);
not not6390(N21380,R5);
not not6391(N21391,in1);
not not6392(N21392,in2);
not not6393(N21393,R1);
not not6394(N21394,R3);
not not6395(N21395,R4);
not not6396(N21405,in0);
not not6397(N21406,in1);
not not6398(N21407,R0);
not not6399(N21408,R5);
not not6400(N21419,in2);
not not6401(N21420,R1);
not not6402(N21421,R3);
not not6403(N21422,R4);
not not6404(N21423,R5);
not not6405(N21433,in0);
not not6406(N21434,in1);
not not6407(N21435,in2);
not not6408(N21436,R2);
not not6409(N21437,R4);
not not6410(N21447,in1);
not not6411(N21448,in2);
not not6412(N21449,R1);
not not6413(N21450,R3);
not not6414(N21451,R5);
not not6415(N21461,in1);
not not6416(N21462,in2);
not not6417(N21463,R3);
not not6418(N21464,R5);
not not6419(N21475,in1);
not not6420(N21476,R0);
not not6421(N21477,R2);
not not6422(N21478,R3);
not not6423(N21489,in2);
not not6424(N21490,R0);
not not6425(N21491,R2);
not not6426(N21492,R3);
not not6427(N21503,in0);
not not6428(N21504,in1);
not not6429(N21505,in2);
not not6430(N21506,R0);
not not6431(N21507,R5);
not not6432(N21517,R1);
not not6433(N21518,R2);
not not6434(N21519,R3);
not not6435(N21520,R4);
not not6436(N21531,in0);
not not6437(N21532,in2);
not not6438(N21533,R5);
not not6439(N21544,in2);
not not6440(N21545,R2);
not not6441(N21546,R3);
not not6442(N21547,R4);
not not6443(N21557,in1);
not not6444(N21558,in2);
not not6445(N21559,R5);
not not6446(N21570,in2);
not not6447(N21571,R1);
not not6448(N21572,R2);
not not6449(N21573,R5);
not not6450(N21583,R0);
not not6451(N21584,R1);
not not6452(N21585,R2);
not not6453(N21596,in0);
not not6454(N21597,in1);
not not6455(N21598,in2);
not not6456(N21599,R2);
not not6457(N21609,in0);
not not6458(N21610,R1);
not not6459(N21611,R2);
not not6460(N21612,R5);
not not6461(N21622,in1);
not not6462(N21623,R1);
not not6463(N21624,R2);
not not6464(N21625,R4);
not not6465(N21635,in1);
not not6466(N21636,R0);
not not6467(N21637,R1);
not not6468(N21638,R4);
not not6469(N21648,in0);
not not6470(N21649,in1);
not not6471(N21650,R2);
not not6472(N21651,R4);
not not6473(N21661,in0);
not not6474(N21662,in2);
not not6475(N21663,R0);
not not6476(N21674,R2);
not not6477(N21675,R4);
not not6478(N21676,R5);
not not6479(N21687,in0);
not not6480(N21688,in1);
not not6481(N21689,R0);
not not6482(N21690,R2);
not not6483(N21691,R5);
not not6484(N21700,in1);
not not6485(N21701,in2);
not not6486(N21702,R3);
not not6487(N21703,R4);
not not6488(N21704,R5);
not not6489(N21713,in1);
not not6490(N21714,in2);
not not6491(N21715,R1);
not not6492(N21716,R4);
not not6493(N21717,R5);
not not6494(N21726,in1);
not not6495(N21727,R0);
not not6496(N21728,R3);
not not6497(N21729,R4);
not not6498(N21739,in0);
not not6499(N21740,in1);
not not6500(N21741,R3);
not not6501(N21742,R4);
not not6502(N21752,in0);
not not6503(N21753,R1);
not not6504(N21754,R2);
not not6505(N21755,R5);
not not6506(N21765,in1);
not not6507(N21766,R0);
not not6508(N21767,R2);
not not6509(N21768,R5);
not not6510(N21778,in2);
not not6511(N21779,R0);
not not6512(N21780,R2);
not not6513(N21781,R5);
not not6514(N21791,in0);
not not6515(N21792,R1);
not not6516(N21793,R2);
not not6517(N21794,R5);
not not6518(N21804,R1);
not not6519(N21805,R3);
not not6520(N21806,R5);
not not6521(N21817,in2);
not not6522(N21818,R0);
not not6523(N21819,R3);
not not6524(N21820,R4);
not not6525(N21830,in2);
not not6526(N21831,R0);
not not6527(N21832,R3);
not not6528(N21833,R4);
not not6529(N21843,in1);
not not6530(N21844,in2);
not not6531(N21845,R0);
not not6532(N21846,R1);
not not6533(N21847,R5);
not not6534(N21856,in1);
not not6535(N21857,in2);
not not6536(N21858,R2);
not not6537(N21859,R3);
not not6538(N21869,R0);
not not6539(N21870,R2);
not not6540(N21871,R3);
not not6541(N21882,in1);
not not6542(N21883,R0);
not not6543(N21884,R3);
not not6544(N21885,R5);
not not6545(N21895,R1);
not not6546(N21896,R2);
not not6547(N21897,R4);
not not6548(N21898,R5);
not not6549(N21908,R1);
not not6550(N21909,R2);
not not6551(N21910,R4);
not not6552(N21911,R5);
not not6553(N21921,R1);
not not6554(N21922,R2);
not not6555(N21923,R4);
not not6556(N21924,R5);
not not6557(N21934,in0);
not not6558(N21935,in2);
not not6559(N21936,R2);
not not6560(N21937,R3);
not not6561(N21938,R5);
not not6562(N21947,in1);
not not6563(N21948,R0);
not not6564(N21949,R1);
not not6565(N21950,R4);
not not6566(N21951,R5);
not not6567(N21960,in1);
not not6568(N21961,R0);
not not6569(N21962,R2);
not not6570(N21963,R3);
not not6571(N21973,in2);
not not6572(N21974,R0);
not not6573(N21975,R2);
not not6574(N21976,R3);
not not6575(N21986,in1);
not not6576(N21987,R0);
not not6577(N21988,R2);
not not6578(N21989,R4);
not not6579(N21999,in2);
not not6580(N22000,R0);
not not6581(N22001,R2);
not not6582(N22002,R4);
not not6583(N22012,R0);
not not6584(N22013,R2);
not not6585(N22014,R4);
not not6586(N22015,R5);
not not6587(N22025,in2);
not not6588(N22026,R0);
not not6589(N22027,R1);
not not6590(N22028,R4);
not not6591(N22038,in1);
not not6592(N22039,R0);
not not6593(N22040,R1);
not not6594(N22041,R4);
not not6595(N22051,in1);
not not6596(N22052,R0);
not not6597(N22053,R1);
not not6598(N22054,R4);
not not6599(N22064,in0);
not not6600(N22065,R1);
not not6601(N22066,R4);
not not6602(N22077,in1);
not not6603(N22078,R0);
not not6604(N22079,R1);
not not6605(N22080,R3);
not not6606(N22090,in1);
not not6607(N22091,R0);
not not6608(N22092,R1);
not not6609(N22093,R3);
not not6610(N22103,in1);
not not6611(N22104,R0);
not not6612(N22105,R3);
not not6613(N22116,R1);
not not6614(N22117,R3);
not not6615(N22118,R4);
not not6616(N22119,R5);
not not6617(N22129,in2);
not not6618(N22130,R0);
not not6619(N22131,R4);
not not6620(N22142,in0);
not not6621(N22143,in2);
not not6622(N22144,R3);
not not6623(N22145,R4);
not not6624(N22155,in1);
not not6625(N22156,R1);
not not6626(N22157,R2);
not not6627(N22158,R4);
not not6628(N22168,R2);
not not6629(N22169,R3);
not not6630(N22170,R4);
not not6631(N22181,R1);
not not6632(N22182,R2);
not not6633(N22183,R3);
not not6634(N22184,R5);
not not6635(N22194,in0);
not not6636(N22195,R0);
not not6637(N22196,R2);
not not6638(N22197,R3);
not not6639(N22207,in0);
not not6640(N22208,R0);
not not6641(N22209,R2);
not not6642(N22210,R3);
not not6643(N22220,R2);
not not6644(N22221,R3);
not not6645(N22222,R5);
not not6646(N22233,in1);
not not6647(N22234,in2);
not not6648(N22235,R0);
not not6649(N22245,in2);
not not6650(N22246,R0);
not not6651(N22257,R1);
not not6652(N22258,R5);
not not6653(N22269,in2);
not not6654(N22270,R0);
not not6655(N22271,R2);
not not6656(N22272,R5);
not not6657(N22281,in1);
not not6658(N22282,R1);
not not6659(N22283,R3);
not not6660(N22293,in2);
not not6661(N22294,R1);
not not6662(N22295,R5);
not not6663(N22305,R0);
not not6664(N22306,R5);
not not6665(N22317,R4);
not not6666(N22318,R5);
not not6667(N22329,in0);
not not6668(N22330,R0);
not not6669(N22331,R4);
not not6670(N22341,R2);
not not6671(N22342,R3);
not not6672(N22343,R4);
not not6673(N22353,in2);
not not6674(N22354,R0);
not not6675(N22355,R3);
not not6676(N22365,in1);
not not6677(N22366,R3);
not not6678(N22367,R4);
not not6679(N22377,in1);
not not6680(N22378,R3);
not not6681(N22379,R4);
not not6682(N22389,R0);
not not6683(N22390,R2);
not not6684(N22391,R3);
not not6685(N22401,in0);
not not6686(N22402,R1);
not not6687(N22403,R2);
not not6688(N22404,R5);
not not6689(N22413,in0);
not not6690(N22414,R0);
not not6691(N22415,R1);
not not6692(N22425,in1);
not not6693(N22426,R2);
not not6694(N22427,R4);
not not6695(N22437,in1);
not not6696(N22438,R1);
not not6697(N22439,R4);
not not6698(N22449,in0);
not not6699(N22450,in2);
not not6700(N22451,R3);
not not6701(N22461,in0);
not not6702(N22462,in1);
not not6703(N22463,R5);
not not6704(N22473,in1);
not not6705(N22474,in2);
not not6706(N22475,R2);
not not6707(N22485,in2);
not not6708(N22486,R2);
not not6709(N22487,R3);
not not6710(N22497,in1);
not not6711(N22498,R2);
not not6712(N22499,R3);
not not6713(N22509,R0);
not not6714(N22510,R1);
not not6715(N22511,R3);
not not6716(N22512,R5);
not not6717(N22521,R0);
not not6718(N22522,R3);
not not6719(N22523,R4);
not not6720(N22533,in1);
not not6721(N22534,in2);
not not6722(N22535,R0);
not not6723(N22545,R0);
not not6724(N22546,R4);
not not6725(N22547,R5);
not not6726(N22557,in1);
not not6727(N22558,R1);
not not6728(N22559,R5);
not not6729(N22569,in2);
not not6730(N22570,R1);
not not6731(N22571,R4);
not not6732(N22581,in1);
not not6733(N22582,R4);
not not6734(N22583,R5);
not not6735(N22593,in1);
not not6736(N22594,in2);
not not6737(N22595,R3);
not not6738(N22605,in0);
not not6739(N22606,in2);
not not6740(N22607,R3);
not not6741(N22617,in2);
not not6742(N22618,R1);
not not6743(N22619,R3);
not not6744(N22629,in2);
not not6745(N22630,R1);
not not6746(N22631,R3);
not not6747(N22641,in1);
not not6748(N22642,R1);
not not6749(N22643,R5);
not not6750(N22653,in2);
not not6751(N22654,R2);
not not6752(N22665,in2);
not not6753(N22666,R2);
not not6754(N22667,R5);
not not6755(N22677,in0);
not not6756(N22678,in1);
not not6757(N22679,R2);
not not6758(N22689,in0);
not not6759(N22690,in1);
not not6760(N22691,R4);
not not6761(N22701,in1);
not not6762(N22702,R1);
not not6763(N22703,R4);
not not6764(N22704,R5);
not not6765(N22713,R0);
not not6766(N22714,R3);
not not6767(N22715,R4);
not not6768(N22725,R1);
not not6769(N22726,R2);
not not6770(N22727,R5);
not not6771(N22737,R0);
not not6772(N22738,R2);
not not6773(N22739,R4);
not not6774(N22749,in1);
not not6775(N22750,R0);
not not6776(N22751,R1);
not not6777(N22752,R5);
not not6778(N22761,in2);
not not6779(N22762,R0);
not not6780(N22763,R1);
not not6781(N22764,R5);
not not6782(N22773,in1);
not not6783(N22774,in2);
not not6784(N22775,R2);
not not6785(N22785,R0);
not not6786(N22786,R1);
not not6787(N22787,R4);
not not6788(N22788,R5);
not not6789(N22797,R0);
not not6790(N22798,R2);
not not6791(N22799,R5);
not not6792(N22809,R0);
not not6793(N22810,R1);
not not6794(N22811,R4);
not not6795(N22821,in1);
not not6796(N22822,in2);
not not6797(N22833,in1);
not not6798(N22844,in2);
not not6799(N22855,in0);
not not6800(N22856,R2);
not not6801(N22866,in0);
not not6802(N22867,R1);
not not6803(N22877,in1);
not not6804(N22878,R2);
not not6805(N22879,R5);
not not6806(N22888,R0);
not not6807(N22889,R1);
not not6808(N22899,R2);
not not6809(N22900,R3);
not not6810(N22901,R5);
not not6811(N22910,R3);
not not6812(N22911,R4);
not not6813(N22921,R3);
not not6814(N22922,R4);
not not6815(N22932,in2);
not not6816(N22933,R3);
not not6817(N22943,in1);
not not6818(N22944,R5);
not not6819(N22954,in2);
not not6820(N22955,R5);
not not6821(N22965,R3);
not not6822(N22966,R4);
not not6823(N22967,R5);
not not6824(N22976,R3);
not not6825(N22977,R4);
not not6826(N22978,R5);
not not6827(N22987,R0);
not not6828(N22988,R1);
not not6829(N22998,in1);
not not6830(N22999,R0);
not not6831(N23000,R4);
not not6832(N23009,in1);
not not6833(N23010,R3);
not not6834(N23020,R2);
not not6835(N23021,R3);
not not6836(N23031,R2);
not not6837(N23032,R3);
not not6838(N23042,in0);
not not6839(N23043,R2);
not not6840(N23044,R5);
not not6841(N23053,in2);
not not6842(N23054,R3);
not not6843(N23064,in1);
not not6844(N23065,R3);
not not6845(N23075,R0);
not not6846(N23076,R5);
not not6847(N23086,R0);
not not6848(N23087,R5);
not not6849(N23097,in1);
not not6850(N23098,in2);
not not6851(N23099,R2);
not not6852(N23108,R1);
not not6853(N23109,R5);
not not6854(N23119,R0);
not not6855(N23120,R3);
not not6856(N23130,in2);
not not6857(N23131,R3);
not not6858(N23141,in2);
not not6859(N23142,R4);
not not6860(N23152,R4);
not not6861(N23153,R5);
not not6862(N23163,in1);
not not6863(N23164,R0);
not not6864(N23165,R3);
not not6865(N23174,in1);
not not6866(N23175,R1);
not not6867(N23185,R2);
not not6868(N23196,in1);
not not6869(N23197,R4);
not not6870(N23207,in1);
not not6871(N23208,R4);
not not6872(N23218,R1);
not not6873(N23219,R3);
not not6874(N23229,R0);
not not6875(N23240,in1);
not not6876(N23241,R2);
not not6877(N23251,R5);
not not6878(N23262,in2);
not not6879(N23263,R2);
not not6880(N23264,R5);
not not6881(N23273,R1);
not not6882(N23274,R2);
not not6883(N23275,R5);
not not6884(N23284,in2);
not not6885(N23285,R0);
not not6886(N23286,R3);
not not6887(N23295,R0);
not not6888(N23296,R3);
not not6889(N23306,R1);
not not6890(N23307,R5);
not not6891(N23317,R1);
not not6892(N23318,R3);
not not6893(N23328,R2);
not not6894(N23329,R3);
not not6895(N23339,in1);
not not6896(N23340,R2);
not not6897(N23350,R0);
not not6898(N23351,R2);
not not6899(N23361,R2);
not not6900(N23362,R4);
not not6901(N23372,R0);
not not6902(N23373,R3);
not not6903(N23383,R3);
not not6904(N23384,R4);
not not6905(N23394,in2);
not not6906(N23395,R0);
not not6907(N23405,R0);
not not6908(N23415,in1);
not not6909(N23425,R2);
not not6910(N23435,in2);
not not6911(N23445,in1);
not not6912(N23455,in2);
not not6913(N23456,R4);
not not6914(N23465,in0);
not not6915(N23466,R4);
not not6916(N23475,in2);
not not6917(N23476,R3);
not not6918(N23485,in0);
not not6919(N23486,R3);
not not6920(N23495,in0);
not not6921(N23496,R3);
not not6922(N23505,in2);
not not6923(N23506,R0);
not not6924(N23515,in1);
not not6925(N23525,in1);
not not6926(N23526,R0);
not not6927(N23535,R0);
not not6928(N23536,R4);
not not6929(N23545,R2);
not not6930(N23555,R1);
not not6931(N23564,R1);
not not6932(N23573,in2);
not not6933(N23591,in1);
not not6934(N23618,in2);
not not6935(N23627,R4);
not not6936(N23643,R0);
not not6937(N23644,R2);
not not6938(N23645,R3);
not not6939(N23646,R4);
not not6940(N23647,R5);
not not6941(N23648,R6);
not not6942(N23649,R7);
not not6943(N23657,in0);
not not6944(N23658,in1);
not not6945(N23659,in2);
not not6946(N23660,R0);
not not6947(N23661,R5);
not not6948(N23662,R6);
not not6949(N23663,R7);
not not6950(N23671,R0);
not not6951(N23672,R1);
not not6952(N23673,R2);
not not6953(N23674,R4);
not not6954(N23675,R5);
not not6955(N23676,R6);
not not6956(N23684,R0);
not not6957(N23685,R1);
not not6958(N23686,R2);
not not6959(N23687,R3);
not not6960(N23688,R5);
not not6961(N23689,R6);
not not6962(N23697,in2);
not not6963(N23698,R0);
not not6964(N23699,R2);
not not6965(N23700,R4);
not not6966(N23701,R5);
not not6967(N23702,R7);
not not6968(N23710,in1);
not not6969(N23711,R2);
not not6970(N23712,R3);
not not6971(N23713,R4);
not not6972(N23714,R5);
not not6973(N23715,R6);
not not6974(N23723,R0);
not not6975(N23724,R1);
not not6976(N23725,R3);
not not6977(N23726,R4);
not not6978(N23727,R6);
not not6979(N23728,R7);
not not6980(N23736,in2);
not not6981(N23737,R0);
not not6982(N23738,R2);
not not6983(N23739,R5);
not not6984(N23740,R6);
not not6985(N23741,R7);
not not6986(N23749,R1);
not not6987(N23750,R4);
not not6988(N23751,R5);
not not6989(N23752,R6);
not not6990(N23753,R7);
not not6991(N23761,R0);
not not6992(N23762,R1);
not not6993(N23763,R3);
not not6994(N23764,R5);
not not6995(N23765,R7);
not not6996(N23773,in2);
not not6997(N23774,R1);
not not6998(N23775,R2);
not not6999(N23776,R4);
not not7000(N23777,R6);
not not7001(N23785,in1);
not not7002(N23786,R2);
not not7003(N23787,R5);
not not7004(N23788,R6);
not not7005(N23789,R7);
not not7006(N23797,in2);
not not7007(N23798,R1);
not not7008(N23799,R2);
not not7009(N23800,R4);
not not7010(N23801,R7);
not not7011(N23809,in1);
not not7012(N23810,R0);
not not7013(N23811,R4);
not not7014(N23812,R5);
not not7015(N23813,R6);
not not7016(N23821,in1);
not not7017(N23822,in2);
not not7018(N23823,R4);
not not7019(N23824,R6);
not not7020(N23825,R7);
not not7021(N23833,R1);
not not7022(N23834,R2);
not not7023(N23835,R3);
not not7024(N23836,R6);
not not7025(N23837,R7);
not not7026(N23845,R0);
not not7027(N23846,R2);
not not7028(N23847,R5);
not not7029(N23848,R6);
not not7030(N23849,R7);
not not7031(N23857,in0);
not not7032(N23858,in2);
not not7033(N23859,R4);
not not7034(N23860,R6);
not not7035(N23868,R2);
not not7036(N23869,R4);
not not7037(N23870,R5);
not not7038(N23871,R7);
not not7039(N23879,in2);
not not7040(N23880,R0);
not not7041(N23881,R1);
not not7042(N23882,R6);
not not7043(N23890,in2);
not not7044(N23891,R0);
not not7045(N23892,R4);
not not7046(N23893,R5);
not not7047(N23901,in1);
not not7048(N23902,R0);
not not7049(N23903,R4);
not not7050(N23904,R5);
not not7051(N23912,R2);
not not7052(N23913,R4);
not not7053(N23914,R5);
not not7054(N23915,R7);
not not7055(N23923,R1);
not not7056(N23924,R2);
not not7057(N23925,R4);
not not7058(N23926,R7);
not not7059(N23934,in1);
not not7060(N23935,R4);
not not7061(N23936,R6);
not not7062(N23937,R7);
not not7063(N23945,R2);
not not7064(N23946,R4);
not not7065(N23947,R6);
not not7066(N23955,in1);
not not7067(N23956,R1);
not not7068(N23957,R7);
not not7069(N23965,in2);
not not7070(N23966,R1);
not not7071(N23967,R6);
not not7072(N23975,R0);
not not7073(N23976,R5);
not not7074(N23977,R6);
not not7075(N23985,R1);
not not7076(N23986,R3);
not not7077(N23987,R5);
not not7078(N23995,R2);
not not7079(N23996,R3);
not not7080(N23997,R5);
not not7081(N24005,R1);
not not7082(N24006,R4);
not not7083(N24007,R6);
not not7084(N24015,R1);
not not7085(N24016,R3);
not not7086(N24017,R6);
not not7087(N24025,in1);
not not7088(N24026,R2);
not not7089(N24027,R4);
not not7090(N24035,in2);
not not7091(N24036,R1);
not not7092(N24037,R6);
not not7093(N24045,in1);
not not7094(N24046,R1);
not not7095(N24054,R3);
not not7096(N24055,R5);
not not7097(N18124,R4);
not not7098(N18125,R5);
not not7099(N18126,R6);
not not7100(N18127,R7);
not not7101(N18142,R4);
not not7102(N18143,R6);
not not7103(N18144,R7);
not not7104(N18159,R4);
not not7105(N18160,R5);
not not7106(N18161,R6);
not not7107(N18176,R4);
not not7108(N18177,R5);
not not7109(N18178,R6);
not not7110(N18193,R4);
not not7111(N18194,R5);
not not7112(N18195,R7);
not not7113(N18211,R6);
not not7114(N18212,R7);
not not7115(N18227,R3);
not not7116(N18228,R5);
not not7117(N18229,R6);
not not7118(N18242,R4);
not not7119(N18243,R5);
not not7120(N18244,R6);
not not7121(N18245,R7);
not not7122(N18260,R6);
not not7123(N18261,R7);
not not7124(N18275,R5);
not not7125(N18276,R6);
not not7126(N18277,R7);
not not7127(N18291,R5);
not not7128(N18292,R6);
not not7129(N18293,R7);
not not7130(N18307,R5);
not not7131(N18308,R6);
not not7132(N18309,R7);
not not7133(N18323,R4);
not not7134(N18324,R5);
not not7135(N18325,R6);
not not7136(N18339,R5);
not not7137(N18340,R6);
not not7138(N18341,R7);
not not7139(N18355,R3);
not not7140(N18356,R5);
not not7141(N18357,R6);
not not7142(N18372,R4);
not not7143(N18373,R5);
not not7144(N18387,R4);
not not7145(N18388,R5);
not not7146(N18389,R7);
not not7147(N18402,R4);
not not7148(N18403,R5);
not not7149(N18404,R6);
not not7150(N18405,R7);
not not7151(N18418,R4);
not not7152(N18419,R5);
not not7153(N18420,R6);
not not7154(N18421,R7);
not not7155(N18435,R5);
not not7156(N18436,R6);
not not7157(N18437,R7);
not not7158(N18451,R4);
not not7159(N18452,R6);
not not7160(N18453,R7);
not not7161(N18467,R4);
not not7162(N18468,R6);
not not7163(N18469,R7);
not not7164(N18483,R4);
not not7165(N18484,R5);
not not7166(N18485,R6);
not not7167(N18499,R3);
not not7168(N18500,R5);
not not7169(N18501,R7);
not not7170(N18515,R3);
not not7171(N18516,R4);
not not7172(N18517,R5);
not not7173(N18531,R3);
not not7174(N18532,R4);
not not7175(N18533,R5);
not not7176(N18548,R5);
not not7177(N18549,R6);
not not7178(N18563,R4);
not not7179(N18564,R7);
not not7180(N18576,R4);
not not7181(N18577,R5);
not not7182(N18578,R6);
not not7183(N18579,R7);
not not7184(N18592,R4);
not not7185(N18593,R5);
not not7186(N18594,R7);
not not7187(N18606,R4);
not not7188(N18607,R5);
not not7189(N18608,R6);
not not7190(N18609,R7);
not not7191(N18623,R4);
not not7192(N18624,R7);
not not7193(N18637,R4);
not not7194(N18638,R5);
not not7195(N18639,R7);
not not7196(N18652,R4);
not not7197(N18653,R6);
not not7198(N18654,R7);
not not7199(N18667,R4);
not not7200(N18668,R6);
not not7201(N18669,R7);
not not7202(N18683,R4);
not not7203(N18684,R7);
not not7204(N18697,R3);
not not7205(N18698,R6);
not not7206(N18699,R7);
not not7207(N18713,R4);
not not7208(N18714,R7);
not not7209(N18728,R4);
not not7210(N18729,R5);
not not7211(N18741,R4);
not not7212(N18742,R5);
not not7213(N18743,R6);
not not7214(N18744,R7);
not not7215(N18756,R4);
not not7216(N18757,R5);
not not7217(N18758,R6);
not not7218(N18759,R7);
not not7219(N18771,R3);
not not7220(N18772,R5);
not not7221(N18773,R6);
not not7222(N18774,R7);
not not7223(N18788,R5);
not not7224(N18789,R6);
not not7225(N18803,R5);
not not7226(N18804,R6);
not not7227(N18818,R4);
not not7228(N18819,R7);
not not7229(N18832,R4);
not not7230(N18833,R6);
not not7231(N18834,R7);
not not7232(N18847,R4);
not not7233(N18848,R5);
not not7234(N18849,R6);
not not7235(N18863,R6);
not not7236(N18864,R7);
not not7237(N18877,R4);
not not7238(N18878,R5);
not not7239(N18879,R7);
not not7240(N18892,R3);
not not7241(N18893,R4);
not not7242(N18894,R6);
not not7243(N18908,R6);
not not7244(N18909,R7);
not not7245(N18921,R5);
not not7246(N18922,R6);
not not7247(N18923,R7);
not not7248(N18935,R5);
not not7249(N18936,R6);
not not7250(N18937,R7);
not not7251(N18949,R4);
not not7252(N18950,R5);
not not7253(N18951,R7);
not not7254(N18963,R4);
not not7255(N18964,R6);
not not7256(N18965,R7);
not not7257(N18977,R5);
not not7258(N18978,R6);
not not7259(N18979,R7);
not not7260(N18992,R6);
not not7261(N18993,R7);
not not7262(N19006,R6);
not not7263(N19007,R7);
not not7264(N19019,R4);
not not7265(N19020,R6);
not not7266(N19021,R7);
not not7267(N19034,R4);
not not7268(N19035,R7);
not not7269(N19048,R5);
not not7270(N19049,R6);
not not7271(N19062,R5);
not not7272(N19063,R6);
not not7273(N19076,R6);
not not7274(N19077,R7);
not not7275(N19090,R6);
not not7276(N19091,R7);
not not7277(N19105,R5);
not not7278(N19118,R4);
not not7279(N19119,R7);
not not7280(N19132,R6);
not not7281(N19133,R7);
not not7282(N19146,R4);
not not7283(N19147,R6);
not not7284(N19161,R6);
not not7285(N19173,R4);
not not7286(N19174,R6);
not not7287(N19175,R7);
not not7288(N19187,R4);
not not7289(N19188,R6);
not not7290(N19189,R7);
not not7291(N19201,R5);
not not7292(N19202,R6);
not not7293(N19203,R7);
not not7294(N19217,R7);
not not7295(N19230,R4);
not not7296(N19231,R5);
not not7297(N19244,R4);
not not7298(N19245,R5);
not not7299(N19258,R4);
not not7300(N19259,R5);
not not7301(N19272,R4);
not not7302(N19273,R6);
not not7303(N19286,R4);
not not7304(N19287,R6);
not not7305(N19300,R4);
not not7306(N19301,R6);
not not7307(N19315,R6);
not not7308(N19328,R4);
not not7309(N19329,R6);
not not7310(N19342,R5);
not not7311(N19343,R6);
not not7312(N19356,R5);
not not7313(N19357,R7);
not not7314(N19369,R5);
not not7315(N19370,R6);
not not7316(N19371,R7);
not not7317(N19384,R4);
not not7318(N19385,R6);
not not7319(N19398,R5);
not not7320(N19399,R7);
not not7321(N19413,R7);
not not7322(N19427,R5);
not not7323(N19441,R5);
not not7324(N19453,R3);
not not7325(N19454,R5);
not not7326(N19455,R6);
not not7327(N19467,R4);
not not7328(N19468,R5);
not not7329(N19469,R6);
not not7330(N19482,R4);
not not7331(N19483,R7);
not not7332(N19495,R4);
not not7333(N19496,R6);
not not7334(N19497,R7);
not not7335(N19510,R5);
not not7336(N19511,R6);
not not7337(N19524,R5);
not not7338(N19525,R6);
not not7339(N19538,R3);
not not7340(N19539,R6);
not not7341(N19552,R5);
not not7342(N19553,R7);
not not7343(N19567,R7);
not not7344(N19580,R6);
not not7345(N19581,R7);
not not7346(N19593,R3);
not not7347(N19594,R4);
not not7348(N19595,R7);
not not7349(N19608,R4);
not not7350(N19609,R5);
not not7351(N19623,R4);
not not7352(N19636,R3);
not not7353(N19637,R5);
not not7354(N19649,R3);
not not7355(N19650,R4);
not not7356(N19651,R7);
not not7357(N19663,R4);
not not7358(N19664,R6);
not not7359(N19665,R7);
not not7360(N19679,R6);
not not7361(N19692,R5);
not not7362(N19693,R6);
not not7363(N19706,R5);
not not7364(N19707,R6);
not not7365(N19720,R5);
not not7366(N19721,R6);
not not7367(N19733,R4);
not not7368(N19734,R5);
not not7369(N19745,R5);
not not7370(N19746,R6);
not not7371(N19747,R7);
not not7372(N19759,R5);
not not7373(N19760,R6);
not not7374(N19785,R4);
not not7375(N19786,R6);
not not7376(N19798,R5);
not not7377(N19799,R6);
not not7378(N19810,R4);
not not7379(N19811,R5);
not not7380(N19812,R7);
not not7381(N19824,R4);
not not7382(N19825,R7);
not not7383(N19837,R4);
not not7384(N19838,R5);
not not7385(N19851,R7);
not not7386(N19862,R4);
not not7387(N19863,R5);
not not7388(N19864,R7);
not not7389(N19877,R7);
not not7390(N19890,R6);
not not7391(N19903,R6);
not not7392(N19915,R6);
not not7393(N19916,R7);
not not7394(N19928,R6);
not not7395(N19929,R7);
not not7396(N19941,R4);
not not7397(N19942,R7);
not not7398(N19955,R7);
not not7399(N19968,R4);
not not7400(N19981,R7);
not not7401(N19993,R5);
not not7402(N19994,R7);
not not7403(N20007,R5);
not not7404(N20020,R5);
not not7405(N20032,R6);
not not7406(N20033,R7);
not not7407(N20045,R5);
not not7408(N20046,R7);
not not7409(N20058,R5);
not not7410(N20059,R7);
not not7411(N20071,R5);
not not7412(N20072,R7);
not not7413(N20084,R5);
not not7414(N20085,R7);
not not7415(N20098,R4);
not not7416(N20110,R4);
not not7417(N20111,R5);
not not7418(N20124,R6);
not not7419(N20137,R6);
not not7420(N20149,R6);
not not7421(N20150,R7);
not not7422(N20163,R5);
not not7423(N20176,R7);
not not7424(N20188,R6);
not not7425(N20189,R7);
not not7426(N20201,R6);
not not7427(N20202,R7);
not not7428(N20214,R6);
not not7429(N20215,R7);
not not7430(N20228,R3);
not not7431(N20240,R5);
not not7432(N20241,R6);
not not7433(N20252,R4);
not not7434(N20253,R7);
not not7435(N20264,R6);
not not7436(N20265,R7);
not not7437(N20277,R6);
not not7438(N20289,R6);
not not7439(N20300,R5);
not not7440(N20301,R6);
not not7441(N20313,R5);
not not7442(N20324,R5);
not not7443(N20325,R7);
not not7444(N20336,R4);
not not7445(N20337,R6);
not not7446(N20349,R7);
not not7447(N20360,R4);
not not7448(N20361,R5);
not not7449(N20373,R6);
not not7450(N20384,R6);
not not7451(N20385,R7);
not not7452(N20395,R4);
not not7453(N20396,R5);
not not7454(N20397,R7);
not not7455(N20408,R4);
not not7456(N20409,R7);
not not7457(N20421,R4);
not not7458(N20433,R4);
not not7459(N20444,R6);
not not7460(N20445,R7);
not not7461(N20455,R4);
not not7462(N20456,R6);
not not7463(N20457,R7);
not not7464(N20468,R4);
not not7465(N20469,R7);
not not7466(N20481,R4);
not not7467(N20504,R4);
not not7468(N20505,R5);
not not7469(N20516,R5);
not not7470(N20517,R6);
not not7471(N20541,R5);
not not7472(N20553,R5);
not not7473(N20565,R6);
not not7474(N20589,R7);
not not7475(N20601,R6);
not not7476(N20613,R5);
not not7477(N20624,R6);
not not7478(N20625,R7);
not not7479(N20636,R4);
not not7480(N20637,R5);
not not7481(N20648,R6);
not not7482(N20649,R7);
not not7483(N20660,R5);
not not7484(N20661,R6);
not not7485(N20671,R4);
not not7486(N20672,R5);
not not7487(N20683,R7);
not not7488(N20694,R5);
not not7489(N20705,R5);
not not7490(N20727,R3);
not not7491(N20737,R3);
not not7492(N20767,R4);
not not7493(N20787,R7);
not not7494(N20797,R6);
not not7495(N20807,R7);
not not7496(N20817,R6);
not not7497(N20837,R5);
not not7498(N20862,R6);
not not7499(N20863,R7);
not not7500(N20878,R5);
not not7501(N20879,R6);
not not7502(N20893,R6);
not not7503(N20894,R7);
not not7504(N20909,R7);
not not7505(N20923,R6);
not not7506(N20924,R7);
not not7507(N20939,R7);
not not7508(N20954,R7);
not not7509(N20968,R6);
not not7510(N20969,R7);
not not7511(N20983,R6);
not not7512(N20984,R7);
not not7513(N20998,R5);
not not7514(N20999,R7);
not not7515(N21013,R5);
not not7516(N21014,R6);
not not7517(N21028,R6);
not not7518(N21029,R7);
not not7519(N21043,R6);
not not7520(N21044,R7);
not not7521(N21059,R7);
not not7522(N21073,R5);
not not7523(N21074,R6);
not not7524(N21087,R6);
not not7525(N21088,R7);
not not7526(N21101,R6);
not not7527(N21102,R7);
not not7528(N21115,R6);
not not7529(N21116,R7);
not not7530(N21129,R6);
not not7531(N21130,R7);
not not7532(N21144,R6);
not not7533(N21158,R6);
not not7534(N21171,R5);
not not7535(N21172,R7);
not not7536(N21185,R6);
not not7537(N21186,R7);
not not7538(N21200,R7);
not not7539(N21214,R7);
not not7540(N21228,R6);
not not7541(N21242,R6);
not not7542(N21256,R7);
not not7543(N21269,R6);
not not7544(N21270,R7);
not not7545(N21283,R6);
not not7546(N21284,R7);
not not7547(N21297,R6);
not not7548(N21298,R7);
not not7549(N21311,R6);
not not7550(N21312,R7);
not not7551(N21326,R6);
not not7552(N21340,R7);
not not7553(N21353,R5);
not not7554(N21354,R6);
not not7555(N21367,R5);
not not7556(N21368,R6);
not not7557(N21381,R6);
not not7558(N21382,R7);
not not7559(N21396,R6);
not not7560(N21409,R6);
not not7561(N21410,R7);
not not7562(N21424,R7);
not not7563(N21438,R6);
not not7564(N21452,R7);
not not7565(N21465,R6);
not not7566(N21466,R7);
not not7567(N21479,R6);
not not7568(N21480,R7);
not not7569(N21493,R6);
not not7570(N21494,R7);
not not7571(N21508,R7);
not not7572(N21521,R6);
not not7573(N21522,R7);
not not7574(N21534,R6);
not not7575(N21535,R7);
not not7576(N21548,R6);
not not7577(N21560,R6);
not not7578(N21561,R7);
not not7579(N21574,R7);
not not7580(N21586,R6);
not not7581(N21587,R7);
not not7582(N21600,R7);
not not7583(N21613,R7);
not not7584(N21626,R7);
not not7585(N21639,R5);
not not7586(N21652,R6);
not not7587(N21664,R5);
not not7588(N21665,R6);
not not7589(N21677,R6);
not not7590(N21678,R7);
not not7591(N21730,R6);
not not7592(N21743,R6);
not not7593(N21756,R7);
not not7594(N21769,R7);
not not7595(N21782,R7);
not not7596(N21795,R7);
not not7597(N21807,R6);
not not7598(N21808,R7);
not not7599(N21821,R7);
not not7600(N21834,R7);
not not7601(N21860,R7);
not not7602(N21872,R6);
not not7603(N21873,R7);
not not7604(N21886,R6);
not not7605(N21899,R6);
not not7606(N21912,R6);
not not7607(N21925,R6);
not not7608(N21964,R5);
not not7609(N21977,R5);
not not7610(N21990,R5);
not not7611(N22003,R5);
not not7612(N22016,R6);
not not7613(N22029,R5);
not not7614(N22042,R6);
not not7615(N22055,R6);
not not7616(N22067,R6);
not not7617(N22068,R7);
not not7618(N22081,R6);
not not7619(N22094,R6);
not not7620(N22106,R6);
not not7621(N22107,R7);
not not7622(N22120,R6);
not not7623(N22132,R6);
not not7624(N22133,R7);
not not7625(N22146,R5);
not not7626(N22159,R6);
not not7627(N22171,R5);
not not7628(N22172,R6);
not not7629(N22185,R7);
not not7630(N22198,R6);
not not7631(N22211,R5);
not not7632(N22223,R6);
not not7633(N22224,R7);
not not7634(N22236,R6);
not not7635(N22247,R5);
not not7636(N22248,R7);
not not7637(N22259,R6);
not not7638(N22260,R7);
not not7639(N22284,R7);
not not7640(N22296,R7);
not not7641(N22307,R6);
not not7642(N22308,R7);
not not7643(N22319,R6);
not not7644(N22320,R7);
not not7645(N22332,R5);
not not7646(N22344,R7);
not not7647(N22356,R5);
not not7648(N22368,R6);
not not7649(N22380,R7);
not not7650(N22392,R7);
not not7651(N22416,R6);
not not7652(N22428,R7);
not not7653(N22440,R6);
not not7654(N22452,R7);
not not7655(N22464,R6);
not not7656(N22476,R6);
not not7657(N22488,R6);
not not7658(N22500,R6);
not not7659(N22524,R5);
not not7660(N22536,R7);
not not7661(N22548,R6);
not not7662(N22560,R6);
not not7663(N22572,R6);
not not7664(N22584,R6);
not not7665(N22596,R7);
not not7666(N22608,R7);
not not7667(N22620,R7);
not not7668(N22632,R7);
not not7669(N22644,R7);
not not7670(N22655,R6);
not not7671(N22656,R7);
not not7672(N22668,R6);
not not7673(N22680,R6);
not not7674(N22692,R6);
not not7675(N22716,R6);
not not7676(N22728,R7);
not not7677(N22740,R7);
not not7678(N22776,R7);
not not7679(N22800,R7);
not not7680(N22812,R6);
not not7681(N22823,R6);
not not7682(N22824,R7);
not not7683(N22834,R5);
not not7684(N22835,R7);
not not7685(N22845,R5);
not not7686(N22846,R7);
not not7687(N22857,R7);
not not7688(N22868,R7);
not not7689(N22890,R7);
not not7690(N22912,R6);
not not7691(N22923,R7);
not not7692(N22934,R7);
not not7693(N22945,R7);
not not7694(N22956,R7);
not not7695(N22989,R6);
not not7696(N23011,R7);
not not7697(N23022,R7);
not not7698(N23033,R7);
not not7699(N23055,R6);
not not7700(N23066,R6);
not not7701(N23077,R6);
not not7702(N23088,R6);
not not7703(N23110,R6);
not not7704(N23121,R6);
not not7705(N23132,R6);
not not7706(N23143,R6);
not not7707(N23154,R6);
not not7708(N23176,R6);
not not7709(N23186,R6);
not not7710(N23187,R7);
not not7711(N23198,R7);
not not7712(N23209,R7);
not not7713(N23220,R6);
not not7714(N23230,R6);
not not7715(N23231,R7);
not not7716(N23242,R5);
not not7717(N23252,R6);
not not7718(N23253,R7);
not not7719(N23297,R7);
not not7720(N23308,R7);
not not7721(N23319,R7);
not not7722(N23330,R6);
not not7723(N23341,R6);
not not7724(N23352,R7);
not not7725(N23363,R7);
not not7726(N23374,R5);
not not7727(N23385,R6);
not not7728(N23396,R7);
not not7729(N23406,R6);
not not7730(N23416,R6);
not not7731(N23426,R6);
not not7732(N23436,R5);
not not7733(N23446,R5);
not not7734(N23516,R7);
not not7735(N23546,R4);
not not7736(N23582,R7);
not not7737(N23600,R7);
not not7738(N23609,R5);
not not7739(N24436,in0);
not not7740(N24437,in1);
not not7741(N24438,in2);
not not7742(N24439,R0);
not not7743(N24440,R1);
not not7744(N24453,in0);
not not7745(N24454,R0);
not not7746(N24455,R1);
not not7747(N24456,R2);
not not7748(N24470,in0);
not not7749(N24471,in1);
not not7750(N24472,R0);
not not7751(N24473,R1);
not not7752(N24474,R2);
not not7753(N24487,in0);
not not7754(N24488,in2);
not not7755(N24489,R0);
not not7756(N24490,R3);
not not7757(N24504,in0);
not not7758(N24505,in1);
not not7759(N24506,R0);
not not7760(N24507,R1);
not not7761(N24521,in0);
not not7762(N24522,in1);
not not7763(N24523,in2);
not not7764(N24524,R1);
not not7765(N24525,R3);
not not7766(N24538,in0);
not not7767(N24539,in1);
not not7768(N24540,in2);
not not7769(N24541,R0);
not not7770(N24542,R2);
not not7771(N24555,in0);
not not7772(N24556,in1);
not not7773(N24557,in2);
not not7774(N24558,R0);
not not7775(N24559,R2);
not not7776(N24572,in0);
not not7777(N24573,in1);
not not7778(N24574,R0);
not not7779(N24575,R2);
not not7780(N24588,in1);
not not7781(N24589,R0);
not not7782(N24590,R1);
not not7783(N24591,R2);
not not7784(N24604,R0);
not not7785(N24605,R1);
not not7786(N24606,R2);
not not7787(N24607,R3);
not not7788(N24620,in1);
not not7789(N24621,R0);
not not7790(N24622,R1);
not not7791(N24623,R2);
not not7792(N24636,in0);
not not7793(N24637,in2);
not not7794(N24638,R1);
not not7795(N24639,R3);
not not7796(N24652,in0);
not not7797(N24653,in2);
not not7798(N24654,R3);
not not7799(N24668,in0);
not not7800(N24669,in1);
not not7801(N24670,R2);
not not7802(N24671,R3);
not not7803(N24684,in0);
not not7804(N24685,in1);
not not7805(N24686,in2);
not not7806(N24687,R0);
not not7807(N24688,R1);
not not7808(N24700,in0);
not not7809(N24701,in1);
not not7810(N24702,R0);
not not7811(N24703,R1);
not not7812(N24704,R3);
not not7813(N24716,in0);
not not7814(N24717,in1);
not not7815(N24718,R0);
not not7816(N24719,R2);
not not7817(N24720,R3);
not not7818(N24732,in0);
not not7819(N24733,in1);
not not7820(N24734,R0);
not not7821(N24735,R2);
not not7822(N24748,in0);
not not7823(N24749,in1);
not not7824(N24750,R2);
not not7825(N24751,R3);
not not7826(N24764,in0);
not not7827(N24765,in1);
not not7828(N24766,R1);
not not7829(N24767,R2);
not not7830(N24780,in0);
not not7831(N24781,in1);
not not7832(N24782,in2);
not not7833(N24783,R0);
not not7834(N24796,in0);
not not7835(N24797,R0);
not not7836(N24798,R1);
not not7837(N24812,in0);
not not7838(N24813,in2);
not not7839(N24814,R0);
not not7840(N24815,R3);
not not7841(N24828,in0);
not not7842(N24829,in1);
not not7843(N24830,R0);
not not7844(N24831,R3);
not not7845(N24844,in0);
not not7846(N24845,R1);
not not7847(N24846,R2);
not not7848(N24860,in0);
not not7849(N24861,in1);
not not7850(N24862,R0);
not not7851(N24863,R3);
not not7852(N24876,in1);
not not7853(N24877,R1);
not not7854(N24891,in1);
not not7855(N24892,in2);
not not7856(N24893,R0);
not not7857(N24894,R2);
not not7858(N24906,in0);
not not7859(N24907,R0);
not not7860(N24908,R1);
not not7861(N24921,in0);
not not7862(N24922,in1);
not not7863(N24923,R1);
not not7864(N24936,in0);
not not7865(N24937,in2);
not not7866(N24938,R1);
not not7867(N24939,R2);
not not7868(N24951,in0);
not not7869(N24952,in2);
not not7870(N24953,R0);
not not7871(N24954,R2);
not not7872(N24966,in0);
not not7873(N24967,in1);
not not7874(N24968,R2);
not not7875(N24969,R3);
not not7876(N24981,in0);
not not7877(N24982,in1);
not not7878(N24983,in2);
not not7879(N24984,R0);
not not7880(N24985,R2);
not not7881(N24996,in1);
not not7882(N24997,in2);
not not7883(N24998,R0);
not not7884(N24999,R3);
not not7885(N25011,in2);
not not7886(N25012,R0);
not not7887(N25013,R1);
not not7888(N25014,R3);
not not7889(N25026,in1);
not not7890(N25027,R0);
not not7891(N25028,R1);
not not7892(N25041,in0);
not not7893(N25042,R0);
not not7894(N25043,R1);
not not7895(N25056,in1);
not not7896(N25057,in2);
not not7897(N25058,R1);
not not7898(N25059,R3);
not not7899(N25071,in0);
not not7900(N25072,in1);
not not7901(N25073,in2);
not not7902(N25074,R1);
not not7903(N25086,R0);
not not7904(N25087,R1);
not not7905(N25088,R2);
not not7906(N25089,R3);
not not7907(N25101,in0);
not not7908(N25102,R0);
not not7909(N25103,R2);
not not7910(N25104,R3);
not not7911(N25116,in0);
not not7912(N25117,in2);
not not7913(N25118,R2);
not not7914(N25119,R3);
not not7915(N25131,in1);
not not7916(N25132,R0);
not not7917(N25133,R1);
not not7918(N25134,R2);
not not7919(N25146,in0);
not not7920(N25147,R0);
not not7921(N25148,R2);
not not7922(N25161,in0);
not not7923(N25162,in2);
not not7924(N25163,R0);
not not7925(N25164,R2);
not not7926(N25176,in0);
not not7927(N25177,in1);
not not7928(N25178,in2);
not not7929(N25179,R0);
not not7930(N25180,R3);
not not7931(N25191,in0);
not not7932(N25192,in1);
not not7933(N25193,in2);
not not7934(N25194,R0);
not not7935(N25195,R1);
not not7936(N25206,in0);
not not7937(N25207,in2);
not not7938(N25208,R0);
not not7939(N25209,R1);
not not7940(N25221,in0);
not not7941(N25222,R1);
not not7942(N25223,R3);
not not7943(N25236,in0);
not not7944(N25237,in2);
not not7945(N25238,R1);
not not7946(N25251,in0);
not not7947(N25252,in1);
not not7948(N25253,in2);
not not7949(N25254,R2);
not not7950(N25266,in1);
not not7951(N25267,in2);
not not7952(N25268,R2);
not not7953(N25280,R0);
not not7954(N25281,R2);
not not7955(N25294,in0);
not not7956(N25295,in2);
not not7957(N25296,R1);
not not7958(N25308,in0);
not not7959(N25309,R0);
not not7960(N25310,R2);
not not7961(N25322,in1);
not not7962(N25323,R0);
not not7963(N25324,R3);
not not7964(N25336,in0);
not not7965(N25337,in2);
not not7966(N25338,R0);
not not7967(N25350,in0);
not not7968(N25351,in2);
not not7969(N25352,R3);
not not7970(N25364,in1);
not not7971(N25365,R0);
not not7972(N25366,R3);
not not7973(N25378,in0);
not not7974(N25379,R1);
not not7975(N25392,in1);
not not7976(N25393,R2);
not not7977(N25406,in0);
not not7978(N25407,R2);
not not7979(N25420,in2);
not not7980(N25421,R0);
not not7981(N25422,R2);
not not7982(N25434,in0);
not not7983(N25435,R0);
not not7984(N25436,R2);
not not7985(N25448,in1);
not not7986(N25449,R0);
not not7987(N25450,R2);
not not7988(N25451,R3);
not not7989(N25462,R0);
not not7990(N25463,R1);
not not7991(N25464,R3);
not not7992(N25476,in0);
not not7993(N25477,in1);
not not7994(N25478,in2);
not not7995(N25479,R1);
not not7996(N25490,in0);
not not7997(N25491,in1);
not not7998(N25492,in2);
not not7999(N25493,R0);
not not8000(N25504,in1);
not not8001(N25505,in2);
not not8002(N25506,R1);
not not8003(N25507,R2);
not not8004(N25518,in0);
not not8005(N25519,R0);
not not8006(N25532,in0);
not not8007(N25533,in1);
not not8008(N25534,R3);
not not8009(N25546,in0);
not not8010(N25547,in2);
not not8011(N25548,R3);
not not8012(N25560,R2);
not not8013(N25561,R3);
not not8014(N25574,in0);
not not8015(N25575,in1);
not not8016(N25576,R1);
not not8017(N25577,R2);
not not8018(N25588,R1);
not not8019(N25589,R2);
not not8020(N25602,R0);
not not8021(N25603,R1);
not not8022(N25616,in2);
not not8023(N25617,R0);
not not8024(N25618,R1);
not not8025(N25630,in0);
not not8026(N25631,in1);
not not8027(N25632,in2);
not not8028(N25633,R2);
not not8029(N25644,in0);
not not8030(N25645,R0);
not not8031(N25658,in2);
not not8032(N25659,R2);
not not8033(N25660,R3);
not not8034(N25672,in0);
not not8035(N25673,in1);
not not8036(N25686,R0);
not not8037(N25687,R1);
not not8038(N25688,R2);
not not8039(N25700,in2);
not not8040(N25701,R1);
not not8041(N25702,R2);
not not8042(N25714,in0);
not not8043(N25715,in1);
not not8044(N25716,R0);
not not8045(N25728,in2);
not not8046(N25729,R0);
not not8047(N25730,R2);
not not8048(N25742,in0);
not not8049(N25743,in2);
not not8050(N25744,R0);
not not8051(N25745,R1);
not not8052(N25756,in0);
not not8053(N25757,in1);
not not8054(N25758,R0);
not not8055(N25759,R1);
not not8056(N25770,R0);
not not8057(N25771,R1);
not not8058(N25772,R3);
not not8059(N25784,in0);
not not8060(N25785,R0);
not not8061(N25786,R3);
not not8062(N25798,R0);
not not8063(N25799,R3);
not not8064(N25812,in0);
not not8065(N25813,in2);
not not8066(N25814,R0);
not not8067(N25815,R1);
not not8068(N25826,in1);
not not8069(N25827,in2);
not not8070(N25828,R1);
not not8071(N25840,in2);
not not8072(N25841,R0);
not not8073(N25854,in0);
not not8074(N25855,R2);
not not8075(N25868,in0);
not not8076(N25869,in1);
not not8077(N25870,in2);
not not8078(N25871,R2);
not not8079(N25882,R0);
not not8080(N25883,R2);
not not8081(N25884,R3);
not not8082(N25896,in0);
not not8083(N25897,R0);
not not8084(N25898,R2);
not not8085(N25899,R3);
not not8086(N25910,in0);
not not8087(N25911,in1);
not not8088(N25912,R0);
not not8089(N25913,R1);
not not8090(N25924,in0);
not not8091(N25925,R0);
not not8092(N25926,R1);
not not8093(N25927,R3);
not not8094(N25938,in0);
not not8095(N25939,in1);
not not8096(N25940,R1);
not not8097(N25952,in0);
not not8098(N25953,in1);
not not8099(N25954,R1);
not not8100(N25966,in0);
not not8101(N25967,R1);
not not8102(N25980,in0);
not not8103(N25981,R2);
not not8104(N25994,in0);
not not8105(N25995,R2);
not not8106(N26008,in0);
not not8107(N26009,in2);
not not8108(N26022,in0);
not not8109(N26023,R1);
not not8110(N26024,R2);
not not8111(N26036,in0);
not not8112(N26037,in1);
not not8113(N26038,R1);
not not8114(N26039,R2);
not not8115(N26050,in0);
not not8116(N26051,in1);
not not8117(N26052,in2);
not not8118(N26064,in0);
not not8119(N26065,in2);
not not8120(N26078,in0);
not not8121(N26079,R0);
not not8122(N26092,in2);
not not8123(N26093,R0);
not not8124(N26106,in1);
not not8125(N26107,in2);
not not8126(N26108,R1);
not not8127(N26120,in1);
not not8128(N26121,R0);
not not8129(N26122,R1);
not not8130(N26134,in2);
not not8131(N26135,R0);
not not8132(N26136,R1);
not not8133(N26148,in0);
not not8134(N26161,in2);
not not8135(N26162,R2);
not not8136(N26174,in2);
not not8137(N26175,R1);
not not8138(N26187,in0);
not not8139(N26188,in1);
not not8140(N26189,R1);
not not8141(N26200,R0);
not not8142(N26201,R3);
not not8143(N26213,in2);
not not8144(N26214,R1);
not not8145(N26226,in0);
not not8146(N26227,in1);
not not8147(N26228,R3);
not not8148(N26239,R0);
not not8149(N26240,R3);
not not8150(N26252,in1);
not not8151(N26253,R1);
not not8152(N26265,R0);
not not8153(N26266,R2);
not not8154(N26267,R3);
not not8155(N26278,R1);
not not8156(N26279,R3);
not not8157(N26291,in0);
not not8158(N26292,R0);
not not8159(N26293,R1);
not not8160(N26304,in1);
not not8161(N26317,in0);
not not8162(N26318,in2);
not not8163(N26319,R2);
not not8164(N26330,in0);
not not8165(N26331,R2);
not not8166(N26332,R3);
not not8167(N26343,in0);
not not8168(N26344,in1);
not not8169(N26345,R1);
not not8170(N26356,in0);
not not8171(N26357,in2);
not not8172(N26358,R1);
not not8173(N26369,in1);
not not8174(N26370,in2);
not not8175(N26371,R2);
not not8176(N26382,in1);
not not8177(N26383,R2);
not not8178(N26395,in0);
not not8179(N26396,in1);
not not8180(N26397,in2);
not not8181(N26408,in2);
not not8182(N26409,R0);
not not8183(N26421,R0);
not not8184(N26422,R2);
not not8185(N26434,in1);
not not8186(N26435,in2);
not not8187(N26436,R0);
not not8188(N26447,in0);
not not8189(N26448,in2);
not not8190(N26449,R0);
not not8191(N26460,in0);
not not8192(N26473,in1);
not not8193(N26474,R3);
not not8194(N26486,R3);
not not8195(N26499,in0);
not not8196(N26500,R0);
not not8197(N26501,R1);
not not8198(N26512,in0);
not not8199(N26513,R2);
not not8200(N26524,R2);
not not8201(N26536,in1);
not not8202(N26537,R2);
not not8203(N26548,in1);
not not8204(N26549,R0);
not not8205(N26560,in0);
not not8206(N26572,in0);
not not8207(N26573,R3);
not not8208(N26584,in0);
not not8209(N26596,R0);
not not8210(N26608,R2);
not not8211(N26620,in2);
not not8212(N26621,R0);
not not8213(N26632,in0);
not not8214(N26633,R1);
not not8215(N26644,R1);
not not8216(N26645,R2);
not not8217(N26656,in2);
not not8218(N26657,R2);
not not8219(N26668,R3);
not not8220(N26680,in0);
not not8221(N26704,R2);
not not8222(N26716,in0);
not not8223(N26728,R1);
not not8224(N26740,in1);
not not8225(N26741,R0);
not not8226(N26742,R1);
not not8227(N26752,R0);
not not8228(N26753,R2);
not not8229(N26764,R0);
not not8230(N26765,R1);
not not8231(N26776,in1);
not not8232(N26788,in0);
not not8233(N26789,R0);
not not8234(N26812,in0);
not not8235(N26813,in2);
not not8236(N26824,in0);
not not8237(N26836,in0);
not not8238(N26837,R3);
not not8239(N26848,in2);
not not8240(N26849,R0);
not not8241(N26860,in1);
not not8242(N26861,R0);
not not8243(N26872,in0);
not not8244(N26873,in2);
not not8245(N26884,in1);
not not8246(N26885,R2);
not not8247(N26896,in2);
not not8248(N26897,R2);
not not8249(N26908,R0);
not not8250(N26909,R2);
not not8251(N26920,in0);
not not8252(N26932,in0);
not not8253(N26933,R0);
not not8254(N26944,R1);
not not8255(N26956,in2);
not not8256(N26968,R1);
not not8257(N26980,in1);
not not8258(N26981,R2);
not not8259(N26991,in2);
not not8260(N26992,R2);
not not8261(N27002,R2);
not not8262(N27013,in2);
not not8263(N27014,R2);
not not8264(N27024,R0);
not not8265(N27025,R1);
not not8266(N27035,in0);
not not8267(N27036,in2);
not not8268(N27057,in0);
not not8269(N27058,in1);
not not8270(N27068,in0);
not not8271(N27069,in2);
not not8272(N27079,in0);
not not8273(N27080,in1);
not not8274(N27090,in1);
not not8275(N27101,in0);
not not8276(N27134,in0);
not not8277(N27145,R0);
not not8278(N27166,R3);
not not8279(N27176,R1);
not not8280(N27186,R1);
not not8281(N27196,R3);
not not8282(N27205,in1);
not not8283(N27206,in2);
not not8284(N27207,R0);
not not8285(N27208,R1);
not not8286(N27209,R2);
not not8287(N27210,R4);
not not8288(N27211,R5);
not not8289(N27221,in0);
not not8290(N27222,in1);
not not8291(N27223,R0);
not not8292(N27224,R2);
not not8293(N27225,R4);
not not8294(N27226,R5);
not not8295(N27237,in0);
not not8296(N27238,in1);
not not8297(N27239,in2);
not not8298(N27240,R2);
not not8299(N27241,R3);
not not8300(N27242,R4);
not not8301(N27253,R0);
not not8302(N27254,R2);
not not8303(N27255,R3);
not not8304(N27256,R4);
not not8305(N27257,R5);
not not8306(N27268,R0);
not not8307(N27269,R2);
not not8308(N27270,R3);
not not8309(N27271,R4);
not not8310(N27272,R5);
not not8311(N27283,in1);
not not8312(N27284,in2);
not not8313(N27285,R0);
not not8314(N27286,R1);
not not8315(N27287,R4);
not not8316(N27298,in1);
not not8317(N27299,R0);
not not8318(N27300,R1);
not not8319(N27301,R2);
not not8320(N27302,R4);
not not8321(N27303,R5);
not not8322(N27313,in0);
not not8323(N27314,in1);
not not8324(N27315,in2);
not not8325(N27316,R1);
not not8326(N27317,R4);
not not8327(N27318,R5);
not not8328(N27328,in2);
not not8329(N27329,R0);
not not8330(N27330,R1);
not not8331(N27331,R2);
not not8332(N27332,R3);
not not8333(N27333,R5);
not not8334(N27343,in0);
not not8335(N27344,in1);
not not8336(N27345,R1);
not not8337(N27346,R2);
not not8338(N27347,R3);
not not8339(N27358,in0);
not not8340(N27359,in2);
not not8341(N27360,R1);
not not8342(N27361,R2);
not not8343(N27362,R4);
not not8344(N27373,in0);
not not8345(N27374,R0);
not not8346(N27375,R2);
not not8347(N27376,R4);
not not8348(N27377,R5);
not not8349(N27388,in2);
not not8350(N27389,R0);
not not8351(N27390,R1);
not not8352(N27391,R2);
not not8353(N27392,R4);
not not8354(N27393,R5);
not not8355(N27403,in0);
not not8356(N27404,in1);
not not8357(N27405,R1);
not not8358(N27406,R3);
not not8359(N27407,R4);
not not8360(N27408,R5);
not not8361(N27418,in0);
not not8362(N27419,R0);
not not8363(N27420,R1);
not not8364(N27421,R2);
not not8365(N27422,R5);
not not8366(N27432,in0);
not not8367(N27433,R0);
not not8368(N27434,R1);
not not8369(N27435,R2);
not not8370(N27446,in2);
not not8371(N27447,R0);
not not8372(N27448,R1);
not not8373(N27449,R5);
not not8374(N27460,R0);
not not8375(N27461,R1);
not not8376(N27462,R3);
not not8377(N27463,R5);
not not8378(N27474,in2);
not not8379(N27475,R0);
not not8380(N27476,R1);
not not8381(N27477,R2);
not not8382(N27488,in0);
not not8383(N27489,R0);
not not8384(N27490,R4);
not not8385(N27491,R5);
not not8386(N27502,R0);
not not8387(N27503,R1);
not not8388(N27504,R3);
not not8389(N27505,R4);
not not8390(N27506,R5);
not not8391(N27516,R0);
not not8392(N27517,R1);
not not8393(N27518,R3);
not not8394(N27519,R4);
not not8395(N27520,R5);
not not8396(N27530,in0);
not not8397(N27531,in2);
not not8398(N27532,R1);
not not8399(N27533,R2);
not not8400(N27534,R4);
not not8401(N27544,in2);
not not8402(N27545,R0);
not not8403(N27546,R2);
not not8404(N27547,R4);
not not8405(N27548,R5);
not not8406(N27558,in0);
not not8407(N27559,in2);
not not8408(N27560,R1);
not not8409(N27561,R2);
not not8410(N27562,R4);
not not8411(N27572,in2);
not not8412(N27573,R2);
not not8413(N27574,R3);
not not8414(N27575,R4);
not not8415(N27586,in1);
not not8416(N27587,R2);
not not8417(N27588,R3);
not not8418(N27589,R4);
not not8419(N27600,in2);
not not8420(N27601,R0);
not not8421(N27602,R1);
not not8422(N27603,R3);
not not8423(N27604,R5);
not not8424(N27614,in1);
not not8425(N27615,R0);
not not8426(N27616,R1);
not not8427(N27617,R3);
not not8428(N27618,R5);
not not8429(N27628,in1);
not not8430(N27629,R2);
not not8431(N27630,R3);
not not8432(N27631,R4);
not not8433(N27642,in2);
not not8434(N27643,R1);
not not8435(N27644,R2);
not not8436(N27645,R4);
not not8437(N27656,in0);
not not8438(N27657,in1);
not not8439(N27658,R1);
not not8440(N27659,R2);
not not8441(N27660,R4);
not not8442(N27670,in0);
not not8443(N27671,in2);
not not8444(N27672,R3);
not not8445(N27673,R5);
not not8446(N27684,in0);
not not8447(N27685,in1);
not not8448(N27686,in2);
not not8449(N27687,R4);
not not8450(N27688,R5);
not not8451(N27698,in0);
not not8452(N27699,in1);
not not8453(N27700,in2);
not not8454(N27701,R3);
not not8455(N27702,R4);
not not8456(N27712,in2);
not not8457(N27713,R2);
not not8458(N27714,R3);
not not8459(N27715,R4);
not not8460(N27726,in0);
not not8461(N27727,in2);
not not8462(N27728,R0);
not not8463(N27729,R2);
not not8464(N27730,R5);
not not8465(N27740,in0);
not not8466(N27741,in2);
not not8467(N27742,R2);
not not8468(N27743,R3);
not not8469(N27754,in1);
not not8470(N27755,R4);
not not8471(N27756,R5);
not not8472(N27767,in1);
not not8473(N27768,R1);
not not8474(N27769,R2);
not not8475(N27770,R4);
not not8476(N27780,in0);
not not8477(N27781,in1);
not not8478(N27782,R1);
not not8479(N27783,R3);
not not8480(N27793,in0);
not not8481(N27794,R1);
not not8482(N27795,R2);
not not8483(N27796,R5);
not not8484(N27806,in1);
not not8485(N27807,R2);
not not8486(N27808,R4);
not not8487(N27809,R5);
not not8488(N27819,in0);
not not8489(N27820,in2);
not not8490(N27821,R2);
not not8491(N27822,R4);
not not8492(N27832,in2);
not not8493(N27833,R1);
not not8494(N27834,R2);
not not8495(N27835,R4);
not not8496(N27845,in0);
not not8497(N27846,in1);
not not8498(N27847,R5);
not not8499(N27858,in2);
not not8500(N27859,R0);
not not8501(N27860,R2);
not not8502(N27861,R3);
not not8503(N27862,R5);
not not8504(N27871,in1);
not not8505(N27872,R0);
not not8506(N27873,R1);
not not8507(N27874,R4);
not not8508(N27884,in1);
not not8509(N27885,R1);
not not8510(N27886,R2);
not not8511(N27887,R4);
not not8512(N27888,R5);
not not8513(N27897,in1);
not not8514(N27898,R0);
not not8515(N27899,R3);
not not8516(N27900,R4);
not not8517(N27910,R0);
not not8518(N27911,R3);
not not8519(N27912,R4);
not not8520(N27913,R5);
not not8521(N27923,R1);
not not8522(N27924,R2);
not not8523(N27925,R3);
not not8524(N27926,R5);
not not8525(N27936,in0);
not not8526(N27937,R0);
not not8527(N27938,R5);
not not8528(N27949,in2);
not not8529(N27950,R0);
not not8530(N27951,R3);
not not8531(N27952,R5);
not not8532(N27962,in0);
not not8533(N27963,R2);
not not8534(N27964,R3);
not not8535(N27965,R5);
not not8536(N27975,in1);
not not8537(N27976,R0);
not not8538(N27977,R3);
not not8539(N27978,R4);
not not8540(N27988,in0);
not not8541(N27989,in1);
not not8542(N27990,R3);
not not8543(N27991,R5);
not not8544(N28001,in0);
not not8545(N28002,in1);
not not8546(N28003,R2);
not not8547(N28004,R3);
not not8548(N28014,in1);
not not8549(N28015,R0);
not not8550(N28016,R1);
not not8551(N28017,R3);
not not8552(N28027,in1);
not not8553(N28028,R0);
not not8554(N28029,R3);
not not8555(N28030,R4);
not not8556(N28040,R2);
not not8557(N28041,R3);
not not8558(N28042,R4);
not not8559(N28053,in1);
not not8560(N28054,R0);
not not8561(N28055,R2);
not not8562(N28056,R4);
not not8563(N28066,R1);
not not8564(N28067,R2);
not not8565(N28068,R4);
not not8566(N28079,in0);
not not8567(N28080,R1);
not not8568(N28081,R2);
not not8569(N28082,R4);
not not8570(N28092,in1);
not not8571(N28093,R0);
not not8572(N28094,R1);
not not8573(N28095,R4);
not not8574(N28096,R5);
not not8575(N28105,in2);
not not8576(N28106,R0);
not not8577(N28107,R3);
not not8578(N28108,R4);
not not8579(N28118,in0);
not not8580(N28119,in2);
not not8581(N28120,R2);
not not8582(N28121,R3);
not not8583(N28131,in0);
not not8584(N28132,in1);
not not8585(N28133,in2);
not not8586(N28134,R2);
not not8587(N28144,in2);
not not8588(N28145,R0);
not not8589(N28146,R1);
not not8590(N28147,R3);
not not8591(N28157,in1);
not not8592(N28158,in2);
not not8593(N28159,R0);
not not8594(N28160,R1);
not not8595(N28170,R0);
not not8596(N28171,R5);
not not8597(N28182,R2);
not not8598(N28183,R3);
not not8599(N28184,R4);
not not8600(N28194,in2);
not not8601(N28195,R5);
not not8602(N28206,R0);
not not8603(N28207,R2);
not not8604(N28218,in0);
not not8605(N28219,in2);
not not8606(N28220,R4);
not not8607(N28230,R0);
not not8608(N28231,R1);
not not8609(N28242,in0);
not not8610(N28243,R0);
not not8611(N28244,R5);
not not8612(N28254,R1);
not not8613(N28255,R2);
not not8614(N28256,R4);
not not8615(N28266,R0);
not not8616(N28267,R2);
not not8617(N28268,R4);
not not8618(N28278,in0);
not not8619(N28279,in2);
not not8620(N28280,R4);
not not8621(N28290,in0);
not not8622(N28291,R3);
not not8623(N28292,R4);
not not8624(N28293,R5);
not not8625(N28302,R0);
not not8626(N28303,R2);
not not8627(N28304,R4);
not not8628(N28305,R5);
not not8629(N28314,R0);
not not8630(N28315,R2);
not not8631(N28316,R4);
not not8632(N28326,in0);
not not8633(N28327,in1);
not not8634(N28328,R5);
not not8635(N28338,R1);
not not8636(N28339,R2);
not not8637(N28340,R4);
not not8638(N28341,R5);
not not8639(N28350,in1);
not not8640(N28351,R1);
not not8641(N28352,R4);
not not8642(N28353,R5);
not not8643(N28362,in1);
not not8644(N28363,R0);
not not8645(N28364,R1);
not not8646(N28374,in2);
not not8647(N28375,R3);
not not8648(N28376,R4);
not not8649(N28386,in0);
not not8650(N28387,in2);
not not8651(N28388,R0);
not not8652(N28389,R2);
not not8653(N28398,in0);
not not8654(N28399,in2);
not not8655(N28400,R3);
not not8656(N28410,in2);
not not8657(N28411,R3);
not not8658(N28412,R5);
not not8659(N28422,in1);
not not8660(N28423,R0);
not not8661(N28424,R4);
not not8662(N28434,in0);
not not8663(N28435,R0);
not not8664(N28436,R5);
not not8665(N28446,in0);
not not8666(N28447,in2);
not not8667(N28448,R1);
not not8668(N28449,R5);
not not8669(N28458,in0);
not not8670(N28459,in1);
not not8671(N28460,R4);
not not8672(N28461,R5);
not not8673(N28470,in0);
not not8674(N28471,in1);
not not8675(N28472,R4);
not not8676(N28482,in2);
not not8677(N28483,R0);
not not8678(N28484,R5);
not not8679(N28494,in1);
not not8680(N28495,R1);
not not8681(N28496,R3);
not not8682(N28506,R0);
not not8683(N28507,R1);
not not8684(N28508,R5);
not not8685(N28518,in2);
not not8686(N28519,R4);
not not8687(N28530,in0);
not not8688(N28531,in1);
not not8689(N28532,R0);
not not8690(N28533,R4);
not not8691(N28542,R0);
not not8692(N28543,R3);
not not8693(N28544,R5);
not not8694(N28554,in0);
not not8695(N28555,in1);
not not8696(N28556,R1);
not not8697(N28566,R1);
not not8698(N28567,R2);
not not8699(N28568,R4);
not not8700(N28578,R2);
not not8701(N28579,R4);
not not8702(N28580,R5);
not not8703(N28590,in2);
not not8704(N28591,R0);
not not8705(N28592,R1);
not not8706(N28602,in0);
not not8707(N28603,in1);
not not8708(N28604,in2);
not not8709(N28614,in2);
not not8710(N28615,R2);
not not8711(N28626,R1);
not not8712(N28627,R3);
not not8713(N28638,in0);
not not8714(N28639,in1);
not not8715(N28650,in1);
not not8716(N28651,in2);
not not8717(N28652,R3);
not not8718(N28662,R5);
not not8719(N28673,R5);
not not8720(N28684,in1);
not not8721(N28685,R0);
not not8722(N28686,R5);
not not8723(N28695,R0);
not not8724(N28696,R2);
not not8725(N28697,R5);
not not8726(N28706,in0);
not not8727(N28707,R1);
not not8728(N28717,in1);
not not8729(N28718,R4);
not not8730(N28728,R1);
not not8731(N28729,R3);
not not8732(N28739,in1);
not not8733(N28740,R5);
not not8734(N28750,R1);
not not8735(N28751,R4);
not not8736(N28761,R3);
not not8737(N28762,R5);
not not8738(N28772,R3);
not not8739(N28773,R5);
not not8740(N28783,in2);
not not8741(N28784,R2);
not not8742(N28794,in1);
not not8743(N28795,R0);
not not8744(N28796,R3);
not not8745(N28805,in0);
not not8746(N28806,R2);
not not8747(N28816,in0);
not not8748(N28817,R4);
not not8749(N28818,R5);
not not8750(N28827,R0);
not not8751(N28828,R4);
not not8752(N28829,R5);
not not8753(N28838,in2);
not not8754(N28839,R3);
not not8755(N28849,in2);
not not8756(N28860,R3);
not not8757(N28861,R4);
not not8758(N28871,R0);
not not8759(N28872,R4);
not not8760(N28882,R2);
not not8761(N28883,R3);
not not8762(N28893,R0);
not not8763(N28894,R5);
not not8764(N28904,R1);
not not8765(N28905,R4);
not not8766(N28915,in0);
not not8767(N28916,in2);
not not8768(N28917,R0);
not not8769(N28926,in2);
not not8770(N28927,R0);
not not8771(N28928,R3);
not not8772(N28937,R0);
not not8773(N28947,R3);
not not8774(N28957,in2);
not not8775(N28958,R1);
not not8776(N28967,in0);
not not8777(N28968,R0);
not not8778(N28977,R1);
not not8779(N28978,R4);
not not8780(N28987,R4);
not not8781(N28988,R5);
not not8782(N28997,in0);
not not8783(N28998,in1);
not not8784(N29007,R1);
not not8785(N29017,in2);
not not8786(N29018,R3);
not not8787(N29027,R4);
not not8788(N29037,in1);
not not8789(N29038,R3);
not not8790(N29047,R0);
not not8791(N29048,R5);
not not8792(N29057,R2);
not not8793(N29065,in0);
not not8794(N29066,R1);
not not8795(N29067,R2);
not not8796(N29068,R3);
not not8797(N29069,R6);
not not8798(N29070,R7);
not not8799(N29078,R0);
not not8800(N29079,R1);
not not8801(N29080,R2);
not not8802(N29081,R4);
not not8803(N29082,R5);
not not8804(N29083,R7);
not not8805(N29091,in1);
not not8806(N29092,R0);
not not8807(N29093,R2);
not not8808(N29094,R4);
not not8809(N29095,R5);
not not8810(N29096,R7);
not not8811(N29104,R0);
not not8812(N29105,R2);
not not8813(N29106,R5);
not not8814(N29107,R6);
not not8815(N29108,R7);
not not8816(N29116,in2);
not not8817(N29117,R2);
not not8818(N29118,R5);
not not8819(N29119,R6);
not not8820(N29120,R7);
not not8821(N29128,R0);
not not8822(N29129,R4);
not not8823(N29130,R5);
not not8824(N29131,R6);
not not8825(N29132,R7);
not not8826(N29140,R1);
not not8827(N29141,R3);
not not8828(N29142,R4);
not not8829(N29143,R5);
not not8830(N29144,R7);
not not8831(N29152,R1);
not not8832(N29153,R2);
not not8833(N29154,R3);
not not8834(N29155,R6);
not not8835(N29156,R7);
not not8836(N29164,R1);
not not8837(N29165,R4);
not not8838(N29166,R5);
not not8839(N29167,R7);
not not8840(N29175,R1);
not not8841(N29176,R4);
not not8842(N29177,R5);
not not8843(N29178,R7);
not not8844(N29186,R3);
not not8845(N29187,R5);
not not8846(N29188,R6);
not not8847(N29189,R7);
not not8848(N29197,R1);
not not8849(N29198,R2);
not not8850(N29199,R5);
not not8851(N29200,R6);
not not8852(N29208,R1);
not not8853(N29209,R2);
not not8854(N29210,R5);
not not8855(N29211,R6);
not not8856(N29219,in1);
not not8857(N29220,R2);
not not8858(N29221,R3);
not not8859(N29222,R7);
not not8860(N29230,in2);
not not8861(N29231,R2);
not not8862(N29232,R3);
not not8863(N29233,R7);
not not8864(N29241,in1);
not not8865(N29242,R3);
not not8866(N29243,R6);
not not8867(N29251,R1);
not not8868(N29252,R5);
not not8869(N29253,R6);
not not8870(N29261,R2);
not not8871(N29262,R6);
not not8872(N29269,R2);
not not8873(N29270,R3);
not not8874(N29271,R5);
not not8875(N29272,R6);
not not8876(N24441,R3);
not not8877(N24442,R6);
not not8878(N24443,R7);
not not8879(N24457,R3);
not not8880(N24458,R4);
not not8881(N24459,R5);
not not8882(N24460,R7);
not not8883(N24475,R3);
not not8884(N24476,R5);
not not8885(N24477,R6);
not not8886(N24491,R4);
not not8887(N24492,R5);
not not8888(N24493,R6);
not not8889(N24494,R7);
not not8890(N24508,R3);
not not8891(N24509,R5);
not not8892(N24510,R6);
not not8893(N24511,R7);
not not8894(N24526,R5);
not not8895(N24527,R6);
not not8896(N24528,R7);
not not8897(N24543,R3);
not not8898(N24544,R5);
not not8899(N24545,R6);
not not8900(N24560,R4);
not not8901(N24561,R6);
not not8902(N24562,R7);
not not8903(N24576,R5);
not not8904(N24577,R6);
not not8905(N24578,R7);
not not8906(N24592,R4);
not not8907(N24593,R5);
not not8908(N24594,R6);
not not8909(N24608,R4);
not not8910(N24609,R5);
not not8911(N24610,R6);
not not8912(N24624,R5);
not not8913(N24625,R6);
not not8914(N24626,R7);
not not8915(N24640,R4);
not not8916(N24641,R5);
not not8917(N24642,R6);
not not8918(N24655,R4);
not not8919(N24656,R5);
not not8920(N24657,R6);
not not8921(N24658,R7);
not not8922(N24672,R4);
not not8923(N24673,R6);
not not8924(N24674,R7);
not not8925(N24689,R4);
not not8926(N24690,R6);
not not8927(N24705,R5);
not not8928(N24706,R7);
not not8929(N24721,R4);
not not8930(N24722,R7);
not not8931(N24736,R3);
not not8932(N24737,R6);
not not8933(N24738,R7);
not not8934(N24752,R5);
not not8935(N24753,R6);
not not8936(N24754,R7);
not not8937(N24768,R4);
not not8938(N24769,R5);
not not8939(N24770,R6);
not not8940(N24784,R3);
not not8941(N24785,R4);
not not8942(N24786,R5);
not not8943(N24799,R4);
not not8944(N24800,R5);
not not8945(N24801,R6);
not not8946(N24802,R7);
not not8947(N24816,R4);
not not8948(N24817,R5);
not not8949(N24818,R6);
not not8950(N24832,R4);
not not8951(N24833,R5);
not not8952(N24834,R6);
not not8953(N24847,R3);
not not8954(N24848,R4);
not not8955(N24849,R6);
not not8956(N24850,R7);
not not8957(N24864,R4);
not not8958(N24865,R6);
not not8959(N24866,R7);
not not8960(N24878,R4);
not not8961(N24879,R5);
not not8962(N24880,R6);
not not8963(N24881,R7);
not not8964(N24895,R4);
not not8965(N24896,R5);
not not8966(N24909,R4);
not not8967(N24910,R6);
not not8968(N24911,R7);
not not8969(N24924,R5);
not not8970(N24925,R6);
not not8971(N24926,R7);
not not8972(N24940,R5);
not not8973(N24941,R7);
not not8974(N24955,R3);
not not8975(N24956,R6);
not not8976(N24970,R5);
not not8977(N24971,R6);
not not8978(N24986,R5);
not not8979(N25000,R6);
not not8980(N25001,R7);
not not8981(N25015,R6);
not not8982(N25016,R7);
not not8983(N25029,R5);
not not8984(N25030,R6);
not not8985(N25031,R7);
not not8986(N25044,R4);
not not8987(N25045,R5);
not not8988(N25046,R7);
not not8989(N25060,R4);
not not8990(N25061,R6);
not not8991(N25075,R4);
not not8992(N25076,R5);
not not8993(N25090,R5);
not not8994(N25091,R7);
not not8995(N25105,R5);
not not8996(N25106,R7);
not not8997(N25120,R4);
not not8998(N25121,R7);
not not8999(N25135,R6);
not not9000(N25136,R7);
not not9001(N25149,R4);
not not9002(N25150,R6);
not not9003(N25151,R7);
not not9004(N25165,R5);
not not9005(N25166,R6);
not not9006(N25181,R5);
not not9007(N25196,R5);
not not9008(N25210,R4);
not not9009(N25211,R6);
not not9010(N25224,R4);
not not9011(N25225,R6);
not not9012(N25226,R7);
not not9013(N25239,R4);
not not9014(N25240,R6);
not not9015(N25241,R7);
not not9016(N25255,R6);
not not9017(N25256,R7);
not not9018(N25269,R4);
not not9019(N25270,R7);
not not9020(N25282,R4);
not not9021(N25283,R5);
not not9022(N25284,R6);
not not9023(N25297,R5);
not not9024(N25298,R6);
not not9025(N25311,R6);
not not9026(N25312,R7);
not not9027(N25325,R5);
not not9028(N25326,R6);
not not9029(N25339,R4);
not not9030(N25340,R5);
not not9031(N25353,R4);
not not9032(N25354,R7);
not not9033(N25367,R6);
not not9034(N25368,R7);
not not9035(N25380,R3);
not not9036(N25381,R4);
not not9037(N25382,R5);
not not9038(N25394,R4);
not not9039(N25395,R5);
not not9040(N25396,R7);
not not9041(N25408,R4);
not not9042(N25409,R5);
not not9043(N25410,R7);
not not9044(N25423,R4);
not not9045(N25424,R5);
not not9046(N25437,R5);
not not9047(N25438,R6);
not not9048(N25452,R5);
not not9049(N25465,R6);
not not9050(N25466,R7);
not not9051(N25480,R7);
not not9052(N25494,R6);
not not9053(N25508,R7);
not not9054(N25520,R4);
not not9055(N25521,R5);
not not9056(N25522,R7);
not not9057(N25535,R4);
not not9058(N25536,R6);
not not9059(N25549,R4);
not not9060(N25550,R6);
not not9061(N25562,R4);
not not9062(N25563,R6);
not not9063(N25564,R7);
not not9064(N25578,R6);
not not9065(N25590,R4);
not not9066(N25591,R5);
not not9067(N25592,R6);
not not9068(N25604,R4);
not not9069(N25605,R6);
not not9070(N25606,R7);
not not9071(N25619,R4);
not not9072(N25620,R6);
not not9073(N25634,R5);
not not9074(N25646,R4);
not not9075(N25647,R6);
not not9076(N25648,R7);
not not9077(N25661,R4);
not not9078(N25662,R6);
not not9079(N25674,R3);
not not9080(N25675,R4);
not not9081(N25676,R7);
not not9082(N25689,R4);
not not9083(N25690,R6);
not not9084(N25703,R4);
not not9085(N25704,R5);
not not9086(N25717,R4);
not not9087(N25718,R6);
not not9088(N25731,R4);
not not9089(N25732,R6);
not not9090(N25746,R6);
not not9091(N25760,R6);
not not9092(N25773,R4);
not not9093(N25774,R6);
not not9094(N25787,R4);
not not9095(N25788,R7);
not not9096(N25800,R4);
not not9097(N25801,R6);
not not9098(N25802,R7);
not not9099(N25816,R5);
not not9100(N25829,R4);
not not9101(N25830,R6);
not not9102(N25842,R4);
not not9103(N25843,R5);
not not9104(N25844,R6);
not not9105(N25856,R5);
not not9106(N25857,R6);
not not9107(N25858,R7);
not not9108(N25872,R7);
not not9109(N25885,R5);
not not9110(N25886,R6);
not not9111(N25900,R6);
not not9112(N25914,R5);
not not9113(N25928,R5);
not not9114(N25941,R4);
not not9115(N25942,R5);
not not9116(N25955,R4);
not not9117(N25956,R6);
not not9118(N25968,R4);
not not9119(N25969,R5);
not not9120(N25970,R6);
not not9121(N25982,R4);
not not9122(N25983,R6);
not not9123(N25984,R7);
not not9124(N25996,R3);
not not9125(N25997,R5);
not not9126(N25998,R7);
not not9127(N26010,R3);
not not9128(N26011,R4);
not not9129(N26012,R5);
not not9130(N26025,R6);
not not9131(N26026,R7);
not not9132(N26040,R6);
not not9133(N26053,R3);
not not9134(N26054,R6);
not not9135(N26066,R3);
not not9136(N26067,R6);
not not9137(N26068,R7);
not not9138(N26080,R3);
not not9139(N26081,R6);
not not9140(N26082,R7);
not not9141(N26094,R3);
not not9142(N26095,R6);
not not9143(N26096,R7);
not not9144(N26109,R6);
not not9145(N26110,R7);
not not9146(N26123,R5);
not not9147(N26124,R6);
not not9148(N26137,R5);
not not9149(N26138,R6);
not not9150(N26149,R5);
not not9151(N26150,R6);
not not9152(N26151,R7);
not not9153(N26163,R4);
not not9154(N26164,R7);
not not9155(N26176,R4);
not not9156(N26177,R6);
not not9157(N26190,R7);
not not9158(N26202,R5);
not not9159(N26203,R7);
not not9160(N26215,R4);
not not9161(N26216,R5);
not not9162(N26229,R6);
not not9163(N26241,R4);
not not9164(N26242,R7);
not not9165(N26254,R4);
not not9166(N26255,R6);
not not9167(N26268,R7);
not not9168(N26280,R4);
not not9169(N26281,R5);
not not9170(N26294,R7);
not not9171(N26305,R4);
not not9172(N26306,R6);
not not9173(N26307,R7);
not not9174(N26320,R5);
not not9175(N26333,R5);
not not9176(N26346,R7);
not not9177(N26359,R7);
not not9178(N26372,R5);
not not9179(N26384,R5);
not not9180(N26385,R7);
not not9181(N26398,R3);
not not9182(N26410,R4);
not not9183(N26411,R5);
not not9184(N26423,R3);
not not9185(N26424,R5);
not not9186(N26437,R6);
not not9187(N26450,R6);
not not9188(N26461,R3);
not not9189(N26462,R4);
not not9190(N26463,R6);
not not9191(N26475,R5);
not not9192(N26476,R7);
not not9193(N26487,R4);
not not9194(N26488,R6);
not not9195(N26489,R7);
not not9196(N26502,R5);
not not9197(N26514,R6);
not not9198(N26525,R4);
not not9199(N26526,R7);
not not9200(N26538,R7);
not not9201(N26550,R6);
not not9202(N26561,R4);
not not9203(N26562,R6);
not not9204(N26574,R5);
not not9205(N26585,R3);
not not9206(N26586,R7);
not not9207(N26597,R3);
not not9208(N26598,R6);
not not9209(N26609,R5);
not not9210(N26610,R7);
not not9211(N26622,R6);
not not9212(N26634,R7);
not not9213(N26646,R7);
not not9214(N26658,R7);
not not9215(N26669,R4);
not not9216(N26670,R6);
not not9217(N26681,R5);
not not9218(N26682,R6);
not not9219(N26692,R4);
not not9220(N26693,R5);
not not9221(N26694,R6);
not not9222(N26705,R3);
not not9223(N26706,R6);
not not9224(N26717,R6);
not not9225(N26718,R7);
not not9226(N26729,R4);
not not9227(N26730,R6);
not not9228(N26754,R6);
not not9229(N26766,R6);
not not9230(N26777,R6);
not not9231(N26778,R7);
not not9232(N26790,R7);
not not9233(N26800,R4);
not not9234(N26801,R6);
not not9235(N26802,R7);
not not9236(N26814,R7);
not not9237(N26825,R5);
not not9238(N26826,R7);
not not9239(N26838,R5);
not not9240(N26850,R7);
not not9241(N26862,R7);
not not9242(N26874,R4);
not not9243(N26886,R6);
not not9244(N26898,R6);
not not9245(N26910,R7);
not not9246(N26921,R3);
not not9247(N26922,R7);
not not9248(N26934,R7);
not not9249(N26945,R6);
not not9250(N26946,R7);
not not9251(N26957,R6);
not not9252(N26958,R7);
not not9253(N26969,R5);
not not9254(N26970,R6);
not not9255(N27003,R5);
not not9256(N27046,R3);
not not9257(N27047,R5);
not not9258(N27091,R3);
not not9259(N27102,R5);
not not9260(N27112,R5);
not not9261(N27113,R6);
not not9262(N27123,R6);
not not9263(N27124,R7);
not not9264(N27135,R4);
not not9265(N27146,R7);
not not9266(N27156,R3);
not not9267(N27212,R6);
not not9268(N27227,R6);
not not9269(N27228,R7);
not not9270(N27243,R5);
not not9271(N27244,R6);
not not9272(N27258,R6);
not not9273(N27259,R7);
not not9274(N27273,R6);
not not9275(N27274,R7);
not not9276(N27288,R6);
not not9277(N27289,R7);
not not9278(N27304,R7);
not not9279(N27319,R7);
not not9280(N27334,R7);
not not9281(N27348,R5);
not not9282(N27349,R7);
not not9283(N27363,R5);
not not9284(N27364,R6);
not not9285(N27378,R6);
not not9286(N27379,R7);
not not9287(N27394,R6);
not not9288(N27409,R7);
not not9289(N27423,R6);
not not9290(N27436,R5);
not not9291(N27437,R6);
not not9292(N27450,R6);
not not9293(N27451,R7);
not not9294(N27464,R6);
not not9295(N27465,R7);
not not9296(N27478,R6);
not not9297(N27479,R7);
not not9298(N27492,R6);
not not9299(N27493,R7);
not not9300(N27507,R6);
not not9301(N27521,R6);
not not9302(N27535,R7);
not not9303(N27549,R7);
not not9304(N27563,R6);
not not9305(N27576,R5);
not not9306(N27577,R6);
not not9307(N27590,R5);
not not9308(N27591,R6);
not not9309(N27605,R7);
not not9310(N27619,R7);
not not9311(N27632,R6);
not not9312(N27633,R7);
not not9313(N27646,R6);
not not9314(N27647,R7);
not not9315(N27661,R7);
not not9316(N27674,R6);
not not9317(N27675,R7);
not not9318(N27689,R6);
not not9319(N27703,R5);
not not9320(N27716,R6);
not not9321(N27717,R7);
not not9322(N27731,R7);
not not9323(N27744,R4);
not not9324(N27745,R5);
not not9325(N27757,R6);
not not9326(N27758,R7);
not not9327(N27771,R6);
not not9328(N27784,R7);
not not9329(N27797,R7);
not not9330(N27810,R6);
not not9331(N27823,R6);
not not9332(N27836,R6);
not not9333(N27848,R6);
not not9334(N27849,R7);
not not9335(N27875,R6);
not not9336(N27901,R6);
not not9337(N27914,R7);
not not9338(N27927,R7);
not not9339(N27939,R6);
not not9340(N27940,R7);
not not9341(N27953,R6);
not not9342(N27966,R6);
not not9343(N27979,R5);
not not9344(N27992,R6);
not not9345(N28005,R7);
not not9346(N28018,R6);
not not9347(N28031,R7);
not not9348(N28043,R5);
not not9349(N28044,R6);
not not9350(N28057,R6);
not not9351(N28069,R6);
not not9352(N28070,R7);
not not9353(N28083,R7);
not not9354(N28109,R5);
not not9355(N28122,R7);
not not9356(N28135,R4);
not not9357(N28148,R6);
not not9358(N28161,R6);
not not9359(N28172,R6);
not not9360(N28173,R7);
not not9361(N28185,R7);
not not9362(N28196,R6);
not not9363(N28197,R7);
not not9364(N28208,R6);
not not9365(N28209,R7);
not not9366(N28221,R6);
not not9367(N28232,R6);
not not9368(N28233,R7);
not not9369(N28245,R7);
not not9370(N28257,R7);
not not9371(N28269,R7);
not not9372(N28281,R7);
not not9373(N28317,R5);
not not9374(N28329,R7);
not not9375(N28365,R7);
not not9376(N28377,R6);
not not9377(N28401,R7);
not not9378(N28413,R7);
not not9379(N28425,R5);
not not9380(N28437,R7);
not not9381(N28473,R6);
not not9382(N28485,R7);
not not9383(N28497,R6);
not not9384(N28509,R7);
not not9385(N28520,R6);
not not9386(N28521,R7);
not not9387(N28545,R6);
not not9388(N28557,R5);
not not9389(N28569,R6);
not not9390(N28581,R6);
not not9391(N28593,R7);
not not9392(N28605,R5);
not not9393(N28616,R5);
not not9394(N28617,R7);
not not9395(N28628,R6);
not not9396(N28629,R7);
not not9397(N28640,R6);
not not9398(N28641,R7);
not not9399(N28653,R5);
not not9400(N28663,R6);
not not9401(N28664,R7);
not not9402(N28674,R6);
not not9403(N28675,R7);
not not9404(N28708,R7);
not not9405(N28719,R7);
not not9406(N28730,R6);
not not9407(N28741,R6);
not not9408(N28752,R7);
not not9409(N28763,R6);
not not9410(N28774,R6);
not not9411(N28785,R7);
not not9412(N28807,R7);
not not9413(N28840,R6);
not not9414(N28850,R5);
not not9415(N28851,R6);
not not9416(N28862,R6);
not not9417(N28873,R5);
not not9418(N28884,R7);
not not9419(N28895,R7);
not not9420(N28906,R5);
not not9421(N28938,R6);
not not9422(N28948,R7);
not not9423(N29008,R6);
not not9424(N29028,R7);
not not9425(N29444,in0);
not not9426(N29445,in2);
not not9427(N29446,R0);
not not9428(N29447,R1);
not not9429(N29462,in0);
not not9430(N29463,in2);
not not9431(N29464,R1);
not not9432(N29480,in0);
not not9433(N29481,in1);
not not9434(N29482,in2);
not not9435(N29497,in0);
not not9436(N29498,in1);
not not9437(N29499,R0);
not not9438(N29514,in0);
not not9439(N29515,in2);
not not9440(N29516,R0);
not not9441(N29517,R1);
not not9442(N29530,in0);
not not9443(N29531,in2);
not not9444(N29532,R0);
not not9445(N29533,R1);
not not9446(N29546,in0);
not not9447(N29547,in1);
not not9448(N29548,R1);
not not9449(N29559,in0);
not not9450(N29560,in1);
not not9451(N29561,in2);
not not9452(N29562,R0);
not not9453(N29563,R1);
not not9454(N29564,R2);
not not9455(N29577,in0);
not not9456(N29578,in1);
not not9457(N29579,in2);
not not9458(N29580,R1);
not not9459(N29581,R2);
not not9460(N29595,in0);
not not9461(N29596,in1);
not not9462(N29597,in2);
not not9463(N29598,R1);
not not9464(N29599,R2);
not not9465(N29613,in0);
not not9466(N29614,in1);
not not9467(N29615,R0);
not not9468(N29616,R3);
not not9469(N29630,in0);
not not9470(N29631,R0);
not not9471(N29632,R1);
not not9472(N29633,R2);
not not9473(N29634,R3);
not not9474(N29647,in0);
not not9475(N29648,in1);
not not9476(N29649,in2);
not not9477(N29650,R0);
not not9478(N29651,R1);
not not9479(N29664,in0);
not not9480(N29665,R0);
not not9481(N29666,R1);
not not9482(N29667,R2);
not not9483(N29681,in0);
not not9484(N29682,R0);
not not9485(N29683,R1);
not not9486(N29684,R2);
not not9487(N29685,R3);
not not9488(N29698,in0);
not not9489(N29699,in2);
not not9490(N29700,R1);
not not9491(N29701,R2);
not not9492(N29702,R3);
not not9493(N29715,in0);
not not9494(N29716,in1);
not not9495(N29717,R0);
not not9496(N29718,R1);
not not9497(N29719,R2);
not not9498(N29731,in0);
not not9499(N29732,in1);
not not9500(N29733,R1);
not not9501(N29734,R2);
not not9502(N29747,in0);
not not9503(N29748,in1);
not not9504(N29749,R0);
not not9505(N29750,R3);
not not9506(N29763,in0);
not not9507(N29764,in1);
not not9508(N29765,in2);
not not9509(N29766,R0);
not not9510(N29767,R3);
not not9511(N29779,in0);
not not9512(N29780,in2);
not not9513(N29781,R1);
not not9514(N29782,R3);
not not9515(N29795,in0);
not not9516(N29796,in1);
not not9517(N29797,R1);
not not9518(N29811,in0);
not not9519(N29812,in1);
not not9520(N29813,R0);
not not9521(N29814,R1);
not not9522(N29815,R3);
not not9523(N29827,in0);
not not9524(N29828,in1);
not not9525(N29829,R0);
not not9526(N29830,R1);
not not9527(N29831,R2);
not not9528(N29843,in0);
not not9529(N29844,in1);
not not9530(N29845,R0);
not not9531(N29846,R2);
not not9532(N29859,in0);
not not9533(N29860,in2);
not not9534(N29861,R2);
not not9535(N29862,R3);
not not9536(N29875,in0);
not not9537(N29876,in1);
not not9538(N29877,in2);
not not9539(N29878,R0);
not not9540(N29879,R2);
not not9541(N29891,in0);
not not9542(N29892,in1);
not not9543(N29893,in2);
not not9544(N29894,R0);
not not9545(N29895,R2);
not not9546(N29907,in0);
not not9547(N29908,in2);
not not9548(N29909,R1);
not not9549(N29910,R3);
not not9550(N29923,in0);
not not9551(N29924,in1);
not not9552(N29925,R0);
not not9553(N29926,R2);
not not9554(N29939,in0);
not not9555(N29940,in1);
not not9556(N29941,in2);
not not9557(N29942,R0);
not not9558(N29943,R3);
not not9559(N29955,in0);
not not9560(N29956,in1);
not not9561(N29957,in2);
not not9562(N29958,R0);
not not9563(N29971,in0);
not not9564(N29972,R0);
not not9565(N29973,R1);
not not9566(N29974,R3);
not not9567(N29987,in0);
not not9568(N29988,R1);
not not9569(N29989,R2);
not not9570(N29990,R3);
not not9571(N30003,in0);
not not9572(N30004,in2);
not not9573(N30005,R0);
not not9574(N30006,R2);
not not9575(N30018,in0);
not not9576(N30019,in2);
not not9577(N30020,R2);
not not9578(N30033,in0);
not not9579(N30034,in1);
not not9580(N30035,R2);
not not9581(N30048,in0);
not not9582(N30049,R0);
not not9583(N30050,R3);
not not9584(N30063,in0);
not not9585(N30064,R0);
not not9586(N30065,R2);
not not9587(N30078,in0);
not not9588(N30079,in1);
not not9589(N30080,R1);
not not9590(N30093,in0);
not not9591(N30094,in1);
not not9592(N30095,in2);
not not9593(N30096,R1);
not not9594(N30097,R2);
not not9595(N30108,in0);
not not9596(N30109,in2);
not not9597(N30110,R0);
not not9598(N30111,R2);
not not9599(N30123,in0);
not not9600(N30124,R0);
not not9601(N30125,R2);
not not9602(N30138,in0);
not not9603(N30139,R3);
not not9604(N30153,in0);
not not9605(N30154,R0);
not not9606(N30155,R1);
not not9607(N30168,in0);
not not9608(N30169,in1);
not not9609(N30170,R2);
not not9610(N30183,in0);
not not9611(N30184,in2);
not not9612(N30185,R0);
not not9613(N30198,in0);
not not9614(N30199,in2);
not not9615(N30200,R3);
not not9616(N30213,in0);
not not9617(N30214,R1);
not not9618(N30215,R2);
not not9619(N30228,in0);
not not9620(N30229,in2);
not not9621(N30230,R0);
not not9622(N30231,R2);
not not9623(N30243,in0);
not not9624(N30244,R0);
not not9625(N30245,R2);
not not9626(N30258,in0);
not not9627(N30259,R0);
not not9628(N30260,R3);
not not9629(N30273,in0);
not not9630(N30274,R1);
not not9631(N30275,R2);
not not9632(N30288,in0);
not not9633(N30289,in1);
not not9634(N30290,R0);
not not9635(N30291,R3);
not not9636(N30303,in0);
not not9637(N30304,in2);
not not9638(N30305,R0);
not not9639(N30306,R3);
not not9640(N30318,in0);
not not9641(N30319,in1);
not not9642(N30320,in2);
not not9643(N30321,R2);
not not9644(N30333,in0);
not not9645(N30334,in1);
not not9646(N30335,R3);
not not9647(N30348,in0);
not not9648(N30349,R0);
not not9649(N30350,R2);
not not9650(N30363,in0);
not not9651(N30364,in1);
not not9652(N30365,in2);
not not9653(N30366,R2);
not not9654(N30378,in0);
not not9655(N30379,R2);
not not9656(N30380,R3);
not not9657(N30393,in0);
not not9658(N30394,in1);
not not9659(N30395,in2);
not not9660(N30396,R3);
not not9661(N30408,in0);
not not9662(N30409,in1);
not not9663(N30410,R3);
not not9664(N30423,in0);
not not9665(N30424,R1);
not not9666(N30425,R3);
not not9667(N30438,in0);
not not9668(N30439,in2);
not not9669(N30440,R2);
not not9670(N30453,in0);
not not9671(N30454,in2);
not not9672(N30455,R3);
not not9673(N30468,in0);
not not9674(N30469,in1);
not not9675(N30470,R0);
not not9676(N30471,R1);
not not9677(N30483,in0);
not not9678(N30484,R2);
not not9679(N30497,in0);
not not9680(N30498,R0);
not not9681(N30499,R3);
not not9682(N30511,in0);
not not9683(N30512,in1);
not not9684(N30513,R3);
not not9685(N30525,in0);
not not9686(N30526,R1);
not not9687(N30527,R2);
not not9688(N30539,in0);
not not9689(N30540,R0);
not not9690(N30541,R1);
not not9691(N30553,in0);
not not9692(N30554,in1);
not not9693(N30555,in2);
not not9694(N30556,R0);
not not9695(N30567,in0);
not not9696(N30568,in1);
not not9697(N30569,R1);
not not9698(N30570,R2);
not not9699(N30581,in0);
not not9700(N30582,R0);
not not9701(N30583,R1);
not not9702(N30595,in0);
not not9703(N30596,in2);
not not9704(N30597,R0);
not not9705(N30609,in0);
not not9706(N30610,R1);
not not9707(N30611,R3);
not not9708(N30623,in0);
not not9709(N30624,in1);
not not9710(N30625,R3);
not not9711(N30637,in0);
not not9712(N30638,R1);
not not9713(N30639,R2);
not not9714(N30651,in0);
not not9715(N30652,in1);
not not9716(N30653,R2);
not not9717(N30665,in0);
not not9718(N30666,R0);
not not9719(N30667,R1);
not not9720(N30668,R3);
not not9721(N30679,in0);
not not9722(N30680,R2);
not not9723(N30681,R3);
not not9724(N30693,in0);
not not9725(N30694,in1);
not not9726(N30707,in0);
not not9727(N30708,in2);
not not9728(N30709,R1);
not not9729(N30721,in0);
not not9730(N30722,in1);
not not9731(N30723,R0);
not not9732(N30724,R2);
not not9733(N30735,in0);
not not9734(N30736,R0);
not not9735(N30737,R2);
not not9736(N30749,in0);
not not9737(N30750,in1);
not not9738(N30751,R0);
not not9739(N30752,R3);
not not9740(N30763,in0);
not not9741(N30764,in2);
not not9742(N30765,R0);
not not9743(N30766,R3);
not not9744(N30777,in0);
not not9745(N30778,R0);
not not9746(N30779,R2);
not not9747(N30791,in0);
not not9748(N30792,in1);
not not9749(N30793,in2);
not not9750(N30794,R0);
not not9751(N30805,in0);
not not9752(N30806,in2);
not not9753(N30807,R1);
not not9754(N30819,in0);
not not9755(N30820,in1);
not not9756(N30821,R1);
not not9757(N30833,in0);
not not9758(N30834,in2);
not not9759(N30847,in0);
not not9760(N30848,R0);
not not9761(N30849,R1);
not not9762(N30861,in0);
not not9763(N30862,in1);
not not9764(N30863,in2);
not not9765(N30864,R1);
not not9766(N30875,in0);
not not9767(N30876,in2);
not not9768(N30877,R1);
not not9769(N30878,R2);
not not9770(N30889,in0);
not not9771(N30890,in1);
not not9772(N30891,R1);
not not9773(N30892,R2);
not not9774(N30903,in0);
not not9775(N30904,in1);
not not9776(N30905,R1);
not not9777(N30917,in0);
not not9778(N30918,in2);
not not9779(N30919,R1);
not not9780(N30931,in0);
not not9781(N30932,R0);
not not9782(N30933,R2);
not not9783(N30945,in0);
not not9784(N30946,in2);
not not9785(N30947,R2);
not not9786(N30959,in0);
not not9787(N30960,R1);
not not9788(N30961,R3);
not not9789(N30973,in0);
not not9790(N30974,in2);
not not9791(N30975,R2);
not not9792(N30986,in0);
not not9793(N30999,in0);
not not9794(N31000,R1);
not not9795(N31001,R2);
not not9796(N31012,in0);
not not9797(N31013,R0);
not not9798(N31025,in0);
not not9799(N31038,in0);
not not9800(N31039,R3);
not not9801(N31051,in0);
not not9802(N31052,R0);
not not9803(N31064,in0);
not not9804(N31065,R0);
not not9805(N31066,R2);
not not9806(N31077,in0);
not not9807(N31078,in2);
not not9808(N31079,R3);
not not9809(N31090,in0);
not not9810(N31091,R0);
not not9811(N31092,R1);
not not9812(N31103,in0);
not not9813(N31104,R0);
not not9814(N31105,R2);
not not9815(N31116,in0);
not not9816(N31117,R2);
not not9817(N31129,in0);
not not9818(N31130,in1);
not not9819(N31131,R1);
not not9820(N31142,in0);
not not9821(N31143,R0);
not not9822(N31155,in0);
not not9823(N31156,in1);
not not9824(N31168,in0);
not not9825(N31169,in1);
not not9826(N31170,R2);
not not9827(N31181,in0);
not not9828(N31182,in2);
not not9829(N31183,R3);
not not9830(N31194,in0);
not not9831(N31195,R1);
not not9832(N31207,in0);
not not9833(N31208,R0);
not not9834(N31209,R1);
not not9835(N31220,in0);
not not9836(N31221,R1);
not not9837(N31233,in0);
not not9838(N31234,in1);
not not9839(N31235,R2);
not not9840(N31246,in0);
not not9841(N31247,in1);
not not9842(N31248,in2);
not not9843(N31258,in0);
not not9844(N31259,in2);
not not9845(N31270,in0);
not not9846(N31282,in0);
not not9847(N31283,R2);
not not9848(N31294,in0);
not not9849(N31306,in0);
not not9850(N31307,in1);
not not9851(N31308,in2);
not not9852(N31318,in0);
not not9853(N31319,R0);
not not9854(N31330,in0);
not not9855(N31331,in1);
not not9856(N31342,in0);
not not9857(N31343,in2);
not not9858(N31354,in0);
not not9859(N31355,R3);
not not9860(N31366,in0);
not not9861(N31376,in0);
not not9862(N31386,in0);
not not9863(N31396,in0);
not not9864(N31406,in0);
not not9865(N31415,in0);
not not9866(N31416,in2);
not not9867(N31417,R0);
not not9868(N31418,R3);
not not9869(N31419,R4);
not not9870(N31420,R5);
not not9871(N31431,in0);
not not9872(N31432,in2);
not not9873(N31433,R0);
not not9874(N31434,R1);
not not9875(N31435,R2);
not not9876(N31436,R4);
not not9877(N31437,R5);
not not9878(N31447,in0);
not not9879(N31448,in1);
not not9880(N31449,R0);
not not9881(N31450,R1);
not not9882(N31451,R3);
not not9883(N31452,R4);
not not9884(N31463,in0);
not not9885(N31464,in2);
not not9886(N31465,R1);
not not9887(N31466,R4);
not not9888(N31467,R5);
not not9889(N31478,in0);
not not9890(N31479,in1);
not not9891(N31480,in2);
not not9892(N31481,R0);
not not9893(N31482,R2);
not not9894(N31493,in0);
not not9895(N31494,in1);
not not9896(N31495,R0);
not not9897(N31496,R2);
not not9898(N31497,R5);
not not9899(N31508,in0);
not not9900(N31509,in2);
not not9901(N31510,R2);
not not9902(N31511,R4);
not not9903(N31522,in0);
not not9904(N31523,in1);
not not9905(N31524,in2);
not not9906(N31525,R1);
not not9907(N31526,R4);
not not9908(N31536,in0);
not not9909(N31537,in2);
not not9910(N31538,R3);
not not9911(N31539,R5);
not not9912(N31550,in0);
not not9913(N31551,in2);
not not9914(N31552,R0);
not not9915(N31553,R4);
not not9916(N31554,R5);
not not9917(N31564,in0);
not not9918(N31565,R0);
not not9919(N31566,R1);
not not9920(N31567,R2);
not not9921(N31568,R4);
not not9922(N31578,in0);
not not9923(N31579,in1);
not not9924(N31580,R2);
not not9925(N31581,R3);
not not9926(N31592,in0);
not not9927(N31593,in1);
not not9928(N31594,R0);
not not9929(N31595,R4);
not not9930(N31605,in0);
not not9931(N31606,in1);
not not9932(N31607,R0);
not not9933(N31608,R4);
not not9934(N31609,R5);
not not9935(N31618,in0);
not not9936(N31619,in1);
not not9937(N31620,in2);
not not9938(N31621,R0);
not not9939(N31631,in0);
not not9940(N31632,in1);
not not9941(N31633,R0);
not not9942(N31634,R4);
not not9943(N31643,in0);
not not9944(N31644,in2);
not not9945(N31645,R4);
not not9946(N31655,in0);
not not9947(N31656,in1);
not not9948(N31657,R5);
not not9949(N31667,in0);
not not9950(N31668,in1);
not not9951(N31669,R2);
not not9952(N31679,in0);
not not9953(N31680,in1);
not not9954(N31681,R0);
not not9955(N31691,in0);
not not9956(N31692,in2);
not not9957(N31693,R0);
not not9958(N31702,in0);
not not9959(N31713,in0);
not not9960(N31724,in0);
not not9961(N31733,in0);
not not9962(N31734,in1);
not not9963(N31735,in2);
not not9964(N31736,R2);
not not9965(N31737,R5);
not not9966(N31738,R6);
not not9967(N31739,R7);
not not9968(N29448,R2);
not not9969(N29449,R3);
not not9970(N29450,R6);
not not9971(N29451,R7);
not not9972(N29465,R2);
not not9973(N29466,R3);
not not9974(N29467,R4);
not not9975(N29468,R6);
not not9976(N29469,R7);
not not9977(N29483,R2);
not not9978(N29484,R3);
not not9979(N29485,R4);
not not9980(N29486,R7);
not not9981(N29500,R2);
not not9982(N29501,R3);
not not9983(N29502,R4);
not not9984(N29503,R7);
not not9985(N29518,R4);
not not9986(N29519,R5);
not not9987(N29534,R5);
not not9988(N29535,R7);
not not9989(N29549,R4);
not not9990(N29565,R4);
not not9991(N29566,R5);
not not9992(N29567,R6);
not not9993(N29582,R3);
not not9994(N29583,R4);
not not9995(N29584,R5);
not not9996(N29585,R7);
not not9997(N29600,R3);
not not9998(N29601,R4);
not not9999(N29602,R5);
not not10000(N29603,R6);
not not10001(N29617,R4);
not not10002(N29618,R5);
not not10003(N29619,R6);
not not10004(N29620,R7);
not not10005(N29635,R4);
not not10006(N29636,R5);
not not10007(N29637,R6);
not not10008(N29652,R5);
not not10009(N29653,R6);
not not10010(N29654,R7);
not not10011(N29668,R3);
not not10012(N29669,R4);
not not10013(N29670,R5);
not not10014(N29671,R7);
not not10015(N29686,R4);
not not10016(N29687,R5);
not not10017(N29688,R7);
not not10018(N29703,R4);
not not10019(N29704,R5);
not not10020(N29705,R7);
not not10021(N29720,R6);
not not10022(N29721,R7);
not not10023(N29735,R4);
not not10024(N29736,R6);
not not10025(N29737,R7);
not not10026(N29751,R5);
not not10027(N29752,R6);
not not10028(N29753,R7);
not not10029(N29768,R6);
not not10030(N29769,R7);
not not10031(N29783,R4);
not not10032(N29784,R5);
not not10033(N29785,R6);
not not10034(N29798,R4);
not not10035(N29799,R5);
not not10036(N29800,R6);
not not10037(N29801,R7);
not not10038(N29816,R4);
not not10039(N29817,R6);
not not10040(N29832,R5);
not not10041(N29833,R6);
not not10042(N29847,R4);
not not10043(N29848,R6);
not not10044(N29849,R7);
not not10045(N29863,R5);
not not10046(N29864,R6);
not not10047(N29865,R7);
not not10048(N29880,R4);
not not10049(N29881,R7);
not not10050(N29896,R3);
not not10051(N29897,R7);
not not10052(N29911,R5);
not not10053(N29912,R6);
not not10054(N29913,R7);
not not10055(N29927,R3);
not not10056(N29928,R4);
not not10057(N29929,R5);
not not10058(N29944,R5);
not not10059(N29945,R6);
not not10060(N29959,R4);
not not10061(N29960,R6);
not not10062(N29961,R7);
not not10063(N29975,R4);
not not10064(N29976,R5);
not not10065(N29977,R7);
not not10066(N29991,R4);
not not10067(N29992,R5);
not not10068(N29993,R6);
not not10069(N30007,R4);
not not10070(N30008,R5);
not not10071(N30021,R3);
not not10072(N30022,R5);
not not10073(N30023,R6);
not not10074(N30036,R4);
not not10075(N30037,R5);
not not10076(N30038,R6);
not not10077(N30051,R4);
not not10078(N30052,R6);
not not10079(N30053,R7);
not not10080(N30066,R4);
not not10081(N30067,R5);
not not10082(N30068,R6);
not not10083(N30081,R5);
not not10084(N30082,R6);
not not10085(N30083,R7);
not not10086(N30098,R5);
not not10087(N30112,R6);
not not10088(N30113,R7);
not not10089(N30126,R5);
not not10090(N30127,R6);
not not10091(N30128,R7);
not not10092(N30140,R4);
not not10093(N30141,R5);
not not10094(N30142,R6);
not not10095(N30143,R7);
not not10096(N30156,R5);
not not10097(N30157,R6);
not not10098(N30158,R7);
not not10099(N30171,R3);
not not10100(N30172,R4);
not not10101(N30173,R6);
not not10102(N30186,R3);
not not10103(N30187,R5);
not not10104(N30188,R6);
not not10105(N30201,R4);
not not10106(N30202,R5);
not not10107(N30203,R7);
not not10108(N30216,R4);
not not10109(N30217,R6);
not not10110(N30218,R7);
not not10111(N30232,R3);
not not10112(N30233,R7);
not not10113(N30246,R3);
not not10114(N30247,R6);
not not10115(N30248,R7);
not not10116(N30261,R5);
not not10117(N30262,R6);
not not10118(N30263,R7);
not not10119(N30276,R5);
not not10120(N30277,R6);
not not10121(N30278,R7);
not not10122(N30292,R5);
not not10123(N30293,R6);
not not10124(N30307,R5);
not not10125(N30308,R6);
not not10126(N30322,R4);
not not10127(N30323,R5);
not not10128(N30336,R4);
not not10129(N30337,R5);
not not10130(N30338,R7);
not not10131(N30351,R4);
not not10132(N30352,R5);
not not10133(N30353,R6);
not not10134(N30367,R6);
not not10135(N30368,R7);
not not10136(N30381,R4);
not not10137(N30382,R5);
not not10138(N30383,R7);
not not10139(N30397,R5);
not not10140(N30398,R7);
not not10141(N30411,R4);
not not10142(N30412,R6);
not not10143(N30413,R7);
not not10144(N30426,R5);
not not10145(N30427,R6);
not not10146(N30428,R7);
not not10147(N30441,R4);
not not10148(N30442,R6);
not not10149(N30443,R7);
not not10150(N30456,R4);
not not10151(N30457,R5);
not not10152(N30458,R6);
not not10153(N30472,R5);
not not10154(N30473,R7);
not not10155(N30485,R5);
not not10156(N30486,R6);
not not10157(N30487,R7);
not not10158(N30500,R6);
not not10159(N30501,R7);
not not10160(N30514,R5);
not not10161(N30515,R7);
not not10162(N30528,R4);
not not10163(N30529,R5);
not not10164(N30542,R6);
not not10165(N30543,R7);
not not10166(N30557,R6);
not not10167(N30571,R6);
not not10168(N30584,R4);
not not10169(N30585,R7);
not not10170(N30598,R6);
not not10171(N30599,R7);
not not10172(N30612,R4);
not not10173(N30613,R6);
not not10174(N30626,R4);
not not10175(N30627,R5);
not not10176(N30640,R4);
not not10177(N30641,R5);
not not10178(N30654,R4);
not not10179(N30655,R6);
not not10180(N30669,R6);
not not10181(N30682,R5);
not not10182(N30683,R7);
not not10183(N30695,R4);
not not10184(N30696,R6);
not not10185(N30697,R7);
not not10186(N30710,R4);
not not10187(N30711,R7);
not not10188(N30725,R5);
not not10189(N30738,R4);
not not10190(N30739,R7);
not not10191(N30753,R5);
not not10192(N30767,R5);
not not10193(N30780,R5);
not not10194(N30781,R7);
not not10195(N30795,R3);
not not10196(N30808,R5);
not not10197(N30809,R6);
not not10198(N30822,R5);
not not10199(N30823,R6);
not not10200(N30835,R3);
not not10201(N30836,R4);
not not10202(N30837,R7);
not not10203(N30850,R5);
not not10204(N30851,R6);
not not10205(N30865,R7);
not not10206(N30879,R6);
not not10207(N30893,R5);
not not10208(N30906,R5);
not not10209(N30907,R6);
not not10210(N30920,R5);
not not10211(N30921,R6);
not not10212(N30934,R3);
not not10213(N30935,R5);
not not10214(N30948,R3);
not not10215(N30949,R6);
not not10216(N30962,R4);
not not10217(N30963,R5);
not not10218(N30976,R5);
not not10219(N30987,R4);
not not10220(N30988,R5);
not not10221(N30989,R6);
not not10222(N31002,R7);
not not10223(N31014,R6);
not not10224(N31015,R7);
not not10225(N31026,R4);
not not10226(N31027,R5);
not not10227(N31028,R6);
not not10228(N31040,R4);
not not10229(N31041,R6);
not not10230(N31053,R3);
not not10231(N31054,R7);
not not10232(N31067,R4);
not not10233(N31080,R7);
not not10234(N31093,R5);
not not10235(N31106,R6);
not not10236(N31118,R4);
not not10237(N31119,R5);
not not10238(N31132,R5);
not not10239(N31144,R3);
not not10240(N31145,R7);
not not10241(N31157,R3);
not not10242(N31158,R6);
not not10243(N31171,R5);
not not10244(N31184,R5);
not not10245(N31196,R5);
not not10246(N31197,R6);
not not10247(N31210,R7);
not not10248(N31222,R3);
not not10249(N31223,R6);
not not10250(N31236,R4);
not not10251(N31260,R4);
not not10252(N31271,R4);
not not10253(N31272,R5);
not not10254(N31284,R5);
not not10255(N31295,R4);
not not10256(N31296,R5);
not not10257(N31320,R6);
not not10258(N31332,R5);
not not10259(N31344,R5);
not not10260(N31356,R5);
not not10261(N31421,R6);
not not10262(N31422,R7);
not not10263(N31438,R7);
not not10264(N31453,R6);
not not10265(N31454,R7);
not not10266(N31468,R6);
not not10267(N31469,R7);
not not10268(N31483,R6);
not not10269(N31484,R7);
not not10270(N31498,R6);
not not10271(N31499,R7);
not not10272(N31512,R5);
not not10273(N31513,R7);
not not10274(N31527,R5);
not not10275(N31540,R6);
not not10276(N31541,R7);
not not10277(N31555,R7);
not not10278(N31569,R6);
not not10279(N31582,R5);
not not10280(N31583,R6);
not not10281(N31596,R5);
not not10282(N31622,R6);
not not10283(N31646,R7);
not not10284(N31658,R7);
not not10285(N31670,R6);
not not10286(N31682,R7);
not not10287(N31703,R6);
not not10288(N31704,R7);
not not10289(N31714,R6);
not not10290(N31715,R7);
not not10291(N31725,R7);
not not10292(N31922,in0);
not not10293(N31923,in1);
not not10294(N31924,in2);
not not10295(N31925,R0);
not not10296(N31926,R1);
not not10297(N31939,in0);
not not10298(N31940,in2);
not not10299(N31941,R1);
not not10300(N31955,in0);
not not10301(N31956,R0);
not not10302(N31970,in0);
not not10303(N31971,R0);
not not10304(N31972,R1);
not not10305(N31984,in0);
not not10306(N31985,in2);
not not10307(N31986,R0);
not not10308(N31987,R2);
not not10309(N31988,R3);
not not10310(N32002,in0);
not not10311(N32003,in1);
not not10312(N32004,in2);
not not10313(N32005,R0);
not not10314(N32006,R1);
not not10315(N32007,R2);
not not10316(N32020,in0);
not not10317(N32021,in1);
not not10318(N32022,R0);
not not10319(N32023,R1);
not not10320(N32024,R2);
not not10321(N32038,in0);
not not10322(N32039,in2);
not not10323(N32040,R0);
not not10324(N32041,R1);
not not10325(N32042,R2);
not not10326(N32043,R3);
not not10327(N32055,in0);
not not10328(N32056,in2);
not not10329(N32057,R0);
not not10330(N32058,R1);
not not10331(N32059,R2);
not not10332(N32072,in0);
not not10333(N32073,in1);
not not10334(N32074,in2);
not not10335(N32075,R3);
not not10336(N32089,in0);
not not10337(N32090,in1);
not not10338(N32091,in2);
not not10339(N32092,R1);
not not10340(N32106,in0);
not not10341(N32107,in1);
not not10342(N32108,in2);
not not10343(N32109,R1);
not not10344(N32110,R2);
not not10345(N32123,in0);
not not10346(N32124,R0);
not not10347(N32125,R1);
not not10348(N32126,R2);
not not10349(N32140,in0);
not not10350(N32141,in1);
not not10351(N32142,in2);
not not10352(N32143,R0);
not not10353(N32144,R2);
not not10354(N32157,in0);
not not10355(N32158,in1);
not not10356(N32159,in2);
not not10357(N32160,R1);
not not10358(N32161,R2);
not not10359(N32174,in0);
not not10360(N32175,in1);
not not10361(N32176,in2);
not not10362(N32177,R1);
not not10363(N32178,R3);
not not10364(N32191,in0);
not not10365(N32192,in1);
not not10366(N32193,in2);
not not10367(N32194,R0);
not not10368(N32195,R1);
not not10369(N32196,R2);
not not10370(N32208,in0);
not not10371(N32209,in1);
not not10372(N32210,R1);
not not10373(N32211,R2);
not not10374(N32225,in0);
not not10375(N32226,in2);
not not10376(N32227,R1);
not not10377(N32228,R2);
not not10378(N32242,in0);
not not10379(N32243,in2);
not not10380(N32244,R0);
not not10381(N32245,R2);
not not10382(N32259,in0);
not not10383(N32260,in1);
not not10384(N32261,R0);
not not10385(N32262,R2);
not not10386(N32275,in0);
not not10387(N32276,in2);
not not10388(N32277,R0);
not not10389(N32278,R2);
not not10390(N32291,in0);
not not10391(N32292,in2);
not not10392(N32293,R0);
not not10393(N32294,R2);
not not10394(N32307,in0);
not not10395(N32308,in1);
not not10396(N32309,R1);
not not10397(N32310,R3);
not not10398(N32323,in0);
not not10399(N32324,in2);
not not10400(N32325,R0);
not not10401(N32326,R1);
not not10402(N32339,in0);
not not10403(N32340,R0);
not not10404(N32341,R1);
not not10405(N32355,in0);
not not10406(N32356,in2);
not not10407(N32357,R0);
not not10408(N32358,R1);
not not10409(N32359,R2);
not not10410(N32371,in0);
not not10411(N32372,in2);
not not10412(N32373,R0);
not not10413(N32374,R1);
not not10414(N32375,R2);
not not10415(N32387,in0);
not not10416(N32388,R0);
not not10417(N32389,R1);
not not10418(N32390,R3);
not not10419(N32403,in0);
not not10420(N32404,in2);
not not10421(N32405,R0);
not not10422(N32406,R3);
not not10423(N32419,in0);
not not10424(N32420,in1);
not not10425(N32421,in2);
not not10426(N32422,R2);
not not10427(N32423,R3);
not not10428(N32435,in0);
not not10429(N32436,in1);
not not10430(N32437,in2);
not not10431(N32438,R0);
not not10432(N32439,R2);
not not10433(N32451,in0);
not not10434(N32452,R1);
not not10435(N32453,R2);
not not10436(N32454,R3);
not not10437(N32467,in0);
not not10438(N32468,in1);
not not10439(N32469,R2);
not not10440(N32470,R3);
not not10441(N32483,in0);
not not10442(N32484,in1);
not not10443(N32485,R0);
not not10444(N32486,R3);
not not10445(N32499,in0);
not not10446(N32500,R0);
not not10447(N32501,R1);
not not10448(N32502,R2);
not not10449(N32515,in0);
not not10450(N32516,in2);
not not10451(N32517,R0);
not not10452(N32518,R2);
not not10453(N32531,in0);
not not10454(N32532,in1);
not not10455(N32533,in2);
not not10456(N32534,R2);
not not10457(N32547,in0);
not not10458(N32548,R1);
not not10459(N32549,R2);
not not10460(N32563,in0);
not not10461(N32564,in1);
not not10462(N32565,R0);
not not10463(N32566,R1);
not not10464(N32567,R3);
not not10465(N32579,in0);
not not10466(N32580,in2);
not not10467(N32581,R0);
not not10468(N32582,R1);
not not10469(N32583,R3);
not not10470(N32595,in0);
not not10471(N32596,in1);
not not10472(N32597,R0);
not not10473(N32598,R1);
not not10474(N32611,in0);
not not10475(N32612,R0);
not not10476(N32613,R1);
not not10477(N32614,R2);
not not10478(N32626,in0);
not not10479(N32627,R1);
not not10480(N32628,R2);
not not10481(N32641,in0);
not not10482(N32642,in2);
not not10483(N32643,R1);
not not10484(N32644,R2);
not not10485(N32656,in0);
not not10486(N32657,in1);
not not10487(N32658,R0);
not not10488(N32659,R2);
not not10489(N32671,in0);
not not10490(N32672,in1);
not not10491(N32673,R1);
not not10492(N32686,in0);
not not10493(N32687,in1);
not not10494(N32688,R0);
not not10495(N32689,R1);
not not10496(N32701,in0);
not not10497(N32702,in2);
not not10498(N32703,R1);
not not10499(N32704,R2);
not not10500(N32716,in0);
not not10501(N32717,in2);
not not10502(N32718,R0);
not not10503(N32719,R2);
not not10504(N32731,in0);
not not10505(N32732,in2);
not not10506(N32733,R2);
not not10507(N32746,in0);
not not10508(N32747,in1);
not not10509(N32748,R0);
not not10510(N32749,R3);
not not10511(N32761,in0);
not not10512(N32762,R0);
not not10513(N32763,R2);
not not10514(N32776,in0);
not not10515(N32777,in2);
not not10516(N32778,R2);
not not10517(N32791,in0);
not not10518(N32792,in1);
not not10519(N32793,R0);
not not10520(N32806,in0);
not not10521(N32807,in1);
not not10522(N32808,in2);
not not10523(N32809,R2);
not not10524(N32821,in0);
not not10525(N32822,in1);
not not10526(N32823,in2);
not not10527(N32824,R3);
not not10528(N32836,in0);
not not10529(N32837,in1);
not not10530(N32838,R0);
not not10531(N32839,R2);
not not10532(N32840,R3);
not not10533(N32851,in0);
not not10534(N32852,R1);
not not10535(N32853,R3);
not not10536(N32866,in0);
not not10537(N32867,in1);
not not10538(N32868,R0);
not not10539(N32869,R2);
not not10540(N32881,in0);
not not10541(N32882,in1);
not not10542(N32883,R0);
not not10543(N32884,R1);
not not10544(N32896,in0);
not not10545(N32897,in2);
not not10546(N32898,R1);
not not10547(N32899,R2);
not not10548(N32911,in0);
not not10549(N32912,in1);
not not10550(N32913,in2);
not not10551(N32914,R1);
not not10552(N32926,in0);
not not10553(N32927,R0);
not not10554(N32928,R2);
not not10555(N32941,in0);
not not10556(N32942,in2);
not not10557(N32943,R1);
not not10558(N32944,R2);
not not10559(N32956,in0);
not not10560(N32957,in1);
not not10561(N32958,R2);
not not10562(N32959,R3);
not not10563(N32971,in0);
not not10564(N32972,in1);
not not10565(N32973,in2);
not not10566(N32974,R3);
not not10567(N32986,in0);
not not10568(N32987,in1);
not not10569(N32988,R0);
not not10570(N32989,R2);
not not10571(N32990,R3);
not not10572(N33001,in0);
not not10573(N33002,in1);
not not10574(N33003,in2);
not not10575(N33016,in0);
not not10576(N33017,in1);
not not10577(N33018,in2);
not not10578(N33031,in0);
not not10579(N33032,in1);
not not10580(N33033,in2);
not not10581(N33034,R2);
not not10582(N33046,in0);
not not10583(N33047,in1);
not not10584(N33048,in2);
not not10585(N33049,R2);
not not10586(N33061,in0);
not not10587(N33062,in2);
not not10588(N33063,R0);
not not10589(N33076,in0);
not not10590(N33077,in1);
not not10591(N33078,R2);
not not10592(N33079,R3);
not not10593(N33091,in0);
not not10594(N33092,in2);
not not10595(N33093,R1);
not not10596(N33094,R2);
not not10597(N33106,in0);
not not10598(N33107,R0);
not not10599(N33108,R1);
not not10600(N33109,R2);
not not10601(N33121,in0);
not not10602(N33122,in2);
not not10603(N33123,R2);
not not10604(N33124,R3);
not not10605(N33136,in0);
not not10606(N33137,R2);
not not10607(N33138,R3);
not not10608(N33150,in0);
not not10609(N33151,R2);
not not10610(N33164,in0);
not not10611(N33165,in1);
not not10612(N33166,R2);
not not10613(N33178,in0);
not not10614(N33179,in1);
not not10615(N33180,R1);
not not10616(N33181,R2);
not not10617(N33192,in0);
not not10618(N33193,in2);
not not10619(N33194,R0);
not not10620(N33195,R2);
not not10621(N33206,in0);
not not10622(N33207,in2);
not not10623(N33208,R0);
not not10624(N33220,in0);
not not10625(N33221,in1);
not not10626(N33222,R2);
not not10627(N33234,in0);
not not10628(N33235,R2);
not not10629(N33248,in0);
not not10630(N33249,R0);
not not10631(N33250,R2);
not not10632(N33262,in0);
not not10633(N33263,in2);
not not10634(N33264,R0);
not not10635(N33265,R2);
not not10636(N33276,in0);
not not10637(N33277,in2);
not not10638(N33278,R1);
not not10639(N33279,R2);
not not10640(N33290,in0);
not not10641(N33291,R0);
not not10642(N33304,in0);
not not10643(N33305,in1);
not not10644(N33306,in2);
not not10645(N33307,R2);
not not10646(N33318,in0);
not not10647(N33319,in1);
not not10648(N33320,in2);
not not10649(N33332,in0);
not not10650(N33333,in1);
not not10651(N33334,R0);
not not10652(N33346,in0);
not not10653(N33347,R2);
not not10654(N33348,R3);
not not10655(N33360,in0);
not not10656(N33361,R2);
not not10657(N33362,R3);
not not10658(N33374,in0);
not not10659(N33375,in2);
not not10660(N33376,R0);
not not10661(N33377,R2);
not not10662(N33388,in0);
not not10663(N33389,in1);
not not10664(N33402,in0);
not not10665(N33403,in1);
not not10666(N33404,R2);
not not10667(N33416,in0);
not not10668(N33417,in1);
not not10669(N33418,in2);
not not10670(N33419,R2);
not not10671(N33430,in0);
not not10672(N33431,in1);
not not10673(N33432,R1);
not not10674(N33433,R3);
not not10675(N33444,in0);
not not10676(N33445,in1);
not not10677(N33446,R0);
not not10678(N33447,R1);
not not10679(N33458,in0);
not not10680(N33459,R0);
not not10681(N33460,R1);
not not10682(N33472,in0);
not not10683(N33473,R0);
not not10684(N33486,in0);
not not10685(N33487,in1);
not not10686(N33488,R1);
not not10687(N33500,in0);
not not10688(N33501,R0);
not not10689(N33502,R1);
not not10690(N33514,in0);
not not10691(N33515,in1);
not not10692(N33516,R2);
not not10693(N33528,in0);
not not10694(N33529,in1);
not not10695(N33542,in0);
not not10696(N33543,in1);
not not10697(N33544,R1);
not not10698(N33545,R2);
not not10699(N33556,in0);
not not10700(N33557,in1);
not not10701(N33558,in2);
not not10702(N33559,R0);
not not10703(N33570,in0);
not not10704(N33571,in2);
not not10705(N33572,R1);
not not10706(N33584,in0);
not not10707(N33585,R0);
not not10708(N33586,R1);
not not10709(N33587,R3);
not not10710(N33598,in0);
not not10711(N33599,in1);
not not10712(N33600,in2);
not not10713(N33601,R2);
not not10714(N33611,in0);
not not10715(N33612,in1);
not not10716(N33613,in2);
not not10717(N33624,in0);
not not10718(N33625,in2);
not not10719(N33637,in0);
not not10720(N33638,R2);
not not10721(N33650,in0);
not not10722(N33651,R1);
not not10723(N33663,in0);
not not10724(N33664,R2);
not not10725(N33676,in0);
not not10726(N33677,R1);
not not10727(N33689,in0);
not not10728(N33690,in1);
not not10729(N33691,R1);
not not10730(N33702,in0);
not not10731(N33703,in2);
not not10732(N33715,in0);
not not10733(N33716,in1);
not not10734(N33717,in2);
not not10735(N33718,R1);
not not10736(N33728,in0);
not not10737(N33729,in1);
not not10738(N33730,in2);
not not10739(N33731,R2);
not not10740(N33741,in0);
not not10741(N33742,R1);
not not10742(N33743,R3);
not not10743(N33754,in0);
not not10744(N33755,in2);
not not10745(N33756,R0);
not not10746(N33767,in0);
not not10747(N33768,R0);
not not10748(N33769,R2);
not not10749(N33780,in0);
not not10750(N33781,in2);
not not10751(N33782,R3);
not not10752(N33793,in0);
not not10753(N33806,in0);
not not10754(N33807,R2);
not not10755(N33819,in0);
not not10756(N33820,R0);
not not10757(N33821,R2);
not not10758(N33832,in0);
not not10759(N33833,in1);
not not10760(N33845,in0);
not not10761(N33846,R2);
not not10762(N33858,in0);
not not10763(N33859,R2);
not not10764(N33871,in0);
not not10765(N33872,in1);
not not10766(N33883,in0);
not not10767(N33884,in2);
not not10768(N33895,in0);
not not10769(N33896,in1);
not not10770(N33897,R3);
not not10771(N33907,in0);
not not10772(N33908,in2);
not not10773(N33909,R0);
not not10774(N33919,in0);
not not10775(N33920,R0);
not not10776(N33931,in0);
not not10777(N33943,in0);
not not10778(N33944,R0);
not not10779(N33945,R1);
not not10780(N33955,in0);
not not10781(N33967,in0);
not not10782(N33979,in0);
not not10783(N33980,R1);
not not10784(N33991,in0);
not not10785(N33992,R0);
not not10786(N34003,in0);
not not10787(N34004,R3);
not not10788(N34015,in0);
not not10789(N34016,R1);
not not10790(N34027,in0);
not not10791(N34039,in0);
not not10792(N34051,in0);
not not10793(N34062,in0);
not not10794(N34063,R1);
not not10795(N34072,in0);
not not10796(N34073,in1);
not not10797(N34074,R0);
not not10798(N34075,R1);
not not10799(N34076,R3);
not not10800(N34077,R4);
not not10801(N34088,in0);
not not10802(N34089,in2);
not not10803(N34090,R0);
not not10804(N34091,R3);
not not10805(N34092,R5);
not not10806(N34103,in0);
not not10807(N34104,in1);
not not10808(N34105,R0);
not not10809(N34106,R1);
not not10810(N34107,R2);
not not10811(N34108,R5);
not not10812(N34118,in0);
not not10813(N34119,in2);
not not10814(N34120,R1);
not not10815(N34121,R3);
not not10816(N34122,R5);
not not10817(N34133,in0);
not not10818(N34134,in1);
not not10819(N34135,R0);
not not10820(N34136,R1);
not not10821(N34137,R5);
not not10822(N34148,in0);
not not10823(N34149,in1);
not not10824(N34150,in2);
not not10825(N34151,R0);
not not10826(N34152,R2);
not not10827(N34162,in0);
not not10828(N34163,in1);
not not10829(N34164,in2);
not not10830(N34165,R3);
not not10831(N34176,in0);
not not10832(N34177,in1);
not not10833(N34178,R0);
not not10834(N34179,R2);
not not10835(N34180,R4);
not not10836(N34190,in0);
not not10837(N34191,R0);
not not10838(N34192,R1);
not not10839(N34193,R2);
not not10840(N34194,R5);
not not10841(N34204,in0);
not not10842(N34205,in2);
not not10843(N34206,R0);
not not10844(N34207,R1);
not not10845(N34208,R4);
not not10846(N34218,in0);
not not10847(N34219,in1);
not not10848(N34220,in2);
not not10849(N34221,R4);
not not10850(N34232,in0);
not not10851(N34233,in1);
not not10852(N34234,R0);
not not10853(N34235,R2);
not not10854(N34236,R5);
not not10855(N34246,in0);
not not10856(N34247,R3);
not not10857(N34248,R5);
not not10858(N34259,in0);
not not10859(N34260,R1);
not not10860(N34261,R3);
not not10861(N34262,R4);
not not10862(N34272,in0);
not not10863(N34273,in1);
not not10864(N34274,R3);
not not10865(N34285,in0);
not not10866(N34286,in1);
not not10867(N34287,R4);
not not10868(N34298,in0);
not not10869(N34299,in2);
not not10870(N34300,R0);
not not10871(N34310,in0);
not not10872(N34311,in2);
not not10873(N34312,R5);
not not10874(N34322,in0);
not not10875(N34323,R1);
not not10876(N34334,in0);
not not10877(N34345,in0);
not not10878(N34346,in2);
not not10879(N34356,in0);
not not10880(N34357,in1);
not not10881(N34367,in0);
not not10882(N34368,in1);
not not10883(N34369,R2);
not not10884(N34378,in0);
not not10885(N34389,in0);
not not10886(N34390,in2);
not not10887(N31927,R5);
not not10888(N31928,R7);
not not10889(N31942,R3);
not not10890(N31943,R4);
not not10891(N31944,R5);
not not10892(N31957,R3);
not not10893(N31958,R5);
not not10894(N31959,R6);
not not10895(N31973,R3);
not not10896(N31974,R6);
not not10897(N31989,R4);
not not10898(N31990,R5);
not not10899(N31991,R6);
not not10900(N31992,R7);
not not10901(N32008,R4);
not not10902(N32009,R5);
not not10903(N32010,R6);
not not10904(N32025,R3);
not not10905(N32026,R4);
not not10906(N32027,R5);
not not10907(N32028,R6);
not not10908(N32044,R6);
not not10909(N32045,R7);
not not10910(N32060,R3);
not not10911(N32061,R5);
not not10912(N32062,R6);
not not10913(N32076,R4);
not not10914(N32077,R5);
not not10915(N32078,R6);
not not10916(N32079,R7);
not not10917(N32093,R4);
not not10918(N32094,R5);
not not10919(N32095,R6);
not not10920(N32096,R7);
not not10921(N32111,R4);
not not10922(N32112,R5);
not not10923(N32113,R7);
not not10924(N32127,R3);
not not10925(N32128,R4);
not not10926(N32129,R5);
not not10927(N32130,R7);
not not10928(N32145,R3);
not not10929(N32146,R4);
not not10930(N32147,R5);
not not10931(N32162,R4);
not not10932(N32163,R6);
not not10933(N32164,R7);
not not10934(N32179,R4);
not not10935(N32180,R5);
not not10936(N32181,R7);
not not10937(N32197,R6);
not not10938(N32198,R7);
not not10939(N32212,R3);
not not10940(N32213,R4);
not not10941(N32214,R5);
not not10942(N32215,R7);
not not10943(N32229,R4);
not not10944(N32230,R5);
not not10945(N32231,R6);
not not10946(N32232,R7);
not not10947(N32246,R3);
not not10948(N32247,R4);
not not10949(N32248,R6);
not not10950(N32249,R7);
not not10951(N32263,R4);
not not10952(N32264,R5);
not not10953(N32265,R7);
not not10954(N32279,R4);
not not10955(N32280,R5);
not not10956(N32281,R6);
not not10957(N32295,R5);
not not10958(N32296,R6);
not not10959(N32297,R7);
not not10960(N32311,R4);
not not10961(N32312,R5);
not not10962(N32313,R6);
not not10963(N32327,R4);
not not10964(N32328,R5);
not not10965(N32329,R6);
not not10966(N32342,R4);
not not10967(N32343,R5);
not not10968(N32344,R6);
not not10969(N32345,R7);
not not10970(N32360,R4);
not not10971(N32361,R6);
not not10972(N32376,R4);
not not10973(N32377,R5);
not not10974(N32391,R4);
not not10975(N32392,R5);
not not10976(N32393,R7);
not not10977(N32407,R4);
not not10978(N32408,R5);
not not10979(N32409,R7);
not not10980(N32424,R5);
not not10981(N32425,R6);
not not10982(N32440,R5);
not not10983(N32441,R6);
not not10984(N32455,R4);
not not10985(N32456,R5);
not not10986(N32457,R6);
not not10987(N32471,R5);
not not10988(N32472,R6);
not not10989(N32473,R7);
not not10990(N32487,R4);
not not10991(N32488,R5);
not not10992(N32489,R6);
not not10993(N32503,R5);
not not10994(N32504,R6);
not not10995(N32505,R7);
not not10996(N32519,R4);
not not10997(N32520,R5);
not not10998(N32521,R6);
not not10999(N32535,R3);
not not11000(N32536,R4);
not not11001(N32537,R7);
not not11002(N32550,R3);
not not11003(N32551,R4);
not not11004(N32552,R6);
not not11005(N32553,R7);
not not11006(N32568,R5);
not not11007(N32569,R6);
not not11008(N32584,R6);
not not11009(N32585,R7);
not not11010(N32599,R3);
not not11011(N32600,R4);
not not11012(N32601,R6);
not not11013(N32615,R5);
not not11014(N32616,R6);
not not11015(N32629,R4);
not not11016(N32630,R6);
not not11017(N32631,R7);
not not11018(N32645,R6);
not not11019(N32646,R7);
not not11020(N32660,R6);
not not11021(N32661,R7);
not not11022(N32674,R4);
not not11023(N32675,R5);
not not11024(N32676,R7);
not not11025(N32690,R6);
not not11026(N32691,R7);
not not11027(N32705,R6);
not not11028(N32706,R7);
not not11029(N32720,R4);
not not11030(N32721,R5);
not not11031(N32734,R4);
not not11032(N32735,R5);
not not11033(N32736,R6);
not not11034(N32750,R6);
not not11035(N32751,R7);
not not11036(N32764,R4);
not not11037(N32765,R5);
not not11038(N32766,R7);
not not11039(N32779,R3);
not not11040(N32780,R6);
not not11041(N32781,R7);
not not11042(N32794,R3);
not not11043(N32795,R5);
not not11044(N32796,R7);
not not11045(N32810,R3);
not not11046(N32811,R6);
not not11047(N32825,R4);
not not11048(N32826,R7);
not not11049(N32841,R7);
not not11050(N32854,R4);
not not11051(N32855,R5);
not not11052(N32856,R7);
not not11053(N32870,R4);
not not11054(N32871,R5);
not not11055(N32885,R6);
not not11056(N32886,R7);
not not11057(N32900,R5);
not not11058(N32901,R7);
not not11059(N32915,R4);
not not11060(N32916,R7);
not not11061(N32929,R3);
not not11062(N32930,R5);
not not11063(N32931,R7);
not not11064(N32945,R5);
not not11065(N32946,R6);
not not11066(N32960,R5);
not not11067(N32961,R6);
not not11068(N32975,R4);
not not11069(N32976,R5);
not not11070(N32991,R6);
not not11071(N33004,R4);
not not11072(N33005,R5);
not not11073(N33006,R6);
not not11074(N33019,R3);
not not11075(N33020,R5);
not not11076(N33021,R6);
not not11077(N33035,R6);
not not11078(N33036,R7);
not not11079(N33050,R6);
not not11080(N33051,R7);
not not11081(N33064,R4);
not not11082(N33065,R6);
not not11083(N33066,R7);
not not11084(N33080,R4);
not not11085(N33081,R6);
not not11086(N33095,R4);
not not11087(N33096,R5);
not not11088(N33110,R5);
not not11089(N33111,R7);
not not11090(N33125,R4);
not not11091(N33126,R5);
not not11092(N33139,R4);
not not11093(N33140,R7);
not not11094(N33152,R4);
not not11095(N33153,R5);
not not11096(N33154,R7);
not not11097(N33167,R5);
not not11098(N33168,R6);
not not11099(N33182,R6);
not not11100(N33196,R5);
not not11101(N33209,R5);
not not11102(N33210,R7);
not not11103(N33223,R4);
not not11104(N33224,R5);
not not11105(N33236,R4);
not not11106(N33237,R5);
not not11107(N33238,R7);
not not11108(N33251,R4);
not not11109(N33252,R5);
not not11110(N33266,R5);
not not11111(N33280,R7);
not not11112(N33292,R4);
not not11113(N33293,R5);
not not11114(N33294,R7);
not not11115(N33308,R5);
not not11116(N33321,R4);
not not11117(N33322,R7);
not not11118(N33335,R3);
not not11119(N33336,R7);
not not11120(N33349,R4);
not not11121(N33350,R7);
not not11122(N33363,R6);
not not11123(N33364,R7);
not not11124(N33378,R5);
not not11125(N33390,R4);
not not11126(N33391,R6);
not not11127(N33392,R7);
not not11128(N33405,R3);
not not11129(N33406,R5);
not not11130(N33420,R5);
not not11131(N33434,R5);
not not11132(N33448,R5);
not not11133(N33461,R4);
not not11134(N33462,R5);
not not11135(N33474,R4);
not not11136(N33475,R5);
not not11137(N33476,R7);
not not11138(N33489,R5);
not not11139(N33490,R6);
not not11140(N33503,R4);
not not11141(N33504,R5);
not not11142(N33517,R6);
not not11143(N33518,R7);
not not11144(N33530,R4);
not not11145(N33531,R5);
not not11146(N33532,R6);
not not11147(N33546,R7);
not not11148(N33560,R7);
not not11149(N33573,R5);
not not11150(N33574,R6);
not not11151(N33588,R5);
not not11152(N33614,R4);
not not11153(N33626,R4);
not not11154(N33627,R5);
not not11155(N33639,R5);
not not11156(N33640,R6);
not not11157(N33652,R4);
not not11158(N33653,R7);
not not11159(N33665,R4);
not not11160(N33666,R6);
not not11161(N33678,R4);
not not11162(N33679,R7);
not not11163(N33692,R7);
not not11164(N33704,R4);
not not11165(N33705,R5);
not not11166(N33744,R7);
not not11167(N33757,R4);
not not11168(N33770,R6);
not not11169(N33783,R6);
not not11170(N33794,R3);
not not11171(N33795,R4);
not not11172(N33796,R5);
not not11173(N33808,R5);
not not11174(N33809,R6);
not not11175(N33822,R5);
not not11176(N33834,R4);
not not11177(N33835,R7);
not not11178(N33847,R3);
not not11179(N33848,R7);
not not11180(N33860,R5);
not not11181(N33861,R7);
not not11182(N33873,R3);
not not11183(N33885,R5);
not not11184(N33921,R4);
not not11185(N33932,R3);
not not11186(N33933,R4);
not not11187(N33956,R6);
not not11188(N33957,R7);
not not11189(N33968,R4);
not not11190(N33969,R5);
not not11191(N33981,R5);
not not11192(N33993,R7);
not not11193(N34005,R4);
not not11194(N34017,R5);
not not11195(N34028,R6);
not not11196(N34029,R7);
not not11197(N34040,R3);
not not11198(N34041,R5);
not not11199(N34052,R6);
not not11200(N34078,R6);
not not11201(N34079,R7);
not not11202(N34093,R6);
not not11203(N34094,R7);
not not11204(N34109,R7);
not not11205(N34123,R6);
not not11206(N34124,R7);
not not11207(N34138,R6);
not not11208(N34139,R7);
not not11209(N34153,R4);
not not11210(N34166,R5);
not not11211(N34167,R7);
not not11212(N34181,R7);
not not11213(N34195,R6);
not not11214(N34209,R7);
not not11215(N34222,R6);
not not11216(N34223,R7);
not not11217(N34237,R7);
not not11218(N34249,R6);
not not11219(N34250,R7);
not not11220(N34263,R6);
not not11221(N34275,R5);
not not11222(N34276,R7);
not not11223(N34288,R6);
not not11224(N34289,R7);
not not11225(N34301,R6);
not not11226(N34313,R7);
not not11227(N34324,R5);
not not11228(N34325,R6);
not not11229(N34335,R6);
not not11230(N34336,R7);
not not11231(N34347,R7);
not not11232(N34358,R6);
not not11233(N34379,R6);
not not11234(N34380,R7);
not not11235(N34391,R5);
not not11236(N34592,in0);
not not11237(N34593,in1);
not not11238(N34594,in2);
not not11239(N34595,R0);
not not11240(N34612,in0);
not not11241(N34613,in1);
not not11242(N34614,R0);
not not11243(N34630,in0);
not not11244(N34631,in1);
not not11245(N34632,in2);
not not11246(N34633,R0);
not not11247(N34634,R1);
not not11248(N34646,in0);
not not11249(N34647,in2);
not not11250(N34648,R0);
not not11251(N34649,R1);
not not11252(N34650,R2);
not not11253(N34651,R3);
not not11254(N34664,in0);
not not11255(N34665,in1);
not not11256(N34666,R0);
not not11257(N34667,R1);
not not11258(N34668,R2);
not not11259(N34682,in0);
not not11260(N34683,in2);
not not11261(N34684,R0);
not not11262(N34685,R1);
not not11263(N34686,R2);
not not11264(N34700,in0);
not not11265(N34701,in1);
not not11266(N34702,in2);
not not11267(N34703,R0);
not not11268(N34704,R1);
not not11269(N34705,R3);
not not11270(N34718,in0);
not not11271(N34719,in1);
not not11272(N34720,in2);
not not11273(N34721,R0);
not not11274(N34722,R1);
not not11275(N34736,in0);
not not11276(N34737,in1);
not not11277(N34738,in2);
not not11278(N34739,R1);
not not11279(N34740,R2);
not not11280(N34753,in0);
not not11281(N34754,in1);
not not11282(N34755,R1);
not not11283(N34756,R2);
not not11284(N34757,R3);
not not11285(N34770,in0);
not not11286(N34771,in1);
not not11287(N34772,R1);
not not11288(N34773,R2);
not not11289(N34787,in0);
not not11290(N34788,in1);
not not11291(N34789,R0);
not not11292(N34790,R2);
not not11293(N34791,R3);
not not11294(N34803,in0);
not not11295(N34804,in2);
not not11296(N34805,R2);
not not11297(N34819,in0);
not not11298(N34820,in1);
not not11299(N34821,R1);
not not11300(N34822,R3);
not not11301(N34835,in0);
not not11302(N34836,in2);
not not11303(N34837,R0);
not not11304(N34838,R3);
not not11305(N34851,in0);
not not11306(N34852,in2);
not not11307(N34853,R1);
not not11308(N34854,R3);
not not11309(N34867,in0);
not not11310(N34868,in1);
not not11311(N34869,R0);
not not11312(N34870,R2);
not not11313(N34883,in0);
not not11314(N34884,in2);
not not11315(N34885,R0);
not not11316(N34886,R2);
not not11317(N34899,in0);
not not11318(N34900,R0);
not not11319(N34901,R1);
not not11320(N34902,R3);
not not11321(N34915,in0);
not not11322(N34916,in1);
not not11323(N34917,R1);
not not11324(N34918,R2);
not not11325(N34931,in0);
not not11326(N34932,in1);
not not11327(N34933,in2);
not not11328(N34934,R0);
not not11329(N34935,R2);
not not11330(N34947,in0);
not not11331(N34948,in1);
not not11332(N34949,in2);
not not11333(N34950,R0);
not not11334(N34951,R3);
not not11335(N34963,in0);
not not11336(N34964,in2);
not not11337(N34965,R1);
not not11338(N34966,R2);
not not11339(N34979,in0);
not not11340(N34980,in1);
not not11341(N34981,R1);
not not11342(N34982,R3);
not not11343(N34995,in0);
not not11344(N34996,R1);
not not11345(N34997,R2);
not not11346(N34998,R3);
not not11347(N35011,in0);
not not11348(N35012,in1);
not not11349(N35013,R0);
not not11350(N35014,R1);
not not11351(N35015,R2);
not not11352(N35027,in0);
not not11353(N35028,in1);
not not11354(N35029,R0);
not not11355(N35030,R1);
not not11356(N35031,R2);
not not11357(N35043,in0);
not not11358(N35044,R0);
not not11359(N35045,R1);
not not11360(N35046,R2);
not not11361(N35047,R3);
not not11362(N35059,in0);
not not11363(N35060,in2);
not not11364(N35061,R0);
not not11365(N35062,R1);
not not11366(N35063,R2);
not not11367(N35075,in0);
not not11368(N35076,R1);
not not11369(N35077,R3);
not not11370(N35091,in0);
not not11371(N35092,R0);
not not11372(N35093,R1);
not not11373(N35107,in0);
not not11374(N35108,in1);
not not11375(N35109,R1);
not not11376(N35110,R2);
not not11377(N35123,in0);
not not11378(N35124,in1);
not not11379(N35125,in2);
not not11380(N35126,R0);
not not11381(N35127,R1);
not not11382(N35139,in0);
not not11383(N35140,in1);
not not11384(N35141,in2);
not not11385(N35142,R3);
not not11386(N35155,in0);
not not11387(N35156,R1);
not not11388(N35170,in0);
not not11389(N35171,in2);
not not11390(N35172,R2);
not not11391(N35173,R3);
not not11392(N35185,in0);
not not11393(N35186,in1);
not not11394(N35187,R2);
not not11395(N35200,in0);
not not11396(N35201,in1);
not not11397(N35202,R1);
not not11398(N35203,R2);
not not11399(N35215,in0);
not not11400(N35216,in2);
not not11401(N35217,R1);
not not11402(N35218,R2);
not not11403(N35230,in0);
not not11404(N35231,in2);
not not11405(N35232,R0);
not not11406(N35233,R2);
not not11407(N35245,in0);
not not11408(N35246,in1);
not not11409(N35247,R1);
not not11410(N35248,R3);
not not11411(N35260,in0);
not not11412(N35261,in1);
not not11413(N35262,in2);
not not11414(N35263,R2);
not not11415(N35275,in0);
not not11416(N35276,in1);
not not11417(N35277,R1);
not not11418(N35278,R3);
not not11419(N35290,in0);
not not11420(N35291,in2);
not not11421(N35292,R3);
not not11422(N35305,in0);
not not11423(N35306,in2);
not not11424(N35307,R1);
not not11425(N35308,R2);
not not11426(N35320,in0);
not not11427(N35321,in1);
not not11428(N35322,in2);
not not11429(N35335,in0);
not not11430(N35336,R1);
not not11431(N35337,R2);
not not11432(N35350,in0);
not not11433(N35351,in1);
not not11434(N35352,in2);
not not11435(N35353,R3);
not not11436(N35365,in1);
not not11437(N35366,in2);
not not11438(N35367,R1);
not not11439(N35368,R2);
not not11440(N35380,in0);
not not11441(N35381,R2);
not not11442(N35395,in0);
not not11443(N35396,in2);
not not11444(N35397,R0);
not not11445(N35398,R2);
not not11446(N35410,in0);
not not11447(N35411,in1);
not not11448(N35412,in2);
not not11449(N35413,R0);
not not11450(N35414,R1);
not not11451(N35425,in0);
not not11452(N35426,in2);
not not11453(N35427,R1);
not not11454(N35428,R2);
not not11455(N35440,in0);
not not11456(N35441,R0);
not not11457(N35442,R1);
not not11458(N35443,R2);
not not11459(N35455,in0);
not not11460(N35456,in2);
not not11461(N35457,R0);
not not11462(N35458,R2);
not not11463(N35470,in0);
not not11464(N35471,in1);
not not11465(N35472,R0);
not not11466(N35473,R2);
not not11467(N35485,in0);
not not11468(N35486,in2);
not not11469(N35487,R0);
not not11470(N35500,in0);
not not11471(N35501,in1);
not not11472(N35502,in2);
not not11473(N35503,R1);
not not11474(N35515,in0);
not not11475(N35516,in2);
not not11476(N35517,R1);
not not11477(N35518,R3);
not not11478(N35530,in0);
not not11479(N35531,in1);
not not11480(N35532,in2);
not not11481(N35533,R2);
not not11482(N35545,in0);
not not11483(N35546,in1);
not not11484(N35547,R0);
not not11485(N35548,R1);
not not11486(N35560,in0);
not not11487(N35561,R0);
not not11488(N35562,R1);
not not11489(N35563,R2);
not not11490(N35575,in0);
not not11491(N35576,in1);
not not11492(N35577,R1);
not not11493(N35590,in0);
not not11494(N35591,in2);
not not11495(N35592,R0);
not not11496(N35605,in0);
not not11497(N35606,R0);
not not11498(N35607,R2);
not not11499(N35619,in0);
not not11500(N35620,in1);
not not11501(N35621,R2);
not not11502(N35633,in0);
not not11503(N35634,R1);
not not11504(N35647,in0);
not not11505(N35648,R1);
not not11506(N35649,R2);
not not11507(N35661,in0);
not not11508(N35662,in2);
not not11509(N35663,R2);
not not11510(N35675,in0);
not not11511(N35676,in1);
not not11512(N35677,in2);
not not11513(N35678,R0);
not not11514(N35689,in0);
not not11515(N35690,R0);
not not11516(N35691,R2);
not not11517(N35703,in0);
not not11518(N35704,in1);
not not11519(N35705,R2);
not not11520(N35717,in0);
not not11521(N35718,in1);
not not11522(N35719,R0);
not not11523(N35731,in0);
not not11524(N35732,in2);
not not11525(N35733,R1);
not not11526(N35745,in0);
not not11527(N35746,in2);
not not11528(N35747,R1);
not not11529(N35759,in0);
not not11530(N35760,in1);
not not11531(N35773,in0);
not not11532(N35774,in1);
not not11533(N35775,in2);
not not11534(N35776,R2);
not not11535(N35787,in0);
not not11536(N35788,R0);
not not11537(N35801,in0);
not not11538(N35802,in1);
not not11539(N35803,R0);
not not11540(N35804,R2);
not not11541(N35815,in0);
not not11542(N35816,in1);
not not11543(N35817,R0);
not not11544(N35829,in0);
not not11545(N35830,in1);
not not11546(N35831,in2);
not not11547(N35832,R1);
not not11548(N35843,in0);
not not11549(N35844,R0);
not not11550(N35845,R1);
not not11551(N35857,in0);
not not11552(N35858,R0);
not not11553(N35871,in0);
not not11554(N35872,R0);
not not11555(N35885,in0);
not not11556(N35886,R1);
not not11557(N35887,R2);
not not11558(N35899,in0);
not not11559(N35900,R0);
not not11560(N35901,R1);
not not11561(N35913,in1);
not not11562(N35914,R1);
not not11563(N35915,R3);
not not11564(N35927,in2);
not not11565(N35928,R1);
not not11566(N35929,R3);
not not11567(N35941,in0);
not not11568(N35942,in1);
not not11569(N35943,R1);
not not11570(N35955,in1);
not not11571(N35956,R0);
not not11572(N35957,R2);
not not11573(N35969,in2);
not not11574(N35970,R0);
not not11575(N35971,R2);
not not11576(N35983,in0);
not not11577(N35984,R0);
not not11578(N35985,R1);
not not11579(N35997,in0);
not not11580(N35998,in1);
not not11581(N35999,in2);
not not11582(N36011,in0);
not not11583(N36012,R0);
not not11584(N36013,R2);
not not11585(N36025,in0);
not not11586(N36026,in1);
not not11587(N36027,in2);
not not11588(N36028,R2);
not not11589(N36039,in0);
not not11590(N36040,R2);
not not11591(N36053,in0);
not not11592(N36054,in1);
not not11593(N36055,R0);
not not11594(N36067,in0);
not not11595(N36068,R2);
not not11596(N36069,R3);
not not11597(N36081,in0);
not not11598(N36082,in2);
not not11599(N36083,R0);
not not11600(N36084,R1);
not not11601(N36095,in0);
not not11602(N36096,R0);
not not11603(N36109,in0);
not not11604(N36110,in2);
not not11605(N36111,R2);
not not11606(N36123,in0);
not not11607(N36124,in1);
not not11608(N36125,in2);
not not11609(N36137,in0);
not not11610(N36138,in2);
not not11611(N36151,in0);
not not11612(N36152,in1);
not not11613(N36153,in2);
not not11614(N36165,in0);
not not11615(N36166,R0);
not not11616(N36167,R1);
not not11617(N36168,R3);
not not11618(N36179,in0);
not not11619(N36180,R1);
not not11620(N36193,in0);
not not11621(N36194,in1);
not not11622(N36195,R1);
not not11623(N36206,in0);
not not11624(N36207,R0);
not not11625(N36219,in0);
not not11626(N36220,R0);
not not11627(N36221,R2);
not not11628(N36232,in0);
not not11629(N36233,in1);
not not11630(N36234,R2);
not not11631(N36245,in0);
not not11632(N36246,in2);
not not11633(N36247,R1);
not not11634(N36258,in0);
not not11635(N36259,in1);
not not11636(N36260,R1);
not not11637(N36271,in0);
not not11638(N36272,in2);
not not11639(N36273,R3);
not not11640(N36284,in0);
not not11641(N36285,in2);
not not11642(N36286,R1);
not not11643(N36297,in0);
not not11644(N36298,in1);
not not11645(N36299,R2);
not not11646(N36310,in0);
not not11647(N36311,R2);
not not11648(N36323,in0);
not not11649(N36336,in0);
not not11650(N36337,in1);
not not11651(N36338,in2);
not not11652(N36339,R1);
not not11653(N36349,R1);
not not11654(N36350,R2);
not not11655(N36362,R1);
not not11656(N36363,R2);
not not11657(N36375,in0);
not not11658(N36376,in1);
not not11659(N36388,in0);
not not11660(N36389,R0);
not not11661(N36401,in0);
not not11662(N36402,in1);
not not11663(N36403,R1);
not not11664(N36414,in0);
not not11665(N36415,in1);
not not11666(N36416,R2);
not not11667(N36427,in0);
not not11668(N36428,in1);
not not11669(N36429,R1);
not not11670(N36440,in0);
not not11671(N36441,in2);
not not11672(N36442,R1);
not not11673(N36453,in0);
not not11674(N36454,R2);
not not11675(N36455,R3);
not not11676(N36466,in0);
not not11677(N36467,in1);
not not11678(N36468,in2);
not not11679(N36479,in0);
not not11680(N36480,in2);
not not11681(N36481,R0);
not not11682(N36482,R2);
not not11683(N36492,in0);
not not11684(N36505,in0);
not not11685(N36506,in1);
not not11686(N36507,R3);
not not11687(N36518,in0);
not not11688(N36519,R0);
not not11689(N36520,R1);
not not11690(N36531,in0);
not not11691(N36532,in2);
not not11692(N36533,R2);
not not11693(N36544,in0);
not not11694(N36545,in1);
not not11695(N36546,R0);
not not11696(N36557,in0);
not not11697(N36558,in2);
not not11698(N36559,R1);
not not11699(N36570,in0);
not not11700(N36571,R1);
not not11701(N36572,R2);
not not11702(N36583,in0);
not not11703(N36584,R2);
not not11704(N36596,in0);
not not11705(N36597,R1);
not not11706(N36598,R2);
not not11707(N36609,R1);
not not11708(N36610,R3);
not not11709(N36622,R0);
not not11710(N36623,R2);
not not11711(N36635,in0);
not not11712(N36636,R2);
not not11713(N36648,in0);
not not11714(N36649,in1);
not not11715(N36650,R2);
not not11716(N36660,in0);
not not11717(N36672,in0);
not not11718(N36673,in1);
not not11719(N36674,R1);
not not11720(N36684,in0);
not not11721(N36685,R3);
not not11722(N36696,in0);
not not11723(N36708,in0);
not not11724(N36709,in1);
not not11725(N36710,R0);
not not11726(N36720,in0);
not not11727(N36721,R0);
not not11728(N36732,in0);
not not11729(N36733,in2);
not not11730(N36744,in0);
not not11731(N36745,in2);
not not11732(N36756,in0);
not not11733(N36757,R3);
not not11734(N36767,in0);
not not11735(N36768,R1);
not not11736(N36778,in0);
not not11737(N36779,R3);
not not11738(N36789,in0);
not not11739(N36800,in0);
not not11740(N36801,R1);
not not11741(N36811,in0);
not not11742(N36821,in0);
not not11743(N36822,in1);
not not11744(N36823,R1);
not not11745(N36824,R2);
not not11746(N36825,R3);
not not11747(N36836,in0);
not not11748(N36837,in1);
not not11749(N36838,in2);
not not11750(N36839,R2);
not not11751(N36840,R5);
not not11752(N36851,in0);
not not11753(N36852,in1);
not not11754(N36853,R1);
not not11755(N36854,R3);
not not11756(N36855,R4);
not not11757(N36856,R5);
not not11758(N36866,in0);
not not11759(N36867,in1);
not not11760(N36868,R1);
not not11761(N36869,R4);
not not11762(N36870,R5);
not not11763(N36881,in0);
not not11764(N36882,in2);
not not11765(N36883,R1);
not not11766(N36884,R3);
not not11767(N36885,R4);
not not11768(N36886,R5);
not not11769(N36896,in0);
not not11770(N36897,R0);
not not11771(N36898,R2);
not not11772(N36899,R5);
not not11773(N36910,in0);
not not11774(N36911,R0);
not not11775(N36912,R1);
not not11776(N36913,R5);
not not11777(N36924,in0);
not not11778(N36925,R0);
not not11779(N36926,R1);
not not11780(N36927,R2);
not not11781(N36938,in0);
not not11782(N36939,in2);
not not11783(N36940,R4);
not not11784(N36941,R5);
not not11785(N36952,R0);
not not11786(N36953,R1);
not not11787(N36954,R3);
not not11788(N36955,R4);
not not11789(N36956,R5);
not not11790(N36966,R0);
not not11791(N36967,R2);
not not11792(N36968,R3);
not not11793(N36969,R4);
not not11794(N36980,R0);
not not11795(N36981,R1);
not not11796(N36982,R2);
not not11797(N36983,R4);
not not11798(N36994,in0);
not not11799(N36995,R1);
not not11800(N36996,R3);
not not11801(N36997,R5);
not not11802(N37008,in0);
not not11803(N37009,in1);
not not11804(N37010,in2);
not not11805(N37011,R2);
not not11806(N37012,R3);
not not11807(N37022,in0);
not not11808(N37023,in2);
not not11809(N37024,R0);
not not11810(N37025,R4);
not not11811(N37036,in0);
not not11812(N37037,in2);
not not11813(N37038,R0);
not not11814(N37039,R1);
not not11815(N37050,in0);
not not11816(N37051,in1);
not not11817(N37052,in2);
not not11818(N37053,R2);
not not11819(N37063,in0);
not not11820(N37064,in2);
not not11821(N37065,R0);
not not11822(N37066,R2);
not not11823(N37076,R1);
not not11824(N37077,R2);
not not11825(N37078,R3);
not not11826(N37079,R5);
not not11827(N37089,R1);
not not11828(N37090,R2);
not not11829(N37091,R3);
not not11830(N37092,R5);
not not11831(N37102,R1);
not not11832(N37103,R2);
not not11833(N37104,R5);
not not11834(N37115,in0);
not not11835(N37116,in2);
not not11836(N37127,in0);
not not11837(N37128,in2);
not not11838(N37129,R0);
not not11839(N37130,R4);
not not11840(N37139,in0);
not not11841(N37140,in2);
not not11842(N37141,R5);
not not11843(N37151,in0);
not not11844(N37152,R3);
not not11845(N37153,R4);
not not11846(N37163,in0);
not not11847(N37164,in2);
not not11848(N37165,R3);
not not11849(N37175,in0);
not not11850(N37176,in1);
not not11851(N37177,R3);
not not11852(N37187,in0);
not not11853(N37188,R0);
not not11854(N37198,in0);
not not11855(N37199,in1);
not not11856(N37200,R0);
not not11857(N37209,in0);
not not11858(N37210,R0);
not not11859(N37220,in0);
not not11860(N37221,in1);
not not11861(N37230,R4);
not not11862(N37231,R5);
not not11863(N37240,in0);
not not11864(N37241,R0);
not not11865(N37249,R0);
not not11866(N37250,R2);
not not11867(N37251,R3);
not not11868(N37252,R5);
not not11869(N37260,R0);
not not11870(N37261,R1);
not not11871(N37262,R3);
not not11872(N37263,R6);
not not11873(N34596,R2);
not not11874(N34597,R3);
not not11875(N34598,R4);
not not11876(N34599,R5);
not not11877(N34600,R6);
not not11878(N34601,R7);
not not11879(N34615,R3);
not not11880(N34616,R4);
not not11881(N34617,R5);
not not11882(N34618,R6);
not not11883(N34619,R7);
not not11884(N34635,R4);
not not11885(N34636,R7);
not not11886(N34652,R4);
not not11887(N34653,R5);
not not11888(N34654,R6);
not not11889(N34669,R3);
not not11890(N34670,R4);
not not11891(N34671,R5);
not not11892(N34672,R7);
not not11893(N34687,R3);
not not11894(N34688,R4);
not not11895(N34689,R5);
not not11896(N34690,R7);
not not11897(N34706,R4);
not not11898(N34707,R5);
not not11899(N34708,R7);
not not11900(N34723,R3);
not not11901(N34724,R5);
not not11902(N34725,R6);
not not11903(N34726,R7);
not not11904(N34741,R4);
not not11905(N34742,R6);
not not11906(N34743,R7);
not not11907(N34758,R4);
not not11908(N34759,R5);
not not11909(N34760,R6);
not not11910(N34774,R3);
not not11911(N34775,R4);
not not11912(N34776,R6);
not not11913(N34777,R7);
not not11914(N34792,R5);
not not11915(N34793,R6);
not not11916(N34806,R4);
not not11917(N34807,R5);
not not11918(N34808,R6);
not not11919(N34809,R7);
not not11920(N34823,R4);
not not11921(N34824,R6);
not not11922(N34825,R7);
not not11923(N34839,R4);
not not11924(N34840,R6);
not not11925(N34841,R7);
not not11926(N34855,R4);
not not11927(N34856,R5);
not not11928(N34857,R7);
not not11929(N34871,R4);
not not11930(N34872,R5);
not not11931(N34873,R6);
not not11932(N34887,R4);
not not11933(N34888,R5);
not not11934(N34889,R6);
not not11935(N34903,R4);
not not11936(N34904,R5);
not not11937(N34905,R6);
not not11938(N34919,R4);
not not11939(N34920,R5);
not not11940(N34921,R7);
not not11941(N34936,R4);
not not11942(N34937,R5);
not not11943(N34952,R6);
not not11944(N34953,R7);
not not11945(N34967,R4);
not not11946(N34968,R5);
not not11947(N34969,R7);
not not11948(N34983,R4);
not not11949(N34984,R5);
not not11950(N34985,R7);
not not11951(N34999,R4);
not not11952(N35000,R5);
not not11953(N35001,R7);
not not11954(N35016,R4);
not not11955(N35017,R6);
not not11956(N35032,R4);
not not11957(N35033,R5);
not not11958(N35048,R5);
not not11959(N35049,R7);
not not11960(N35064,R5);
not not11961(N35065,R7);
not not11962(N35078,R4);
not not11963(N35079,R5);
not not11964(N35080,R6);
not not11965(N35081,R7);
not not11966(N35094,R3);
not not11967(N35095,R5);
not not11968(N35096,R6);
not not11969(N35097,R7);
not not11970(N35111,R5);
not not11971(N35112,R6);
not not11972(N35113,R7);
not not11973(N35128,R4);
not not11974(N35129,R5);
not not11975(N35143,R4);
not not11976(N35144,R6);
not not11977(N35145,R7);
not not11978(N35157,R4);
not not11979(N35158,R5);
not not11980(N35159,R6);
not not11981(N35160,R7);
not not11982(N35174,R4);
not not11983(N35175,R7);
not not11984(N35188,R4);
not not11985(N35189,R5);
not not11986(N35190,R6);
not not11987(N35204,R4);
not not11988(N35205,R7);
not not11989(N35219,R4);
not not11990(N35220,R6);
not not11991(N35234,R6);
not not11992(N35235,R7);
not not11993(N35249,R5);
not not11994(N35250,R7);
not not11995(N35264,R4);
not not11996(N35265,R7);
not not11997(N35279,R5);
not not11998(N35280,R7);
not not11999(N35293,R5);
not not12000(N35294,R6);
not not12001(N35295,R7);
not not12002(N35309,R4);
not not12003(N35310,R6);
not not12004(N35323,R3);
not not12005(N35324,R4);
not not12006(N35325,R7);
not not12007(N35338,R4);
not not12008(N35339,R5);
not not12009(N35340,R7);
not not12010(N35354,R4);
not not12011(N35355,R5);
not not12012(N35369,R4);
not not12013(N35370,R5);
not not12014(N35382,R3);
not not12015(N35383,R5);
not not12016(N35384,R6);
not not12017(N35385,R7);
not not12018(N35399,R3);
not not12019(N35400,R7);
not not12020(N35415,R5);
not not12021(N35429,R5);
not not12022(N35430,R7);
not not12023(N35444,R4);
not not12024(N35445,R7);
not not12025(N35459,R5);
not not12026(N35460,R7);
not not12027(N35474,R5);
not not12028(N35475,R7);
not not12029(N35488,R3);
not not12030(N35489,R5);
not not12031(N35490,R6);
not not12032(N35504,R5);
not not12033(N35505,R6);
not not12034(N35519,R6);
not not12035(N35520,R7);
not not12036(N35534,R3);
not not12037(N35535,R7);
not not12038(N35549,R3);
not not12039(N35550,R6);
not not12040(N35564,R6);
not not12041(N35565,R7);
not not12042(N35578,R3);
not not12043(N35579,R4);
not not12044(N35580,R6);
not not12045(N35593,R3);
not not12046(N35594,R5);
not not12047(N35595,R7);
not not12048(N35608,R4);
not not12049(N35609,R5);
not not12050(N35622,R3);
not not12051(N35623,R7);
not not12052(N35635,R3);
not not12053(N35636,R5);
not not12054(N35637,R7);
not not12055(N35650,R5);
not not12056(N35651,R7);
not not12057(N35664,R4);
not not12058(N35665,R6);
not not12059(N35679,R3);
not not12060(N35692,R4);
not not12061(N35693,R7);
not not12062(N35706,R3);
not not12063(N35707,R6);
not not12064(N35720,R6);
not not12065(N35721,R7);
not not12066(N35734,R3);
not not12067(N35735,R5);
not not12068(N35748,R4);
not not12069(N35749,R7);
not not12070(N35761,R4);
not not12071(N35762,R5);
not not12072(N35763,R7);
not not12073(N35777,R5);
not not12074(N35789,R4);
not not12075(N35790,R5);
not not12076(N35791,R7);
not not12077(N35805,R7);
not not12078(N35818,R4);
not not12079(N35819,R6);
not not12080(N35833,R6);
not not12081(N35846,R4);
not not12082(N35847,R7);
not not12083(N35859,R3);
not not12084(N35860,R5);
not not12085(N35861,R6);
not not12086(N35873,R4);
not not12087(N35874,R6);
not not12088(N35875,R7);
not not12089(N35888,R4);
not not12090(N35889,R6);
not not12091(N35902,R4);
not not12092(N35903,R5);
not not12093(N35916,R4);
not not12094(N35917,R5);
not not12095(N35930,R4);
not not12096(N35931,R5);
not not12097(N35944,R3);
not not12098(N35945,R5);
not not12099(N35958,R4);
not not12100(N35959,R6);
not not12101(N35972,R4);
not not12102(N35973,R6);
not not12103(N35986,R4);
not not12104(N35987,R6);
not not12105(N36000,R4);
not not12106(N36001,R6);
not not12107(N36014,R4);
not not12108(N36015,R7);
not not12109(N36029,R5);
not not12110(N36041,R5);
not not12111(N36042,R6);
not not12112(N36043,R7);
not not12113(N36056,R5);
not not12114(N36057,R7);
not not12115(N36070,R4);
not not12116(N36071,R5);
not not12117(N36085,R5);
not not12118(N36097,R3);
not not12119(N36098,R4);
not not12120(N36099,R5);
not not12121(N36112,R6);
not not12122(N36113,R7);
not not12123(N36126,R4);
not not12124(N36127,R5);
not not12125(N36139,R4);
not not12126(N36140,R5);
not not12127(N36141,R7);
not not12128(N36154,R3);
not not12129(N36155,R4);
not not12130(N36169,R5);
not not12131(N36181,R3);
not not12132(N36182,R6);
not not12133(N36183,R7);
not not12134(N36196,R5);
not not12135(N36208,R4);
not not12136(N36209,R5);
not not12137(N36222,R5);
not not12138(N36235,R5);
not not12139(N36248,R4);
not not12140(N36261,R6);
not not12141(N36274,R6);
not not12142(N36287,R5);
not not12143(N36300,R5);
not not12144(N36312,R4);
not not12145(N36313,R6);
not not12146(N36324,R3);
not not12147(N36325,R4);
not not12148(N36326,R7);
not not12149(N36351,R4);
not not12150(N36352,R5);
not not12151(N36364,R4);
not not12152(N36365,R5);
not not12153(N36377,R3);
not not12154(N36378,R5);
not not12155(N36390,R4);
not not12156(N36391,R6);
not not12157(N36404,R7);
not not12158(N36417,R5);
not not12159(N36430,R7);
not not12160(N36443,R7);
not not12161(N36456,R6);
not not12162(N36469,R5);
not not12163(N36493,R4);
not not12164(N36494,R5);
not not12165(N36495,R6);
not not12166(N36508,R6);
not not12167(N36521,R7);
not not12168(N36534,R4);
not not12169(N36547,R4);
not not12170(N36560,R7);
not not12171(N36573,R6);
not not12172(N36585,R6);
not not12173(N36586,R7);
not not12174(N36599,R7);
not not12175(N36611,R4);
not not12176(N36612,R5);
not not12177(N36624,R4);
not not12178(N36625,R6);
not not12179(N36637,R4);
not not12180(N36638,R5);
not not12181(N36661,R4);
not not12182(N36662,R6);
not not12183(N36686,R5);
not not12184(N36697,R3);
not not12185(N36698,R6);
not not12186(N36722,R6);
not not12187(N36734,R5);
not not12188(N36746,R7);
not not12189(N36790,R3);
not not12190(N36812,R6);
not not12191(N36826,R6);
not not12192(N36827,R7);
not not12193(N36841,R6);
not not12194(N36842,R7);
not not12195(N36857,R6);
not not12196(N36871,R6);
not not12197(N36872,R7);
not not12198(N36887,R6);
not not12199(N36900,R6);
not not12200(N36901,R7);
not not12201(N36914,R6);
not not12202(N36915,R7);
not not12203(N36928,R5);
not not12204(N36929,R6);
not not12205(N36942,R6);
not not12206(N36943,R7);
not not12207(N36957,R7);
not not12208(N36970,R6);
not not12209(N36971,R7);
not not12210(N36984,R6);
not not12211(N36985,R7);
not not12212(N36998,R6);
not not12213(N36999,R7);
not not12214(N37013,R6);
not not12215(N37026,R5);
not not12216(N37027,R7);
not not12217(N37040,R5);
not not12218(N37041,R6);
not not12219(N37054,R7);
not not12220(N37067,R7);
not not12221(N37080,R6);
not not12222(N37093,R7);
not not12223(N37105,R6);
not not12224(N37106,R7);
not not12225(N37117,R6);
not not12226(N37118,R7);
not not12227(N37142,R6);
not not12228(N37154,R5);
not not12229(N37166,R6);
not not12230(N37178,R6);
not not12231(N37189,R5);
not not12232(N37211,R7);
not not12233(N37338,R0);
not not12234(N37350,R0);
not not12235(N37362,R0);
not not12236(N37374,R0);
not not12237(N37386,R0);
not not12238(N37398,R0);
not not12239(N37421,R0);
not not12240(N37432,R1);
not not12241(N37454,R0);
not not12242(N37465,R0);
not not12243(N37476,R0);
not not12244(N37487,R0);
not not12245(N37509,R0);
not not12246(N37520,R0);
not not12247(N37531,R1);
not not12248(N37542,R0);
not not12249(N37552,R0);
not not12250(N37572,R0);
not not12251(N37582,R0);
not not12252(N37592,R0);
not not12253(N37602,R0);
not not12254(N37612,R0);
not not12255(N37622,R0);
not not12256(N37632,R0);
not not12257(N37687,R0);
not not12258(N37741,R0);
not not12259(N37750,R1);
not not12260(N37776,R0);
not not12261(N37800,R0);
not not12262(N37816,R0);
not not12263(N37872,R2);
not not12264(N37881,R2);
not not12265(N37329,R1);
not not12266(N37330,R3);
not not12267(N37331,R7);
not not12268(N37339,R3);
not not12269(N37340,R4);
not not12270(N37341,R5);
not not12271(N37342,R6);
not not12272(N37343,R7);
not not12273(N37351,R1);
not not12274(N37352,R2);
not not12275(N37353,R3);
not not12276(N37354,R5);
not not12277(N37355,R6);
not not12278(N37363,R2);
not not12279(N37364,R3);
not not12280(N37365,R4);
not not12281(N37366,R5);
not not12282(N37367,R7);
not not12283(N37375,R1);
not not12284(N37376,R2);
not not12285(N37377,R3);
not not12286(N37378,R6);
not not12287(N37379,R7);
not not12288(N37387,R1);
not not12289(N37388,R3);
not not12290(N37389,R4);
not not12291(N37390,R6);
not not12292(N37391,R7);
not not12293(N37399,R1);
not not12294(N37400,R3);
not not12295(N37401,R4);
not not12296(N37402,R5);
not not12297(N37403,R6);
not not12298(N37410,R1);
not not12299(N37411,R2);
not not12300(N37412,R4);
not not12301(N37413,R6);
not not12302(N37414,R7);
not not12303(N37422,R1);
not not12304(N37423,R2);
not not12305(N37424,R4);
not not12306(N37425,R6);
not not12307(N37433,R4);
not not12308(N37434,R5);
not not12309(N37435,R6);
not not12310(N37436,R7);
not not12311(N37443,R1);
not not12312(N37444,R3);
not not12313(N37445,R4);
not not12314(N37446,R5);
not not12315(N37447,R7);
not not12316(N37455,R1);
not not12317(N37456,R3);
not not12318(N37457,R5);
not not12319(N37458,R7);
not not12320(N37466,R2);
not not12321(N37467,R3);
not not12322(N37468,R4);
not not12323(N37469,R7);
not not12324(N37477,R1);
not not12325(N37478,R2);
not not12326(N37479,R4);
not not12327(N37480,R7);
not not12328(N37488,R2);
not not12329(N37489,R5);
not not12330(N37490,R6);
not not12331(N37491,R7);
not not12332(N37498,R2);
not not12333(N37499,R3);
not not12334(N37500,R4);
not not12335(N37501,R5);
not not12336(N37502,R6);
not not12337(N37510,R1);
not not12338(N37511,R5);
not not12339(N37512,R6);
not not12340(N37513,R7);
not not12341(N37521,R1);
not not12342(N37522,R3);
not not12343(N37523,R6);
not not12344(N37524,R7);
not not12345(N37532,R2);
not not12346(N37533,R3);
not not12347(N37534,R6);
not not12348(N37535,R7);
not not12349(N37543,R4);
not not12350(N37544,R5);
not not12351(N37545,R6);
not not12352(N37553,R1);
not not12353(N37554,R4);
not not12354(N37555,R5);
not not12355(N37562,R3);
not not12356(N37563,R5);
not not12357(N37564,R6);
not not12358(N37565,R7);
not not12359(N37573,R2);
not not12360(N37574,R4);
not not12361(N37575,R5);
not not12362(N37583,R1);
not not12363(N37584,R2);
not not12364(N37585,R5);
not not12365(N37593,R2);
not not12366(N37594,R5);
not not12367(N37595,R6);
not not12368(N37603,R2);
not not12369(N37604,R3);
not not12370(N37605,R5);
not not12371(N37613,R3);
not not12372(N37614,R4);
not not12373(N37615,R5);
not not12374(N37623,R2);
not not12375(N37624,R3);
not not12376(N37625,R7);
not not12377(N37633,R3);
not not12378(N37634,R4);
not not12379(N37635,R7);
not not12380(N37642,R2);
not not12381(N37643,R4);
not not12382(N37644,R7);
not not12383(N37651,R1);
not not12384(N37652,R4);
not not12385(N37653,R6);
not not12386(N37660,R1);
not not12387(N37661,R4);
not not12388(N37662,R7);
not not12389(N37669,R3);
not not12390(N37670,R4);
not not12391(N37671,R6);
not not12392(N37678,R4);
not not12393(N37679,R5);
not not12394(N37680,R7);
not not12395(N37688,R1);
not not12396(N37689,R6);
not not12397(N37696,R3);
not not12398(N37697,R4);
not not12399(N37698,R6);
not not12400(N37705,R1);
not not12401(N37706,R3);
not not12402(N37707,R5);
not not12403(N37714,R1);
not not12404(N37715,R4);
not not12405(N37716,R6);
not not12406(N37723,R2);
not not12407(N37724,R3);
not not12408(N37725,R5);
not not12409(N37732,R2);
not not12410(N37733,R3);
not not12411(N37734,R5);
not not12412(N37742,R2);
not not12413(N37743,R6);
not not12414(N37751,R3);
not not12415(N37752,R5);
not not12416(N37759,R5);
not not12417(N37760,R6);
not not12418(N37761,R7);
not not12419(N37768,R1);
not not12420(N37769,R5);
not not12421(N37777,R1);
not not12422(N37784,R2);
not not12423(N37785,R6);
not not12424(N37792,R4);
not not12425(N37793,R5);
not not12426(N37801,R7);
not not12427(N37808,R1);
not not12428(N37809,R5);
not not12429(N37817,R4);
not not12430(N37824,R3);
not not12431(N37831,R3);
not not12432(N37838,R1);
not not12433(N37845,R3);
not not12434(N37852,R5);
not not12435(N37859,R7);
not not12436(N37866,R6);
not not12437(N37873,R5);
not not12438(N37874,R6);
not not12439(N37875,R7);
not not12440(N37934,R0);
not not12441(N37945,R0);
not not12442(N37956,R1);
not not12443(N37967,R0);
not not12444(N38019,R0);
not not12445(N38029,R0);
not not12446(N38039,R0);
not not12447(N38058,R0);
not not12448(N38094,R0);
not not12449(N38130,R0);
not not12450(N38139,R0);
not not12451(N38187,R0);
not not12452(N38210,R0);
not not12453(N37920,R0);
not not12454(N37921,R1);
not not12455(N37922,R2);
not not12456(N37923,R3);
not not12457(N37924,R4);
not not12458(N37925,R5);
not not12459(N37926,R6);
not not12460(N37927,R7);
not not12461(N37935,R2);
not not12462(N37936,R4);
not not12463(N37937,R5);
not not12464(N37938,R7);
not not12465(N37946,R1);
not not12466(N37947,R2);
not not12467(N37948,R6);
not not12468(N37949,R7);
not not12469(N37957,R3);
not not12470(N37958,R5);
not not12471(N37959,R6);
not not12472(N37960,R7);
not not12473(N37968,R2);
not not12474(N37969,R4);
not not12475(N37970,R5);
not not12476(N37971,R7);
not not12477(N37978,R1);
not not12478(N37979,R3);
not not12479(N37980,R5);
not not12480(N37981,R6);
not not12481(N37982,R7);
not not12482(N37989,R2);
not not12483(N37990,R4);
not not12484(N37991,R5);
not not12485(N37992,R6);
not not12486(N37999,R3);
not not12487(N38000,R4);
not not12488(N38001,R6);
not not12489(N38002,R7);
not not12490(N38009,R1);
not not12491(N38010,R2);
not not12492(N38011,R5);
not not12493(N38012,R6);
not not12494(N38020,R1);
not not12495(N38021,R4);
not not12496(N38022,R7);
not not12497(N38030,R3);
not not12498(N38031,R5);
not not12499(N38032,R6);
not not12500(N38040,R1);
not not12501(N38041,R5);
not not12502(N38042,R6);
not not12503(N38049,R4);
not not12504(N38050,R6);
not not12505(N38051,R7);
not not12506(N38059,R2);
not not12507(N38060,R7);
not not12508(N38067,R2);
not not12509(N38068,R3);
not not12510(N38069,R6);
not not12511(N38076,R1);
not not12512(N38077,R4);
not not12513(N38078,R5);
not not12514(N38085,R2);
not not12515(N38086,R5);
not not12516(N38087,R7);
not not12517(N38095,R2);
not not12518(N38096,R7);
not not12519(N38103,R1);
not not12520(N38104,R3);
not not12521(N38105,R6);
not not12522(N38112,R3);
not not12523(N38113,R5);
not not12524(N38114,R7);
not not12525(N38121,R1);
not not12526(N38122,R6);
not not12527(N38123,R7);
not not12528(N38131,R5);
not not12529(N38132,R7);
not not12530(N38140,R5);
not not12531(N38147,R2);
not not12532(N38148,R5);
not not12533(N38155,R2);
not not12534(N38156,R7);
not not12535(N38163,R1);
not not12536(N38164,R6);
not not12537(N38171,R2);
not not12538(N38172,R5);
not not12539(N38179,R3);
not not12540(N38180,R5);
not not12541(N38188,R6);
not not12542(N38195,R3);
not not12543(N38196,R7);
not not12544(N38203,R6);
not not12545(N38204,R7);
not not12546(N38211,R3);
not not12547(N38212,R6);
not not12548(N38349,R1);
not not12549(N38360,R0);
not not12550(N38232,R0);
not not12551(N38233,R3);
not not12552(N38234,R5);
not not12553(N38235,R6);
not not12554(N38236,R7);
not not12555(N38244,R1);
not not12556(N38245,R2);
not not12557(N38246,R3);
not not12558(N38247,R5);
not not12559(N38248,R6);
not not12560(N38256,R0);
not not12561(N38257,R4);
not not12562(N38258,R5);
not not12563(N38259,R7);
not not12564(N38267,R0);
not not12565(N38268,R4);
not not12566(N38269,R6);
not not12567(N38270,R7);
not not12568(N38278,R1);
not not12569(N38279,R2);
not not12570(N38280,R4);
not not12571(N38281,R5);
not not12572(N38289,R0);
not not12573(N38290,R1);
not not12574(N38291,R6);
not not12575(N38292,R7);
not not12576(N38300,R0);
not not12577(N38301,R2);
not not12578(N38302,R4);
not not12579(N38303,R6);
not not12580(N38311,R2);
not not12581(N38312,R3);
not not12582(N38313,R7);
not not12583(N38321,R5);
not not12584(N38322,R6);
not not12585(N38330,R4);
not not12586(N38331,R7);
not not12587(N38338,R3);
not not12588(N38339,R4);
not not12589(N38340,R5);
not not12590(N38341,R6);
not not12591(N38342,R7);
not not12592(N38350,R2);
not not12593(N38351,R3);
not not12594(N38352,R5);
not not12595(N38353,R7);
not not12596(N38361,R1);
not not12597(N38362,R3);
not not12598(N38363,R6);
not not12599(N38424,R0);
not not12600(N38435,R0);
not not12601(N38446,R0);
not not12602(N38457,R1);
not not12603(N38488,R0);
not not12604(N38498,R0);
not not12605(N38508,R0);
not not12606(N38518,R0);
not not12607(N38528,R0);
not not12608(N38547,R0);
not not12609(N38583,R0);
not not12610(N38592,R0);
not not12611(N38610,R1);
not not12612(N38619,R1);
not not12613(N38637,R0);
not not12614(N38695,R0);
not not12615(N38727,R0);
not not12616(N38742,R0);
not not12617(N38760,R1);
not not12618(N38769,R1);
not not12619(N38410,R0);
not not12620(N38411,R1);
not not12621(N38412,R2);
not not12622(N38413,R3);
not not12623(N38414,R4);
not not12624(N38415,R5);
not not12625(N38416,R6);
not not12626(N38417,R7);
not not12627(N38425,R2);
not not12628(N38426,R4);
not not12629(N38427,R5);
not not12630(N38428,R7);
not not12631(N38436,R1);
not not12632(N38437,R2);
not not12633(N38438,R6);
not not12634(N38439,R7);
not not12635(N38447,R2);
not not12636(N38448,R4);
not not12637(N38449,R5);
not not12638(N38450,R7);
not not12639(N38458,R2);
not not12640(N38459,R3);
not not12641(N38460,R5);
not not12642(N38461,R7);
not not12643(N38468,R2);
not not12644(N38469,R4);
not not12645(N38470,R5);
not not12646(N38471,R6);
not not12647(N38478,R1);
not not12648(N38479,R2);
not not12649(N38480,R4);
not not12650(N38481,R5);
not not12651(N38489,R1);
not not12652(N38490,R4);
not not12653(N38491,R7);
not not12654(N38499,R3);
not not12655(N38500,R4);
not not12656(N38501,R6);
not not12657(N38509,R3);
not not12658(N38510,R6);
not not12659(N38511,R7);
not not12660(N38519,R2);
not not12661(N38520,R4);
not not12662(N38521,R6);
not not12663(N38529,R1);
not not12664(N38530,R5);
not not12665(N38531,R6);
not not12666(N38538,R4);
not not12667(N38539,R6);
not not12668(N38540,R7);
not not12669(N38548,R2);
not not12670(N38549,R7);
not not12671(N38556,R2);
not not12672(N38557,R3);
not not12673(N38558,R6);
not not12674(N38565,R1);
not not12675(N38566,R4);
not not12676(N38567,R5);
not not12677(N38574,R2);
not not12678(N38575,R5);
not not12679(N38576,R7);
not not12680(N38584,R2);
not not12681(N38585,R7);
not not12682(N38593,R4);
not not12683(N38594,R5);
not not12684(N38601,R4);
not not12685(N38602,R6);
not not12686(N38603,R7);
not not12687(N38611,R6);
not not12688(N38612,R7);
not not12689(N38620,R3);
not not12690(N38621,R6);
not not12691(N38628,R3);
not not12692(N38629,R5);
not not12693(N38630,R7);
not not12694(N38638,R5);
not not12695(N38639,R7);
not not12696(N38646,R1);
not not12697(N38647,R2);
not not12698(N38648,R6);
not not12699(N38655,R2);
not not12700(N38656,R5);
not not12701(N38663,R2);
not not12702(N38664,R7);
not not12703(N38671,R2);
not not12704(N38672,R5);
not not12705(N38679,R3);
not not12706(N38680,R7);
not not12707(N38687,R5);
not not12708(N38688,R6);
not not12709(N38696,R6);
not not12710(N38703,R4);
not not12711(N38704,R7);
not not12712(N38711,R6);
not not12713(N38712,R7);
not not12714(N38719,R1);
not not12715(N38720,R6);
not not12716(N38728,R5);
not not12717(N38735,R3);
not not12718(N38736,R5);
not not12719(N38743,R3);
not not12720(N38744,R5);
not not12721(N38745,R6);
not not12722(N38751,R3);
not not12723(N38752,R4);
not not12724(N38753,R6);
not not12725(N38754,R7);
not not12726(N38761,R3);
not not12727(N38762,R5);
not not12728(N38763,R6);
not not12729(N38770,R3);
not not12730(N38771,R6);
not not12731(N38982,R0);
not not12732(N38994,R0);
not not12733(N39017,R0);
not not12734(N38801,R0);
not not12735(N38802,R2);
not not12736(N38803,R3);
not not12737(N38804,R4);
not not12738(N38805,R6);
not not12739(N38806,R7);
not not12740(N38814,R0);
not not12741(N38815,R1);
not not12742(N38816,R2);
not not12743(N38817,R4);
not not12744(N38818,R6);
not not12745(N38819,R7);
not not12746(N38827,R1);
not not12747(N38828,R2);
not not12748(N38829,R3);
not not12749(N38830,R4);
not not12750(N38831,R5);
not not12751(N38832,R6);
not not12752(N38840,R1);
not not12753(N38841,R2);
not not12754(N38842,R5);
not not12755(N38843,R6);
not not12756(N38844,R7);
not not12757(N38852,R0);
not not12758(N38853,R1);
not not12759(N38854,R2);
not not12760(N38855,R5);
not not12761(N38863,R1);
not not12762(N38864,R4);
not not12763(N38865,R6);
not not12764(N38866,R7);
not not12765(N38874,R2);
not not12766(N38875,R3);
not not12767(N38876,R5);
not not12768(N38877,R7);
not not12769(N38885,R0);
not not12770(N38886,R2);
not not12771(N38887,R5);
not not12772(N38888,R6);
not not12773(N38896,R2);
not not12774(N38897,R3);
not not12775(N38898,R4);
not not12776(N38899,R5);
not not12777(N38907,R0);
not not12778(N38908,R2);
not not12779(N38909,R3);
not not12780(N38910,R6);
not not12781(N38918,R0);
not not12782(N38919,R1);
not not12783(N38920,R3);
not not12784(N38921,R5);
not not12785(N38929,R1);
not not12786(N38930,R5);
not not12787(N38931,R7);
not not12788(N38939,R1);
not not12789(N38940,R3);
not not12790(N38941,R7);
not not12791(N38949,R2);
not not12792(N38950,R4);
not not12793(N38958,R0);
not not12794(N38959,R2);
not not12795(N38967,R7);
not not12796(N38975,R6);
not not12797(N38983,R1);
not not12798(N38984,R2);
not not12799(N38985,R3);
not not12800(N38986,R6);
not not12801(N38987,R7);
not not12802(N38995,R2);
not not12803(N38996,R3);
not not12804(N38997,R5);
not not12805(N38998,R6);
not not12806(N38999,R7);
not not12807(N39006,R1);
not not12808(N39007,R2);
not not12809(N39008,R3);
not not12810(N39009,R6);
not not12811(N39010,R7);
not not12812(N39018,R4);
not not12813(N39019,R5);
not not12814(N39020,R6);
not not12815(N39027,R5);
not not12816(N39034,R3);
not not12817(N39105,R0);
not not12818(N39117,R0);
not not12819(N39129,R0);
not not12820(N39141,R0);
not not12821(N39153,R0);
not not12822(N39165,R0);
not not12823(N39176,R1);
not not12824(N39209,R0);
not not12825(N39220,R0);
not not12826(N39231,R0);
not not12827(N39242,R0);
not not12828(N39283,R0);
not not12829(N39303,R0);
not not12830(N39313,R0);
not not12831(N39333,R1);
not not12832(N39343,R0);
not not12833(N39353,R0);
not not12834(N39363,R0);
not not12835(N39373,R0);
not not12836(N39392,R1);
not not12837(N39454,R0);
not not12838(N39478,R0);
not not12839(N39486,R0);
not not12840(N39494,R0);
not not12841(N39525,R1);
not not12842(N39087,R4);
not not12843(N39088,R5);
not not12844(N39089,R6);
not not12845(N39097,R0);
not not12846(N39098,R3);
not not12847(N39106,R3);
not not12848(N39107,R4);
not not12849(N39108,R5);
not not12850(N39109,R6);
not not12851(N39110,R7);
not not12852(N39118,R1);
not not12853(N39119,R2);
not not12854(N39120,R3);
not not12855(N39121,R5);
not not12856(N39122,R6);
not not12857(N39130,R2);
not not12858(N39131,R3);
not not12859(N39132,R4);
not not12860(N39133,R5);
not not12861(N39134,R7);
not not12862(N39142,R1);
not not12863(N39143,R3);
not not12864(N39144,R4);
not not12865(N39145,R6);
not not12866(N39146,R7);
not not12867(N39154,R1);
not not12868(N39155,R3);
not not12869(N39156,R4);
not not12870(N39157,R5);
not not12871(N39158,R6);
not not12872(N39166,R1);
not not12873(N39167,R2);
not not12874(N39168,R4);
not not12875(N39169,R6);
not not12876(N39177,R4);
not not12877(N39178,R5);
not not12878(N39179,R6);
not not12879(N39180,R7);
not not12880(N39187,R2);
not not12881(N39188,R4);
not not12882(N39189,R5);
not not12883(N39190,R6);
not not12884(N39191,R7);
not not12885(N39198,R1);
not not12886(N39199,R3);
not not12887(N39200,R4);
not not12888(N39201,R5);
not not12889(N39202,R7);
not not12890(N39210,R1);
not not12891(N39211,R3);
not not12892(N39212,R5);
not not12893(N39213,R7);
not not12894(N39221,R1);
not not12895(N39222,R5);
not not12896(N39223,R6);
not not12897(N39224,R7);
not not12898(N39232,R1);
not not12899(N39233,R3);
not not12900(N39234,R6);
not not12901(N39235,R7);
not not12902(N39243,R1);
not not12903(N39244,R2);
not not12904(N39245,R5);
not not12905(N39246,R6);
not not12906(N39253,R2);
not not12907(N39254,R5);
not not12908(N39255,R6);
not not12909(N39256,R7);
not not12910(N39263,R2);
not not12911(N39264,R3);
not not12912(N39265,R4);
not not12913(N39266,R6);
not not12914(N39273,R1);
not not12915(N39274,R2);
not not12916(N39275,R4);
not not12917(N39276,R6);
not not12918(N39284,R1);
not not12919(N39285,R4);
not not12920(N39286,R5);
not not12921(N39293,R3);
not not12922(N39294,R5);
not not12923(N39295,R6);
not not12924(N39296,R7);
not not12925(N39304,R2);
not not12926(N39305,R4);
not not12927(N39306,R5);
not not12928(N39314,R2);
not not12929(N39315,R4);
not not12930(N39316,R5);
not not12931(N39323,R2);
not not12932(N39324,R3);
not not12933(N39325,R4);
not not12934(N39326,R7);
not not12935(N39334,R2);
not not12936(N39335,R4);
not not12937(N39336,R7);
not not12938(N39344,R2);
not not12939(N39345,R3);
not not12940(N39346,R5);
not not12941(N39354,R3);
not not12942(N39355,R4);
not not12943(N39356,R5);
not not12944(N39364,R2);
not not12945(N39365,R3);
not not12946(N39366,R7);
not not12947(N39374,R3);
not not12948(N39375,R4);
not not12949(N39376,R7);
not not12950(N39383,R4);
not not12951(N39384,R5);
not not12952(N39385,R7);
not not12953(N39393,R4);
not not12954(N39394,R6);
not not12955(N39401,R3);
not not12956(N39402,R4);
not not12957(N39403,R6);
not not12958(N39410,R1);
not not12959(N39411,R3);
not not12960(N39412,R5);
not not12961(N39419,R5);
not not12962(N39420,R6);
not not12963(N39421,R7);
not not12964(N39428,R2);
not not12965(N39429,R4);
not not12966(N39430,R7);
not not12967(N39437,R2);
not not12968(N39438,R3);
not not12969(N39439,R5);
not not12970(N39446,R1);
not not12971(N39447,R5);
not not12972(N39455,R1);
not not12973(N39462,R1);
not not12974(N39463,R4);
not not12975(N39470,R2);
not not12976(N39471,R6);
not not12977(N39479,R1);
not not12978(N39487,R7);
not not12979(N39495,R4);
not not12980(N39502,R2);
not not12981(N39503,R6);
not not12982(N39510,R3);
not not12983(N39511,R6);
not not12984(N39518,R2);

endmodule